
module mem_32_512_0 ( clk, addr_rd, wr_ena, data_rd, addr_wr, data_wr );
  input [8:0] addr_rd;
  output [31:0] data_rd;
  input [8:0] addr_wr;
  input [31:0] data_wr;
  input clk, wr_ena;

  wire   [8:0] int_addr;

  SRAM32x512_1rw SRAM_HM_01 ( .I(data_wr), .O(data_rd), .A(int_addr), .CE(1'b0), .CSB(1'b0), .WEB(wr_ena), .OEB(1'b0) );
  MUX21X1 U3 ( .IN1(addr_rd[0]), .IN2(addr_wr[0]), .S(wr_ena), .Q(int_addr[0])
         );
  MUX21X1 U4 ( .IN1(addr_rd[1]), .IN2(addr_wr[1]), .S(wr_ena), .Q(int_addr[1])
         );
  MUX21X1 U5 ( .IN1(addr_rd[2]), .IN2(addr_wr[2]), .S(wr_ena), .Q(int_addr[2])
         );
  MUX21X1 U6 ( .IN1(addr_rd[3]), .IN2(addr_wr[3]), .S(wr_ena), .Q(int_addr[3])
         );
  MUX21X1 U7 ( .IN1(addr_rd[4]), .IN2(addr_wr[4]), .S(wr_ena), .Q(int_addr[4])
         );
  MUX21X1 U8 ( .IN1(addr_rd[5]), .IN2(addr_wr[5]), .S(wr_ena), .Q(int_addr[5])
         );
  MUX21X1 U9 ( .IN1(addr_rd[6]), .IN2(addr_wr[6]), .S(wr_ena), .Q(int_addr[6])
         );
  MUX21X1 U10 ( .IN1(addr_rd[7]), .IN2(addr_wr[7]), .S(wr_ena), .Q(int_addr[7]) );
  MUX21X1 U11 ( .IN1(addr_rd[8]), .IN2(addr_wr[8]), .S(wr_ena), .Q(int_addr[8]) );
endmodule


module mem_32_512_4 ( clk, addr_rd, wr_ena, data_rd, addr_wr, data_wr );
  input [8:0] addr_rd;
  output [31:0] data_rd;
  input [8:0] addr_wr;
  input [31:0] data_wr;
  input clk, wr_ena;

  wire   [8:0] int_addr;

  SRAM32x512_1rw SRAM_HM_01 ( .I(data_wr), .O(data_rd), .A(int_addr), .CE(1'b0), .CSB(1'b0), .WEB(wr_ena), .OEB(1'b0) );
  MUX21X1 U3 ( .IN1(addr_rd[0]), .IN2(addr_wr[0]), .S(wr_ena), .Q(int_addr[0])
         );
  MUX21X1 U4 ( .IN1(addr_rd[1]), .IN2(addr_wr[1]), .S(wr_ena), .Q(int_addr[1])
         );
  MUX21X1 U5 ( .IN1(addr_rd[2]), .IN2(addr_wr[2]), .S(wr_ena), .Q(int_addr[2])
         );
  MUX21X1 U6 ( .IN1(addr_rd[3]), .IN2(addr_wr[3]), .S(wr_ena), .Q(int_addr[3])
         );
  MUX21X1 U7 ( .IN1(addr_rd[4]), .IN2(addr_wr[4]), .S(wr_ena), .Q(int_addr[4])
         );
  MUX21X1 U8 ( .IN1(addr_rd[5]), .IN2(addr_wr[5]), .S(wr_ena), .Q(int_addr[5])
         );
  MUX21X1 U9 ( .IN1(addr_rd[6]), .IN2(addr_wr[6]), .S(wr_ena), .Q(int_addr[6])
         );
  MUX21X1 U10 ( .IN1(addr_rd[7]), .IN2(addr_wr[7]), .S(wr_ena), .Q(int_addr[7]) );
  MUX21X1 U11 ( .IN1(addr_rd[8]), .IN2(addr_wr[8]), .S(wr_ena), .Q(int_addr[8]) );
endmodule


module mem_int ( clk, addr_rd, wr_ena, data_rd, addr_wr, data_wr );
  input [19:0] addr_rd;
  output [31:0] data_rd;
  input [19:0] addr_wr;
  input [31:0] data_wr;
  input clk, wr_ena;
  wire   wr_0, wr_1, n1;
  wire   [31:0] data_rd_1;
  wire   [31:0] data_rd_0;

  mem_32_512_0 mem_0 ( .clk(clk), .addr_rd(addr_rd[8:0]), .wr_ena(wr_0), 
        .data_rd(data_rd_0), .addr_wr(addr_wr[8:0]), .data_wr(data_wr) );
  mem_32_512_4 mem_1 ( .clk(clk), .addr_rd(addr_rd[8:0]), .wr_ena(wr_1), 
        .data_rd(data_rd_1), .addr_wr(addr_wr[8:0]), .data_wr(data_wr) );
  NOR2X0 U1 ( .IN1(addr_wr[9]), .IN2(n1), .QN(wr_0) );
  AND2X1 U2 ( .IN1(addr_wr[9]), .IN2(wr_ena), .Q(wr_1) );
  MUX21X1 U3 ( .IN1(data_rd_0[0]), .IN2(data_rd_1[0]), .S(addr_rd[9]), .Q(
        data_rd[0]) );
  MUX21X1 U4 ( .IN1(data_rd_0[10]), .IN2(data_rd_1[10]), .S(addr_rd[9]), .Q(
        data_rd[10]) );
  MUX21X1 U5 ( .IN1(data_rd_0[11]), .IN2(data_rd_1[11]), .S(addr_rd[9]), .Q(
        data_rd[11]) );
  MUX21X1 U6 ( .IN1(data_rd_0[12]), .IN2(data_rd_1[12]), .S(addr_rd[9]), .Q(
        data_rd[12]) );
  MUX21X1 U7 ( .IN1(data_rd_0[13]), .IN2(data_rd_1[13]), .S(addr_rd[9]), .Q(
        data_rd[13]) );
  MUX21X1 U8 ( .IN1(data_rd_0[14]), .IN2(data_rd_1[14]), .S(addr_rd[9]), .Q(
        data_rd[14]) );
  MUX21X1 U9 ( .IN1(data_rd_0[15]), .IN2(data_rd_1[15]), .S(addr_rd[9]), .Q(
        data_rd[15]) );
  MUX21X1 U10 ( .IN1(data_rd_0[16]), .IN2(data_rd_1[16]), .S(addr_rd[9]), .Q(
        data_rd[16]) );
  MUX21X1 U11 ( .IN1(data_rd_0[17]), .IN2(data_rd_1[17]), .S(addr_rd[9]), .Q(
        data_rd[17]) );
  MUX21X1 U12 ( .IN1(data_rd_0[18]), .IN2(data_rd_1[18]), .S(addr_rd[9]), .Q(
        data_rd[18]) );
  MUX21X1 U13 ( .IN1(data_rd_0[19]), .IN2(data_rd_1[19]), .S(addr_rd[9]), .Q(
        data_rd[19]) );
  MUX21X1 U14 ( .IN1(data_rd_0[1]), .IN2(data_rd_1[1]), .S(addr_rd[9]), .Q(
        data_rd[1]) );
  MUX21X1 U15 ( .IN1(data_rd_0[20]), .IN2(data_rd_1[20]), .S(addr_rd[9]), .Q(
        data_rd[20]) );
  MUX21X1 U16 ( .IN1(data_rd_0[21]), .IN2(data_rd_1[21]), .S(addr_rd[9]), .Q(
        data_rd[21]) );
  MUX21X1 U17 ( .IN1(data_rd_0[22]), .IN2(data_rd_1[22]), .S(addr_rd[9]), .Q(
        data_rd[22]) );
  MUX21X1 U18 ( .IN1(data_rd_0[23]), .IN2(data_rd_1[23]), .S(addr_rd[9]), .Q(
        data_rd[23]) );
  MUX21X1 U19 ( .IN1(data_rd_0[24]), .IN2(data_rd_1[24]), .S(addr_rd[9]), .Q(
        data_rd[24]) );
  MUX21X1 U20 ( .IN1(data_rd_0[25]), .IN2(data_rd_1[25]), .S(addr_rd[9]), .Q(
        data_rd[25]) );
  MUX21X1 U21 ( .IN1(data_rd_0[26]), .IN2(data_rd_1[26]), .S(addr_rd[9]), .Q(
        data_rd[26]) );
  MUX21X1 U22 ( .IN1(data_rd_0[27]), .IN2(data_rd_1[27]), .S(addr_rd[9]), .Q(
        data_rd[27]) );
  MUX21X1 U23 ( .IN1(data_rd_0[28]), .IN2(data_rd_1[28]), .S(addr_rd[9]), .Q(
        data_rd[28]) );
  MUX21X1 U24 ( .IN1(data_rd_0[29]), .IN2(data_rd_1[29]), .S(addr_rd[9]), .Q(
        data_rd[29]) );
  MUX21X1 U25 ( .IN1(data_rd_0[2]), .IN2(data_rd_1[2]), .S(addr_rd[9]), .Q(
        data_rd[2]) );
  MUX21X1 U26 ( .IN1(data_rd_0[30]), .IN2(data_rd_1[30]), .S(addr_rd[9]), .Q(
        data_rd[30]) );
  MUX21X1 U27 ( .IN1(data_rd_0[31]), .IN2(data_rd_1[31]), .S(addr_rd[9]), .Q(
        data_rd[31]) );
  MUX21X1 U28 ( .IN1(data_rd_0[3]), .IN2(data_rd_1[3]), .S(addr_rd[9]), .Q(
        data_rd[3]) );
  MUX21X1 U29 ( .IN1(data_rd_0[4]), .IN2(data_rd_1[4]), .S(addr_rd[9]), .Q(
        data_rd[4]) );
  MUX21X1 U30 ( .IN1(data_rd_0[5]), .IN2(data_rd_1[5]), .S(addr_rd[9]), .Q(
        data_rd[5]) );
  MUX21X1 U31 ( .IN1(data_rd_0[6]), .IN2(data_rd_1[6]), .S(addr_rd[9]), .Q(
        data_rd[6]) );
  MUX21X1 U32 ( .IN1(data_rd_0[7]), .IN2(data_rd_1[7]), .S(addr_rd[9]), .Q(
        data_rd[7]) );
  MUX21X1 U33 ( .IN1(data_rd_0[8]), .IN2(data_rd_1[8]), .S(addr_rd[9]), .Q(
        data_rd[8]) );
  MUX21X1 U34 ( .IN1(data_rd_0[9]), .IN2(data_rd_1[9]), .S(addr_rd[9]), .Q(
        data_rd[9]) );
  INVX0 U35 ( .INP(wr_ena), .ZN(n1) );
endmodule


module mem_32_512_2 ( clk, addr_rd, wr_ena, data_rd, addr_wr, data_wr );
  input [8:0] addr_rd;
  output [31:0] data_rd;
  input [8:0] addr_wr;
  input [31:0] data_wr;
  input clk, wr_ena;
  wire   SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20;
  wire   [8:0] int_addr;

  SRAM32x512_1rw SRAM_HM_01 ( .I(data_wr), .O({SYNOPSYS_UNCONNECTED_20, 
        SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_18, 
        SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_16, 
        SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_14, 
        SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_12, 
        SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_10, 
        SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_7, 
        SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_4, 
        SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_1, 
        data_rd[11:0]}), .A(int_addr), .CE(1'b0), .CSB(1'b0), .WEB(wr_ena), 
        .OEB(1'b0) );
  MUX21X1 U3 ( .IN1(addr_rd[0]), .IN2(addr_wr[0]), .S(wr_ena), .Q(int_addr[0])
         );
  MUX21X1 U4 ( .IN1(addr_rd[1]), .IN2(addr_wr[1]), .S(wr_ena), .Q(int_addr[1])
         );
  MUX21X1 U5 ( .IN1(addr_rd[2]), .IN2(addr_wr[2]), .S(wr_ena), .Q(int_addr[2])
         );
  MUX21X1 U6 ( .IN1(addr_rd[3]), .IN2(addr_wr[3]), .S(wr_ena), .Q(int_addr[3])
         );
  MUX21X1 U7 ( .IN1(addr_rd[4]), .IN2(addr_wr[4]), .S(wr_ena), .Q(int_addr[4])
         );
  MUX21X1 U8 ( .IN1(addr_rd[5]), .IN2(addr_wr[5]), .S(wr_ena), .Q(int_addr[5])
         );
  MUX21X1 U9 ( .IN1(addr_rd[6]), .IN2(addr_wr[6]), .S(wr_ena), .Q(int_addr[6])
         );
  MUX21X1 U10 ( .IN1(addr_rd[7]), .IN2(addr_wr[7]), .S(wr_ena), .Q(int_addr[7]) );
  MUX21X1 U11 ( .IN1(addr_rd[8]), .IN2(addr_wr[8]), .S(wr_ena), .Q(int_addr[8]) );
endmodule


module mem_32_512_3 ( clk, addr_rd, wr_ena, data_rd, addr_wr, data_wr );
  input [8:0] addr_rd;
  output [31:0] data_rd;
  input [8:0] addr_wr;
  input [31:0] data_wr;
  input clk, wr_ena;
  wire   SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20;
  wire   [8:0] int_addr;

  SRAM32x512_1rw SRAM_HM_01 ( .I(data_wr), .O({SYNOPSYS_UNCONNECTED_20, 
        SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_18, 
        SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_16, 
        SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_14, 
        SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_12, 
        SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_10, 
        SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_7, 
        SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_4, 
        SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_1, 
        data_rd[11:0]}), .A(int_addr), .CE(1'b0), .CSB(1'b0), .WEB(wr_ena), 
        .OEB(1'b0) );
  MUX21X1 U3 ( .IN1(addr_rd[0]), .IN2(addr_wr[0]), .S(wr_ena), .Q(int_addr[0])
         );
  MUX21X1 U4 ( .IN1(addr_rd[1]), .IN2(addr_wr[1]), .S(wr_ena), .Q(int_addr[1])
         );
  MUX21X1 U5 ( .IN1(addr_rd[2]), .IN2(addr_wr[2]), .S(wr_ena), .Q(int_addr[2])
         );
  MUX21X1 U6 ( .IN1(addr_rd[3]), .IN2(addr_wr[3]), .S(wr_ena), .Q(int_addr[3])
         );
  MUX21X1 U7 ( .IN1(addr_rd[4]), .IN2(addr_wr[4]), .S(wr_ena), .Q(int_addr[4])
         );
  MUX21X1 U8 ( .IN1(addr_rd[5]), .IN2(addr_wr[5]), .S(wr_ena), .Q(int_addr[5])
         );
  MUX21X1 U9 ( .IN1(addr_rd[6]), .IN2(addr_wr[6]), .S(wr_ena), .Q(int_addr[6])
         );
  MUX21X1 U10 ( .IN1(addr_rd[7]), .IN2(addr_wr[7]), .S(wr_ena), .Q(int_addr[7]) );
  MUX21X1 U11 ( .IN1(addr_rd[8]), .IN2(addr_wr[8]), .S(wr_ena), .Q(int_addr[8]) );
endmodule


module mem_interface ( clk, addr_rd, wr_ena, data_rd, addr_wr, data_wr );
  input [19:0] addr_rd;
  output [31:0] data_rd;
  input [19:0] addr_wr;
  input [31:0] data_wr;
  input clk, wr_ena;
  wire   wr_0, wr_1, n1, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22,
         SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24,
         SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26,
         SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28,
         SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30,
         SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32,
         SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34,
         SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36,
         SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38,
         SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40;
  wire   [11:0] data_rd_1;
  wire   [11:0] data_rd_0;

  mem_32_512_3 mem_0 ( .clk(clk), .addr_rd(addr_rd[8:0]), .wr_ena(wr_0), 
        .data_rd({SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, 
        SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, 
        SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, 
        SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10, 
        SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12, 
        SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14, 
        SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16, 
        SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18, 
        SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20, data_rd_0}), 
        .addr_wr(addr_wr[8:0]), .data_wr(data_wr) );
  mem_32_512_2 mem_1 ( .clk(clk), .addr_rd(addr_rd[8:0]), .wr_ena(wr_1), 
        .data_rd({SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22, 
        SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24, 
        SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26, 
        SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28, 
        SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30, 
        SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32, 
        SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34, 
        SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36, 
        SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38, 
        SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40, data_rd_1}), 
        .addr_wr(addr_wr[8:0]), .data_wr(data_wr) );
  NOR2X0 U1 ( .IN1(addr_wr[9]), .IN2(n1), .QN(wr_0) );
  AND2X1 U2 ( .IN1(addr_wr[9]), .IN2(wr_ena), .Q(wr_1) );
  MUX21X1 U3 ( .IN1(data_rd_0[0]), .IN2(data_rd_1[0]), .S(addr_rd[9]), .Q(
        data_rd[0]) );
  MUX21X1 U4 ( .IN1(data_rd_0[10]), .IN2(data_rd_1[10]), .S(addr_rd[9]), .Q(
        data_rd[10]) );
  MUX21X1 U5 ( .IN1(data_rd_0[11]), .IN2(data_rd_1[11]), .S(addr_rd[9]), .Q(
        data_rd[11]) );
  MUX21X1 U6 ( .IN1(data_rd_0[1]), .IN2(data_rd_1[1]), .S(addr_rd[9]), .Q(
        data_rd[1]) );
  MUX21X1 U7 ( .IN1(data_rd_0[2]), .IN2(data_rd_1[2]), .S(addr_rd[9]), .Q(
        data_rd[2]) );
  MUX21X1 U8 ( .IN1(data_rd_0[3]), .IN2(data_rd_1[3]), .S(addr_rd[9]), .Q(
        data_rd[3]) );
  MUX21X1 U9 ( .IN1(data_rd_0[4]), .IN2(data_rd_1[4]), .S(addr_rd[9]), .Q(
        data_rd[4]) );
  MUX21X1 U10 ( .IN1(data_rd_0[5]), .IN2(data_rd_1[5]), .S(addr_rd[9]), .Q(
        data_rd[5]) );
  MUX21X1 U11 ( .IN1(data_rd_0[6]), .IN2(data_rd_1[6]), .S(addr_rd[9]), .Q(
        data_rd[6]) );
  MUX21X1 U12 ( .IN1(data_rd_0[7]), .IN2(data_rd_1[7]), .S(addr_rd[9]), .Q(
        data_rd[7]) );
  MUX21X1 U13 ( .IN1(data_rd_0[8]), .IN2(data_rd_1[8]), .S(addr_rd[9]), .Q(
        data_rd[8]) );
  MUX21X1 U14 ( .IN1(data_rd_0[9]), .IN2(data_rd_1[9]), .S(addr_rd[9]), .Q(
        data_rd[9]) );
  INVX0 U15 ( .INP(wr_ena), .ZN(n1) );
endmodule


module mem_32_512_1 ( clk, addr_rd, wr_ena, data_rd, addr_wr, data_wr );
  input [8:0] addr_rd;
  output [31:0] data_rd;
  input [8:0] addr_wr;
  input [31:0] data_wr;
  input clk, wr_ena;


  SRAM32x512_1rw SRAM_HM_01 ( .I({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .O(data_rd), .A(addr_rd), .CE(1'b0), .CSB(1'b0), .WEB(1'b0), 
        .OEB(1'b0) );
endmodule


module mem_mfcc ( clk, addr, wr_ena, data );
  input [19:0] addr;
  output [31:0] data;
  input clk, wr_ena;


  mem_32_512_1 mem_0 ( .clk(clk), .addr_rd(addr[8:0]), .wr_ena(1'b0), 
        .data_rd(data), .addr_wr({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .data_wr({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
endmodule


module input_mac_controller ( clk, rst_n, is_odd_layer, is_first_layer, 
        ena_mac, ena_mac_wait, ena_mul_add, ena_mac_delay, w_addr, 
        input_or_int_mem_addr );
  output [19:0] w_addr;
  output [19:0] input_or_int_mem_addr;
  input clk, rst_n, is_odd_layer, is_first_layer, ena_mac, ena_mac_wait;
  output ena_mul_add, ena_mac_delay;
  wire   N19, N20, N21, N22, ena_rd_input_mac, N23, N142, N143, N144, N145,
         N146, n1, n2, n3, n4, n10, n13, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n5, n6, n7, n8, n9, n11, n12, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161;
  wire   [3:0] counter_rd_input_mac;
  wire   [9:0] addr_mem_back;
  wire   [9:0] addr_mem_front;
  wire   [3:0] counter_mul_add;

  DFFARX1 counter_rd_input_mac_reg_0_ ( .D(N19), .CLK(clk), .RSTB(rst_n), .Q(
        counter_rd_input_mac[0]) );
  DFFARX1 counter_rd_input_mac_reg_2_ ( .D(N21), .CLK(clk), .RSTB(rst_n), .Q(
        counter_rd_input_mac[2]), .QN(n34) );
  DFFARX1 counter_rd_input_mac_reg_3_ ( .D(N22), .CLK(clk), .RSTB(rst_n), .Q(
        counter_rd_input_mac[3]), .QN(n18) );
  DFFARX1 counter_rd_input_mac_reg_1_ ( .D(N20), .CLK(clk), .RSTB(rst_n), .Q(
        n8) );
  DFFARX1 ena_rd_input_mac_reg ( .D(N23), .CLK(clk), .RSTB(rst_n), .Q(
        ena_rd_input_mac), .QN(n7) );
  DFFARX1 w_addr_reg_19_ ( .D(n75), .CLK(clk), .RSTB(rst_n), .Q(w_addr[19]) );
  DFFARX1 w_addr_reg_18_ ( .D(n76), .CLK(clk), .RSTB(rst_n), .Q(w_addr[18]), 
        .QN(n9) );
  DFFARX1 w_addr_reg_17_ ( .D(n77), .CLK(clk), .RSTB(rst_n), .Q(w_addr[17]) );
  DFFARX1 w_addr_reg_16_ ( .D(n78), .CLK(clk), .RSTB(rst_n), .Q(w_addr[16]), 
        .QN(n17) );
  DFFARX1 w_addr_reg_15_ ( .D(n79), .CLK(clk), .RSTB(rst_n), .Q(w_addr[15]) );
  DFFARX1 w_addr_reg_14_ ( .D(n80), .CLK(clk), .RSTB(rst_n), .Q(w_addr[14]), 
        .QN(n16) );
  DFFARX1 w_addr_reg_13_ ( .D(n81), .CLK(clk), .RSTB(rst_n), .Q(w_addr[13]) );
  DFFARX1 w_addr_reg_12_ ( .D(n82), .CLK(clk), .RSTB(rst_n), .Q(w_addr[12]), 
        .QN(n15) );
  DFFARX1 w_addr_reg_11_ ( .D(n83), .CLK(clk), .RSTB(rst_n), .Q(w_addr[11]) );
  DFFARX1 w_addr_reg_10_ ( .D(n84), .CLK(clk), .RSTB(rst_n), .Q(w_addr[10]), 
        .QN(n14) );
  DFFARX1 w_addr_reg_9_ ( .D(n85), .CLK(clk), .RSTB(rst_n), .Q(w_addr[9]) );
  DFFARX1 w_addr_reg_8_ ( .D(n86), .CLK(clk), .RSTB(rst_n), .Q(w_addr[8]), 
        .QN(n12) );
  DFFARX1 w_addr_reg_7_ ( .D(n87), .CLK(clk), .RSTB(rst_n), .Q(w_addr[7]) );
  DFFARX1 w_addr_reg_6_ ( .D(n88), .CLK(clk), .RSTB(rst_n), .Q(w_addr[6]), 
        .QN(n11) );
  DFFARX1 w_addr_reg_5_ ( .D(n89), .CLK(clk), .RSTB(rst_n), .Q(w_addr[5]) );
  DFFARX1 w_addr_reg_4_ ( .D(n90), .CLK(clk), .RSTB(rst_n), .Q(w_addr[4]), 
        .QN(n30) );
  DFFARX1 w_addr_reg_3_ ( .D(n91), .CLK(clk), .RSTB(rst_n), .Q(w_addr[3]), 
        .QN(n22) );
  DFFARX1 w_addr_reg_2_ ( .D(n92), .CLK(clk), .RSTB(rst_n), .Q(w_addr[2]), 
        .QN(n32) );
  DFFARX1 w_addr_reg_1_ ( .D(n93), .CLK(clk), .RSTB(rst_n), .Q(w_addr[1]), 
        .QN(n23) );
  DFFARX1 w_addr_reg_0_ ( .D(n94), .CLK(clk), .RSTB(rst_n), .Q(w_addr[0]) );
  DFFASX1 addr_mem_back_reg_9_ ( .D(n65), .CLK(clk), .SETB(rst_n), .Q(
        addr_mem_back[9]), .QN(n33) );
  DFFARX1 addr_mem_back_reg_8_ ( .D(n66), .CLK(clk), .RSTB(rst_n), .Q(
        addr_mem_back[8]), .QN(n29) );
  DFFARX1 addr_mem_back_reg_7_ ( .D(n67), .CLK(clk), .RSTB(rst_n), .Q(
        addr_mem_back[7]) );
  DFFARX1 addr_mem_back_reg_6_ ( .D(n68), .CLK(clk), .RSTB(rst_n), .Q(
        addr_mem_back[6]), .QN(n25) );
  DFFARX1 addr_mem_back_reg_5_ ( .D(n69), .CLK(clk), .RSTB(rst_n), .Q(
        addr_mem_back[5]) );
  DFFARX1 addr_mem_back_reg_4_ ( .D(n70), .CLK(clk), .RSTB(rst_n), .Q(
        addr_mem_back[4]), .QN(n24) );
  DFFARX1 addr_mem_back_reg_3_ ( .D(n71), .CLK(clk), .RSTB(rst_n), .Q(
        addr_mem_back[3]) );
  DFFARX1 addr_mem_back_reg_2_ ( .D(n72), .CLK(clk), .RSTB(rst_n), .Q(
        addr_mem_back[2]) );
  DFFARX1 addr_mem_back_reg_1_ ( .D(n73), .CLK(clk), .RSTB(rst_n), .Q(
        addr_mem_back[1]) );
  DFFARX1 addr_mem_back_reg_0_ ( .D(n74), .CLK(clk), .RSTB(rst_n), .Q(
        addr_mem_back[0]), .QN(n19) );
  DFFARX1 addr_mem_front_reg_9_ ( .D(n45), .CLK(clk), .RSTB(rst_n), .Q(
        addr_mem_front[9]) );
  DFFARX1 addr_mem_front_reg_8_ ( .D(n46), .CLK(clk), .RSTB(rst_n), .Q(
        addr_mem_front[8]), .QN(n28) );
  DFFARX1 addr_mem_front_reg_7_ ( .D(n47), .CLK(clk), .RSTB(rst_n), .Q(
        addr_mem_front[7]) );
  DFFARX1 addr_mem_front_reg_6_ ( .D(n48), .CLK(clk), .RSTB(rst_n), .Q(
        addr_mem_front[6]), .QN(n27) );
  DFFARX1 addr_mem_front_reg_5_ ( .D(n49), .CLK(clk), .RSTB(rst_n), .Q(
        addr_mem_front[5]) );
  DFFARX1 addr_mem_front_reg_4_ ( .D(n50), .CLK(clk), .RSTB(rst_n), .Q(
        addr_mem_front[4]), .QN(n26) );
  DFFARX1 addr_mem_front_reg_3_ ( .D(n51), .CLK(clk), .RSTB(rst_n), .Q(
        addr_mem_front[3]) );
  DFFARX1 addr_mem_front_reg_2_ ( .D(n52), .CLK(clk), .RSTB(rst_n), .Q(
        addr_mem_front[2]) );
  DFFARX1 addr_mem_front_reg_1_ ( .D(n53), .CLK(clk), .RSTB(rst_n), .Q(
        addr_mem_front[1]) );
  DFFARX1 addr_mem_front_reg_0_ ( .D(n54), .CLK(clk), .RSTB(rst_n), .Q(
        addr_mem_front[0]), .QN(n20) );
  DFFASX1 ena_mac_w1_reg ( .D(n13), .CLK(clk), .SETB(rst_n), .Q(n4) );
  DFFASX1 ena_mac_w2_reg ( .D(n4), .CLK(clk), .SETB(rst_n), .Q(n3) );
  DFFASX1 ena_mac_w3_reg ( .D(n3), .CLK(clk), .SETB(rst_n), .Q(n2) );
  DFFASX1 ena_mac_w4_reg ( .D(n2), .CLK(clk), .SETB(rst_n), .Q(n1) );
  DFFASX1 ena_mac_delay_reg ( .D(n1), .CLK(clk), .SETB(rst_n), .QN(
        ena_mac_delay) );
  DFFARX1 counter_mul_add_reg_0_ ( .D(N142), .CLK(clk), .RSTB(rst_n), .Q(
        counter_mul_add[0]), .QN(n5) );
  DFFARX1 counter_mul_add_reg_2_ ( .D(N144), .CLK(clk), .RSTB(rst_n), .Q(
        counter_mul_add[2]), .QN(n6) );
  DFFARX1 counter_mul_add_reg_3_ ( .D(N145), .CLK(clk), .RSTB(rst_n), .Q(
        counter_mul_add[3]), .QN(n21) );
  DFFARX1 counter_mul_add_reg_1_ ( .D(N143), .CLK(clk), .RSTB(rst_n), .Q(n31), 
        .QN(n10) );
  DFFARX1 ena_mul_add_reg ( .D(N146), .CLK(clk), .RSTB(rst_n), .Q(ena_mul_add)
         );
  NAND2X0 U3 ( .IN1(counter_mul_add[2]), .IN2(n39), .QN(n41) );
  NAND2X0 U4 ( .IN1(n160), .IN2(n20), .QN(n135) );
  NAND2X0 U5 ( .IN1(n159), .IN2(n135), .QN(n138) );
  NAND2X0 U6 ( .IN1(n160), .IN2(n19), .QN(n113) );
  NAND2X0 U7 ( .IN1(n159), .IN2(n113), .QN(n116) );
  NAND2X0 U8 ( .IN1(n7), .IN2(ena_mac), .QN(n159) );
  NAND2X0 U9 ( .IN1(n160), .IN2(w_addr[0]), .QN(n62) );
  NAND2X0 U10 ( .IN1(w_addr[5]), .IN2(n98), .QN(n99) );
  NAND2X0 U11 ( .IN1(n100), .IN2(w_addr[7]), .QN(n101) );
  NAND2X0 U12 ( .IN1(n102), .IN2(w_addr[9]), .QN(n103) );
  NAND2X0 U13 ( .IN1(n104), .IN2(w_addr[11]), .QN(n105) );
  NAND2X0 U14 ( .IN1(n106), .IN2(w_addr[13]), .QN(n107) );
  NAND2X0 U15 ( .IN1(n108), .IN2(w_addr[15]), .QN(n109) );
  NAND2X0 U16 ( .IN1(n110), .IN2(w_addr[17]), .QN(n111) );
  NAND2X0 U17 ( .IN1(n43), .IN2(ena_mac), .QN(n58) );
  NAND2X0 U18 ( .IN1(n41), .IN2(n40), .QN(n36) );
  NAND2X0 U19 ( .IN1(addr_mem_front[1]), .IN2(addr_mem_front[0]), .QN(n136) );
  NAND2X0 U20 ( .IN1(addr_mem_back[1]), .IN2(addr_mem_back[0]), .QN(n114) );
  NAND2X0 U21 ( .IN1(ena_mac), .IN2(n133), .QN(n65) );
  NAND2X0 U22 ( .IN1(n160), .IN2(n96), .QN(n64) );
  NAND2X0 U23 ( .IN1(counter_rd_input_mac[2]), .IN2(n55), .QN(n56) );
  NAND2X0 U24 ( .IN1(ena_mac), .IN2(ena_rd_input_mac), .QN(n161) );
  NOR2X0 U25 ( .IN1(is_first_layer), .IN2(n60), .QN(n61) );
  INVX0 U26 ( .INP(n161), .ZN(n160) );
  NOR2X0 U27 ( .IN1(n35), .IN2(n36), .QN(N144) );
  NOR2X0 U28 ( .IN1(n39), .IN2(counter_mul_add[2]), .QN(n35) );
  NOR2X0 U29 ( .IN1(ena_mac_wait), .IN2(ena_mac_delay), .QN(n37) );
  NOR2X0 U30 ( .IN1(n37), .IN2(counter_mul_add[0]), .QN(N142) );
  NAND4X0 U31 ( .IN1(counter_mul_add[3]), .IN2(counter_mul_add[0]), .IN3(n10), 
        .IN4(n6), .QN(n38) );
  OA21X1 U32 ( .IN1(ena_mac_wait), .IN2(ena_mac_delay), .IN3(n38), .Q(n40) );
  OA221X1 U33 ( .IN1(counter_mul_add[0]), .IN2(n31), .IN3(n5), .IN4(n10), 
        .IN5(n40), .Q(N143) );
  NOR2X0 U34 ( .IN1(n10), .IN2(n5), .QN(n39) );
  INVX0 U35 ( .INP(n41), .ZN(n42) );
  OA221X1 U36 ( .IN1(counter_mul_add[3]), .IN2(n42), .IN3(n21), .IN4(n41), 
        .IN5(n40), .Q(N145) );
  AND4X1 U37 ( .IN1(n10), .IN2(N142), .IN3(n21), .IN4(n6), .Q(N146) );
  INVX0 U38 ( .INP(ena_mac), .ZN(n13) );
  NOR2X0 U39 ( .IN1(counter_rd_input_mac[0]), .IN2(n13), .QN(N19) );
  NOR2X0 U40 ( .IN1(counter_rd_input_mac[2]), .IN2(n8), .QN(n59) );
  NAND3X0 U41 ( .IN1(n59), .IN2(counter_rd_input_mac[3]), .IN3(
        counter_rd_input_mac[0]), .QN(n43) );
  AND2X1 U42 ( .IN1(n8), .IN2(counter_rd_input_mac[0]), .Q(n55) );
  NOR2X0 U43 ( .IN1(n58), .IN2(n55), .QN(n44) );
  OA21X1 U44 ( .IN1(counter_rd_input_mac[0]), .IN2(n8), .IN3(n44), .Q(N20) );
  OA222X1 U45 ( .IN1(counter_rd_input_mac[2]), .IN2(ena_mac), .IN3(
        counter_rd_input_mac[2]), .IN4(n55), .IN5(n44), .IN6(n34), .Q(N21) );
  MUX21X1 U46 ( .IN1(counter_rd_input_mac[3]), .IN2(n18), .S(n56), .Q(n57) );
  NOR2X0 U47 ( .IN1(n58), .IN2(n57), .QN(N22) );
  AND3X1 U48 ( .IN1(N19), .IN2(n59), .IN3(n18), .Q(N23) );
  INVX0 U49 ( .INP(is_odd_layer), .ZN(n60) );
  MUX21X1 U50 ( .IN1(addr_mem_front[0]), .IN2(addr_mem_back[0]), .S(n61), .Q(
        input_or_int_mem_addr[0]) );
  MUX21X1 U51 ( .IN1(addr_mem_front[1]), .IN2(addr_mem_back[1]), .S(n61), .Q(
        input_or_int_mem_addr[1]) );
  MUX21X1 U52 ( .IN1(addr_mem_front[2]), .IN2(addr_mem_back[2]), .S(n61), .Q(
        input_or_int_mem_addr[2]) );
  MUX21X1 U53 ( .IN1(addr_mem_front[3]), .IN2(addr_mem_back[3]), .S(n61), .Q(
        input_or_int_mem_addr[3]) );
  MUX21X1 U54 ( .IN1(addr_mem_front[4]), .IN2(addr_mem_back[4]), .S(n61), .Q(
        input_or_int_mem_addr[4]) );
  MUX21X1 U55 ( .IN1(addr_mem_front[5]), .IN2(addr_mem_back[5]), .S(n61), .Q(
        input_or_int_mem_addr[5]) );
  MUX21X1 U56 ( .IN1(addr_mem_front[6]), .IN2(addr_mem_back[6]), .S(n61), .Q(
        input_or_int_mem_addr[6]) );
  MUX21X1 U57 ( .IN1(addr_mem_front[7]), .IN2(addr_mem_back[7]), .S(n61), .Q(
        input_or_int_mem_addr[7]) );
  MUX21X1 U58 ( .IN1(addr_mem_front[8]), .IN2(addr_mem_back[8]), .S(n61), .Q(
        input_or_int_mem_addr[8]) );
  MUX21X1 U59 ( .IN1(addr_mem_front[9]), .IN2(addr_mem_back[9]), .S(n61), .Q(
        input_or_int_mem_addr[9]) );
  OA21X1 U60 ( .IN1(n160), .IN2(w_addr[0]), .IN3(n62), .Q(n94) );
  MUX21X1 U61 ( .IN1(n23), .IN2(w_addr[1]), .S(n62), .Q(n93) );
  NAND3X0 U62 ( .IN1(n160), .IN2(w_addr[1]), .IN3(w_addr[0]), .QN(n63) );
  MUX21X1 U63 ( .IN1(n32), .IN2(w_addr[2]), .S(n63), .Q(n92) );
  AND3X1 U64 ( .IN1(w_addr[2]), .IN2(w_addr[1]), .IN3(w_addr[0]), .Q(n96) );
  MUX21X1 U65 ( .IN1(n22), .IN2(w_addr[3]), .S(n64), .Q(n91) );
  NAND3X0 U66 ( .IN1(n160), .IN2(n96), .IN3(w_addr[3]), .QN(n95) );
  MUX21X1 U67 ( .IN1(n30), .IN2(w_addr[4]), .S(n95), .Q(n90) );
  NAND3X0 U68 ( .IN1(n96), .IN2(w_addr[4]), .IN3(w_addr[3]), .QN(n97) );
  NOR2X0 U69 ( .IN1(n161), .IN2(n97), .QN(n98) );
  OA21X1 U70 ( .IN1(w_addr[5]), .IN2(n98), .IN3(n99), .Q(n89) );
  MUX21X1 U71 ( .IN1(n11), .IN2(w_addr[6]), .S(n99), .Q(n88) );
  NOR2X0 U72 ( .IN1(n11), .IN2(n99), .QN(n100) );
  OA21X1 U73 ( .IN1(n100), .IN2(w_addr[7]), .IN3(n101), .Q(n87) );
  MUX21X1 U74 ( .IN1(n12), .IN2(w_addr[8]), .S(n101), .Q(n86) );
  NOR2X0 U75 ( .IN1(n12), .IN2(n101), .QN(n102) );
  OA21X1 U76 ( .IN1(n102), .IN2(w_addr[9]), .IN3(n103), .Q(n85) );
  MUX21X1 U77 ( .IN1(n14), .IN2(w_addr[10]), .S(n103), .Q(n84) );
  NOR2X0 U78 ( .IN1(n103), .IN2(n14), .QN(n104) );
  OA21X1 U79 ( .IN1(n104), .IN2(w_addr[11]), .IN3(n105), .Q(n83) );
  MUX21X1 U80 ( .IN1(n15), .IN2(w_addr[12]), .S(n105), .Q(n82) );
  NOR2X0 U81 ( .IN1(n105), .IN2(n15), .QN(n106) );
  OA21X1 U82 ( .IN1(n106), .IN2(w_addr[13]), .IN3(n107), .Q(n81) );
  MUX21X1 U83 ( .IN1(n16), .IN2(w_addr[14]), .S(n107), .Q(n80) );
  NOR2X0 U84 ( .IN1(n107), .IN2(n16), .QN(n108) );
  OA21X1 U85 ( .IN1(n108), .IN2(w_addr[15]), .IN3(n109), .Q(n79) );
  MUX21X1 U86 ( .IN1(n17), .IN2(w_addr[16]), .S(n109), .Q(n78) );
  NOR2X0 U87 ( .IN1(n109), .IN2(n17), .QN(n110) );
  OA21X1 U88 ( .IN1(n110), .IN2(w_addr[17]), .IN3(n111), .Q(n77) );
  MUX21X1 U89 ( .IN1(n9), .IN2(w_addr[18]), .S(n111), .Q(n76) );
  OR2X1 U90 ( .IN1(n111), .IN2(n9), .Q(n112) );
  XNOR2X1 U91 ( .IN1(w_addr[19]), .IN2(n112), .Q(n75) );
  OAI21X1 U92 ( .IN1(n19), .IN2(n159), .IN3(n113), .QN(n74) );
  NOR2X0 U93 ( .IN1(addr_mem_back[1]), .IN2(n161), .QN(n117) );
  AO22X1 U94 ( .IN1(addr_mem_back[1]), .IN2(n116), .IN3(addr_mem_back[0]), 
        .IN4(n117), .Q(n73) );
  NOR3X0 U95 ( .IN1(addr_mem_back[2]), .IN2(n114), .IN3(n161), .QN(n115) );
  AO221X1 U96 ( .IN1(addr_mem_back[2]), .IN2(n117), .IN3(addr_mem_back[2]), 
        .IN4(n116), .IN5(n115), .Q(n72) );
  NAND3X0 U97 ( .IN1(addr_mem_back[1]), .IN2(addr_mem_back[0]), .IN3(
        addr_mem_back[2]), .QN(n118) );
  INVX0 U98 ( .INP(n118), .ZN(n122) );
  NOR2X0 U99 ( .IN1(addr_mem_back[3]), .IN2(n161), .QN(n121) );
  OA21X1 U100 ( .IN1(n7), .IN2(n118), .IN3(ena_mac), .Q(n120) );
  AO22X1 U101 ( .IN1(n122), .IN2(n121), .IN3(addr_mem_back[3]), .IN4(n120), 
        .Q(n71) );
  AND3X1 U102 ( .IN1(n160), .IN2(n122), .IN3(addr_mem_back[3]), .Q(n119) );
  AO222X1 U103 ( .IN1(addr_mem_back[4]), .IN2(n121), .IN3(addr_mem_back[4]), 
        .IN4(n120), .IN5(n119), .IN6(n24), .Q(n70) );
  NAND3X0 U104 ( .IN1(n122), .IN2(addr_mem_back[4]), .IN3(addr_mem_back[3]), 
        .QN(n123) );
  INVX0 U105 ( .INP(n123), .ZN(n127) );
  NOR2X0 U106 ( .IN1(addr_mem_back[5]), .IN2(n161), .QN(n126) );
  OA21X1 U107 ( .IN1(n7), .IN2(n123), .IN3(ena_mac), .Q(n125) );
  AO22X1 U108 ( .IN1(n127), .IN2(n126), .IN3(addr_mem_back[5]), .IN4(n125), 
        .Q(n69) );
  AND3X1 U109 ( .IN1(n160), .IN2(n127), .IN3(addr_mem_back[5]), .Q(n124) );
  AO222X1 U110 ( .IN1(addr_mem_back[6]), .IN2(n126), .IN3(addr_mem_back[6]), 
        .IN4(n125), .IN5(n124), .IN6(n25), .Q(n68) );
  NAND3X0 U111 ( .IN1(n127), .IN2(addr_mem_back[6]), .IN3(addr_mem_back[5]), 
        .QN(n128) );
  INVX0 U112 ( .INP(n128), .ZN(n134) );
  NOR2X0 U113 ( .IN1(addr_mem_back[7]), .IN2(n161), .QN(n131) );
  OA21X1 U114 ( .IN1(n7), .IN2(n128), .IN3(ena_mac), .Q(n130) );
  AO22X1 U115 ( .IN1(n134), .IN2(n131), .IN3(addr_mem_back[7]), .IN4(n130), 
        .Q(n67) );
  AND3X1 U116 ( .IN1(n160), .IN2(n134), .IN3(addr_mem_back[7]), .Q(n129) );
  AO222X1 U117 ( .IN1(addr_mem_back[8]), .IN2(n131), .IN3(addr_mem_back[8]), 
        .IN4(n130), .IN5(n129), .IN6(n29), .Q(n66) );
  NAND4X0 U118 ( .IN1(n134), .IN2(addr_mem_back[8]), .IN3(addr_mem_back[7]), 
        .IN4(n159), .QN(n132) );
  MUX21X1 U119 ( .IN1(addr_mem_back[9]), .IN2(n33), .S(n132), .Q(n133) );
  OAI21X1 U120 ( .IN1(n20), .IN2(n159), .IN3(n135), .QN(n54) );
  NOR2X0 U121 ( .IN1(addr_mem_front[1]), .IN2(n161), .QN(n139) );
  AO22X1 U122 ( .IN1(addr_mem_front[1]), .IN2(n138), .IN3(addr_mem_front[0]), 
        .IN4(n139), .Q(n53) );
  NOR3X0 U123 ( .IN1(addr_mem_front[2]), .IN2(n136), .IN3(n161), .QN(n137) );
  AO221X1 U124 ( .IN1(addr_mem_front[2]), .IN2(n139), .IN3(addr_mem_front[2]), 
        .IN4(n138), .IN5(n137), .Q(n52) );
  NAND3X0 U125 ( .IN1(addr_mem_front[1]), .IN2(addr_mem_front[0]), .IN3(
        addr_mem_front[2]), .QN(n140) );
  INVX0 U126 ( .INP(n140), .ZN(n144) );
  NOR2X0 U127 ( .IN1(addr_mem_front[3]), .IN2(n161), .QN(n143) );
  OA21X1 U128 ( .IN1(n7), .IN2(n140), .IN3(ena_mac), .Q(n142) );
  AO22X1 U129 ( .IN1(n144), .IN2(n143), .IN3(addr_mem_front[3]), .IN4(n142), 
        .Q(n51) );
  AND3X1 U130 ( .IN1(n160), .IN2(n144), .IN3(addr_mem_front[3]), .Q(n141) );
  AO222X1 U131 ( .IN1(addr_mem_front[4]), .IN2(n143), .IN3(addr_mem_front[4]), 
        .IN4(n142), .IN5(n141), .IN6(n26), .Q(n50) );
  NAND3X0 U132 ( .IN1(n144), .IN2(addr_mem_front[4]), .IN3(addr_mem_front[3]), 
        .QN(n145) );
  INVX0 U133 ( .INP(n145), .ZN(n149) );
  NOR2X0 U134 ( .IN1(addr_mem_front[5]), .IN2(n161), .QN(n148) );
  OA21X1 U135 ( .IN1(n7), .IN2(n145), .IN3(ena_mac), .Q(n147) );
  AO22X1 U136 ( .IN1(n149), .IN2(n148), .IN3(addr_mem_front[5]), .IN4(n147), 
        .Q(n49) );
  AND3X1 U137 ( .IN1(n160), .IN2(n149), .IN3(addr_mem_front[5]), .Q(n146) );
  AO222X1 U138 ( .IN1(addr_mem_front[6]), .IN2(n148), .IN3(addr_mem_front[6]), 
        .IN4(n147), .IN5(n146), .IN6(n27), .Q(n48) );
  NAND3X0 U139 ( .IN1(n149), .IN2(addr_mem_front[6]), .IN3(addr_mem_front[5]), 
        .QN(n150) );
  INVX0 U140 ( .INP(n150), .ZN(n154) );
  NOR2X0 U141 ( .IN1(addr_mem_front[7]), .IN2(n161), .QN(n153) );
  OA21X1 U142 ( .IN1(n7), .IN2(n150), .IN3(ena_mac), .Q(n152) );
  AO22X1 U143 ( .IN1(n154), .IN2(n153), .IN3(addr_mem_front[7]), .IN4(n152), 
        .Q(n47) );
  AND3X1 U144 ( .IN1(n160), .IN2(n154), .IN3(addr_mem_front[7]), .Q(n151) );
  AO222X1 U145 ( .IN1(addr_mem_front[8]), .IN2(n153), .IN3(addr_mem_front[8]), 
        .IN4(n152), .IN5(n151), .IN6(n28), .Q(n46) );
  NAND3X0 U146 ( .IN1(n154), .IN2(addr_mem_front[8]), .IN3(addr_mem_front[7]), 
        .QN(n155) );
  INVX0 U147 ( .INP(n155), .ZN(n158) );
  NOR2X0 U148 ( .IN1(addr_mem_front[9]), .IN2(n161), .QN(n157) );
  OA21X1 U149 ( .IN1(n7), .IN2(n155), .IN3(ena_mac), .Q(n156) );
  AO22X1 U150 ( .IN1(n158), .IN2(n157), .IN3(addr_mem_front[9]), .IN4(n156), 
        .Q(n45) );
endmodule


module booth27_0 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93;

  NAND2X0 U3 ( .IN1(n27), .IN2(n26), .QN(n29) );
  NAND2X0 U4 ( .IN1(n32), .IN2(n31), .QN(n34) );
  NAND2X0 U5 ( .IN1(n37), .IN2(n36), .QN(n39) );
  NAND2X0 U6 ( .IN1(n42), .IN2(n41), .QN(n47) );
  NAND2X0 U7 ( .IN1(n78), .IN2(n12), .QN(n82) );
  NAND2X0 U8 ( .IN1(n22), .IN2(n21), .QN(n24) );
  NAND2X0 U9 ( .IN1(in1[2]), .IN2(n47), .QN(n44) );
  NAND2X0 U10 ( .IN1(n52), .IN2(n6), .QN(n55) );
  NAND2X0 U11 ( .IN1(in1[2]), .IN2(n55), .QN(n51) );
  NAND2X0 U12 ( .IN1(n60), .IN2(n8), .QN(n63) );
  NAND2X0 U13 ( .IN1(in1[2]), .IN2(n63), .QN(n59) );
  NAND2X0 U14 ( .IN1(n68), .IN2(n10), .QN(n71) );
  NAND2X0 U15 ( .IN1(in1[2]), .IN2(n71), .QN(n67) );
  NAND2X0 U16 ( .IN1(in1[2]), .IN2(n82), .QN(n77) );
  NAND2X0 U17 ( .IN1(in2[21]), .IN2(n82), .QN(n83) );
  NAND2X0 U18 ( .IN1(n75), .IN2(in1[2]), .QN(n86) );
  NAND2X0 U19 ( .IN1(n3), .IN2(n4), .QN(n17) );
  NAND2X0 U20 ( .IN1(n18), .IN2(n17), .QN(out1[2]) );
  INVX0 U21 ( .INP(n86), .ZN(n89) );
  NAND2X0 U22 ( .IN1(in2[1]), .IN2(in2[0]), .QN(n4) );
  NOR2X0 U23 ( .IN1(n16), .IN2(n86), .QN(n3) );
  NOR2X0 U24 ( .IN1(in1[2]), .IN2(n75), .QN(n90) );
  NOR2X0 U25 ( .IN1(n75), .IN2(n72), .QN(n92) );
  NBUFFX2 U26 ( .INP(in1[2]), .Z(out1[26]) );
  NBUFFX2 U27 ( .INP(in1[2]), .Z(out1[25]) );
  INVX0 U28 ( .INP(in2[13]), .ZN(n5) );
  INVX0 U29 ( .INP(in2[14]), .ZN(n6) );
  INVX0 U30 ( .INP(in2[15]), .ZN(n7) );
  INVX0 U31 ( .INP(in2[16]), .ZN(n8) );
  INVX0 U32 ( .INP(in2[17]), .ZN(n9) );
  INVX0 U33 ( .INP(in2[18]), .ZN(n10) );
  INVX0 U34 ( .INP(in2[19]), .ZN(n11) );
  INVX0 U35 ( .INP(in2[20]), .ZN(n12) );
  INVX0 U36 ( .INP(in2[21]), .ZN(n13) );
  INVX0 U37 ( .INP(in2[22]), .ZN(n14) );
  INVX0 U38 ( .INP(in1[1]), .ZN(n75) );
  INVX0 U39 ( .INP(in1[2]), .ZN(n72) );
  NOR2X0 U40 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n16) );
  INVX0 U41 ( .INP(in2[2]), .ZN(n15) );
  OR3X1 U42 ( .IN1(in2[2]), .IN2(in2[0]), .IN3(in2[1]), .Q(n19) );
  OA21X1 U43 ( .IN1(n16), .IN2(n15), .IN3(n19), .Q(n20) );
  AOI22X1 U44 ( .IN1(in2[2]), .IN2(n90), .IN3(n92), .IN4(n20), .QN(n18) );
  NOR2X0 U45 ( .IN1(in2[3]), .IN2(n19), .QN(n22) );
  AOI21X1 U46 ( .IN1(in2[3]), .IN2(n19), .IN3(n22), .QN(n23) );
  AO222X1 U47 ( .IN1(in2[3]), .IN2(n90), .IN3(n92), .IN4(n23), .IN5(n89), 
        .IN6(n20), .Q(out1[3]) );
  INVX0 U48 ( .INP(in2[4]), .ZN(n21) );
  OA21X1 U49 ( .IN1(n22), .IN2(n21), .IN3(n24), .Q(n25) );
  AO222X1 U50 ( .IN1(in2[4]), .IN2(n90), .IN3(n92), .IN4(n25), .IN5(n89), 
        .IN6(n23), .Q(out1[4]) );
  NOR2X0 U51 ( .IN1(in2[5]), .IN2(n24), .QN(n27) );
  AOI21X1 U52 ( .IN1(in2[5]), .IN2(n24), .IN3(n27), .QN(n28) );
  AO222X1 U53 ( .IN1(in2[5]), .IN2(n90), .IN3(n92), .IN4(n28), .IN5(n89), 
        .IN6(n25), .Q(out1[5]) );
  INVX0 U54 ( .INP(in2[6]), .ZN(n26) );
  OA21X1 U55 ( .IN1(n27), .IN2(n26), .IN3(n29), .Q(n30) );
  AO222X1 U56 ( .IN1(in2[6]), .IN2(n90), .IN3(n92), .IN4(n30), .IN5(n89), 
        .IN6(n28), .Q(out1[6]) );
  NOR2X0 U57 ( .IN1(in2[7]), .IN2(n29), .QN(n32) );
  AOI21X1 U58 ( .IN1(in2[7]), .IN2(n29), .IN3(n32), .QN(n33) );
  AO222X1 U59 ( .IN1(in2[7]), .IN2(n90), .IN3(n92), .IN4(n33), .IN5(n89), 
        .IN6(n30), .Q(out1[7]) );
  INVX0 U60 ( .INP(in2[8]), .ZN(n31) );
  OA21X1 U61 ( .IN1(n32), .IN2(n31), .IN3(n34), .Q(n35) );
  AO222X1 U62 ( .IN1(in2[8]), .IN2(n90), .IN3(n92), .IN4(n35), .IN5(n89), 
        .IN6(n33), .Q(out1[8]) );
  NOR2X0 U63 ( .IN1(in2[9]), .IN2(n34), .QN(n37) );
  AOI21X1 U64 ( .IN1(in2[9]), .IN2(n34), .IN3(n37), .QN(n38) );
  AO222X1 U65 ( .IN1(in2[9]), .IN2(n90), .IN3(n92), .IN4(n38), .IN5(n89), 
        .IN6(n35), .Q(out1[9]) );
  INVX0 U66 ( .INP(in2[10]), .ZN(n36) );
  OA21X1 U67 ( .IN1(n37), .IN2(n36), .IN3(n39), .Q(n40) );
  AO222X1 U68 ( .IN1(in2[10]), .IN2(n90), .IN3(n92), .IN4(n40), .IN5(n89), 
        .IN6(n38), .Q(out1[10]) );
  NOR2X0 U69 ( .IN1(in2[11]), .IN2(n39), .QN(n42) );
  AOI21X1 U70 ( .IN1(in2[11]), .IN2(n39), .IN3(n42), .QN(n43) );
  AO222X1 U71 ( .IN1(in2[11]), .IN2(n90), .IN3(n92), .IN4(n43), .IN5(n89), 
        .IN6(n40), .Q(out1[11]) );
  INVX0 U72 ( .INP(in2[12]), .ZN(n41) );
  OA21X1 U73 ( .IN1(n42), .IN2(n41), .IN3(n47), .Q(n45) );
  AO222X1 U74 ( .IN1(in2[12]), .IN2(n90), .IN3(n92), .IN4(n45), .IN5(n89), 
        .IN6(n43), .Q(out1[12]) );
  MUX21X1 U75 ( .IN1(n5), .IN2(in2[13]), .S(n44), .Q(n46) );
  AO22X1 U76 ( .IN1(in1[1]), .IN2(n46), .IN3(n89), .IN4(n45), .Q(out1[13]) );
  NOR2X0 U77 ( .IN1(in2[13]), .IN2(n47), .QN(n52) );
  AO21X1 U78 ( .IN1(in2[13]), .IN2(n47), .IN3(n86), .Q(n50) );
  NOR2X0 U79 ( .IN1(n52), .IN2(n72), .QN(n48) );
  MUX21X1 U80 ( .IN1(n6), .IN2(in2[14]), .S(n48), .Q(n49) );
  OAI22X1 U81 ( .IN1(n52), .IN2(n50), .IN3(n75), .IN4(n49), .QN(out1[14]) );
  MUX21X1 U82 ( .IN1(n7), .IN2(in2[15]), .S(n51), .Q(n54) );
  OA21X1 U83 ( .IN1(n52), .IN2(n6), .IN3(n89), .Q(n53) );
  AO22X1 U84 ( .IN1(in1[1]), .IN2(n54), .IN3(n53), .IN4(n55), .Q(out1[15]) );
  NOR2X0 U85 ( .IN1(in2[15]), .IN2(n55), .QN(n60) );
  AO21X1 U86 ( .IN1(in2[15]), .IN2(n55), .IN3(n86), .Q(n58) );
  NOR2X0 U87 ( .IN1(n60), .IN2(n72), .QN(n56) );
  MUX21X1 U88 ( .IN1(n8), .IN2(in2[16]), .S(n56), .Q(n57) );
  OAI22X1 U89 ( .IN1(n60), .IN2(n58), .IN3(n75), .IN4(n57), .QN(out1[16]) );
  MUX21X1 U90 ( .IN1(n9), .IN2(in2[17]), .S(n59), .Q(n62) );
  OA21X1 U91 ( .IN1(n60), .IN2(n8), .IN3(n89), .Q(n61) );
  AO22X1 U92 ( .IN1(in1[1]), .IN2(n62), .IN3(n61), .IN4(n63), .Q(out1[17]) );
  NOR2X0 U93 ( .IN1(in2[17]), .IN2(n63), .QN(n68) );
  AO21X1 U94 ( .IN1(in2[17]), .IN2(n63), .IN3(n86), .Q(n66) );
  NOR2X0 U95 ( .IN1(n68), .IN2(n72), .QN(n64) );
  MUX21X1 U96 ( .IN1(n10), .IN2(in2[18]), .S(n64), .Q(n65) );
  OAI22X1 U97 ( .IN1(n68), .IN2(n66), .IN3(n75), .IN4(n65), .QN(out1[18]) );
  MUX21X1 U98 ( .IN1(n11), .IN2(in2[19]), .S(n67), .Q(n70) );
  OA21X1 U99 ( .IN1(n68), .IN2(n10), .IN3(n89), .Q(n69) );
  AO22X1 U100 ( .IN1(in1[1]), .IN2(n70), .IN3(n69), .IN4(n71), .Q(out1[19]) );
  NOR2X0 U101 ( .IN1(in2[19]), .IN2(n71), .QN(n78) );
  AO21X1 U102 ( .IN1(in2[19]), .IN2(n71), .IN3(n86), .Q(n76) );
  NOR2X0 U103 ( .IN1(n78), .IN2(n72), .QN(n73) );
  MUX21X1 U104 ( .IN1(n12), .IN2(in2[20]), .S(n73), .Q(n74) );
  OAI22X1 U105 ( .IN1(n78), .IN2(n76), .IN3(n75), .IN4(n74), .QN(out1[20]) );
  MUX21X1 U106 ( .IN1(n13), .IN2(in2[21]), .S(n77), .Q(n80) );
  MUX21X1 U107 ( .IN1(n12), .IN2(in2[20]), .S(n78), .Q(n79) );
  AO22X1 U108 ( .IN1(in1[1]), .IN2(n80), .IN3(n89), .IN4(n79), .Q(out1[21]) );
  INVX0 U109 ( .INP(n92), .ZN(n81) );
  OR2X1 U110 ( .IN1(n82), .IN2(in2[21]), .Q(n88) );
  NOR2X0 U111 ( .IN1(n81), .IN2(n88), .QN(n87) );
  NOR2X0 U112 ( .IN1(in2[22]), .IN2(n81), .QN(n84) );
  OA221X1 U113 ( .IN1(n84), .IN2(n89), .IN3(n84), .IN4(n83), .IN5(n88), .Q(n85) );
  AO221X1 U114 ( .IN1(in2[22]), .IN2(n87), .IN3(in2[22]), .IN4(n90), .IN5(n85), 
        .Q(out1[22]) );
  NOR2X0 U115 ( .IN1(n86), .IN2(n88), .QN(n93) );
  AO21X1 U116 ( .IN1(n89), .IN2(n88), .IN3(n87), .Q(n91) );
  AO221X1 U117 ( .IN1(in2[22]), .IN2(n93), .IN3(n14), .IN4(n91), .IN5(n90), 
        .Q(out1[23]) );
  AO21X1 U118 ( .IN1(n93), .IN2(n14), .IN3(n92), .Q(out1[24]) );
endmodule


module csa51squ_0 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n2, n3, n4, n5;

  NBUFFX2 U1 ( .INP(in3[31]), .Z(sumout[31]) );
  AND2X1 U2 ( .IN1(in2[2]), .IN2(in1[2]), .Q(cout[2]) );
  AND2X1 U3 ( .IN1(in2[3]), .IN2(in1[3]), .Q(cout[3]) );
  NOR2X0 U4 ( .IN1(in2[3]), .IN2(in1[3]), .QN(n2) );
  NOR2X0 U5 ( .IN1(n2), .IN2(cout[3]), .QN(sumout[3]) );
  AND2X1 U6 ( .IN1(in2[28]), .IN2(in3[28]), .Q(cout[28]) );
  NOR2X0 U7 ( .IN1(in2[28]), .IN2(in3[28]), .QN(n3) );
  NOR2X0 U8 ( .IN1(n3), .IN2(cout[28]), .QN(sumout[28]) );
  INVX0 U9 ( .INP(in3[29]), .ZN(n4) );
  NOR2X0 U10 ( .IN1(in2[28]), .IN2(n4), .QN(cout[29]) );
  MUX21X1 U11 ( .IN1(n4), .IN2(in3[29]), .S(in2[28]), .Q(sumout[29]) );
  INVX0 U12 ( .INP(in1[26]), .ZN(n5) );
  FADDX1 U13 ( .A(in1[10]), .B(in2[10]), .CI(in3[10]), .CO(cout[10]), .S(
        sumout[10]) );
  FADDX1 U14 ( .A(in1[11]), .B(in2[11]), .CI(in3[11]), .CO(cout[11]), .S(
        sumout[11]) );
  FADDX1 U15 ( .A(in1[12]), .B(in2[12]), .CI(in3[12]), .CO(cout[12]), .S(
        sumout[12]) );
  FADDX1 U16 ( .A(in1[13]), .B(in2[13]), .CI(in3[13]), .CO(cout[13]), .S(
        sumout[13]) );
  FADDX1 U17 ( .A(in1[14]), .B(in2[14]), .CI(in3[14]), .CO(cout[14]), .S(
        sumout[14]) );
  FADDX1 U18 ( .A(in1[15]), .B(in2[15]), .CI(in3[15]), .CO(cout[15]), .S(
        sumout[15]) );
  FADDX1 U19 ( .A(in1[16]), .B(in2[16]), .CI(in3[16]), .CO(cout[16]), .S(
        sumout[16]) );
  FADDX1 U20 ( .A(in1[17]), .B(in2[17]), .CI(in3[17]), .CO(cout[17]), .S(
        sumout[17]) );
  FADDX1 U21 ( .A(in1[18]), .B(in2[18]), .CI(in3[18]), .CO(cout[18]), .S(
        sumout[18]) );
  FADDX1 U22 ( .A(in1[19]), .B(in2[19]), .CI(in3[19]), .CO(cout[19]), .S(
        sumout[19]) );
  FADDX1 U23 ( .A(in1[20]), .B(in2[20]), .CI(in3[20]), .CO(cout[20]), .S(
        sumout[20]) );
  FADDX1 U24 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U25 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U26 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U27 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U28 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U29 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U30 ( .A(in2[27]), .B(in3[27]), .CI(n5), .CO(cout[27]), .S(sumout[27]) );
  FADDX1 U31 ( .A(in1[4]), .B(in2[4]), .CI(in3[4]), .CO(cout[4]), .S(sumout[4]) );
  FADDX1 U32 ( .A(in1[5]), .B(in2[5]), .CI(in3[5]), .CO(cout[5]), .S(sumout[5]) );
  FADDX1 U33 ( .A(in1[6]), .B(in2[6]), .CI(in3[6]), .CO(cout[6]), .S(sumout[6]) );
  FADDX1 U34 ( .A(in1[7]), .B(in2[7]), .CI(in3[7]), .CO(cout[7]), .S(sumout[7]) );
  FADDX1 U35 ( .A(in1[8]), .B(in2[8]), .CI(in3[8]), .CO(cout[8]), .S(sumout[8]) );
  FADDX1 U36 ( .A(in1[9]), .B(in2[9]), .CI(in3[9]), .CO(cout[9]), .S(sumout[9]) );
endmodule


module cla51squ_0 ( out, a, b );
  output [50:0] out;
  input [50:0] a;
  input [50:0] b;
  wire   intadd_0_CI, intadd_0_n24, intadd_0_n23, intadd_0_n22, intadd_0_n21,
         intadd_0_n20, intadd_0_n19, intadd_0_n18, intadd_0_n17, intadd_0_n16,
         intadd_0_n15, intadd_0_n14, intadd_0_n13, intadd_0_n12, intadd_0_n11,
         intadd_0_n10, intadd_0_n9, intadd_0_n8, intadd_0_n7, intadd_0_n6,
         intadd_0_n5, intadd_0_n4, intadd_0_n3, intadd_0_n2, intadd_0_n1, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14;

  FADDX1 intadd_0_U25 ( .A(b[23]), .B(a[23]), .CI(intadd_0_CI), .CO(
        intadd_0_n24), .S(out[23]) );
  FADDX1 intadd_0_U24 ( .A(b[24]), .B(a[24]), .CI(intadd_0_n24), .CO(
        intadd_0_n23), .S(out[24]) );
  FADDX1 intadd_0_U23 ( .A(b[25]), .B(a[25]), .CI(intadd_0_n23), .CO(
        intadd_0_n22), .S(out[25]) );
  FADDX1 intadd_0_U22 ( .A(b[26]), .B(a[26]), .CI(intadd_0_n22), .CO(
        intadd_0_n21), .S(out[26]) );
  FADDX1 intadd_0_U21 ( .A(b[27]), .B(a[27]), .CI(intadd_0_n21), .CO(
        intadd_0_n20), .S(out[27]) );
  FADDX1 intadd_0_U20 ( .A(b[28]), .B(a[28]), .CI(intadd_0_n20), .CO(
        intadd_0_n19), .S(out[28]) );
  FADDX1 intadd_0_U19 ( .A(b[29]), .B(a[29]), .CI(intadd_0_n19), .CO(
        intadd_0_n18), .S(out[29]) );
  FADDX1 intadd_0_U18 ( .A(b[30]), .B(a[30]), .CI(intadd_0_n18), .CO(
        intadd_0_n17), .S(out[30]) );
  FADDX1 intadd_0_U17 ( .A(b[31]), .B(a[31]), .CI(intadd_0_n17), .CO(
        intadd_0_n16), .S(out[31]) );
  FADDX1 intadd_0_U16 ( .A(b[32]), .B(a[32]), .CI(intadd_0_n16), .CO(
        intadd_0_n15), .S(out[32]) );
  FADDX1 intadd_0_U15 ( .A(b[33]), .B(a[33]), .CI(intadd_0_n15), .CO(
        intadd_0_n14), .S(out[33]) );
  FADDX1 intadd_0_U14 ( .A(b[34]), .B(a[34]), .CI(intadd_0_n14), .CO(
        intadd_0_n13), .S(out[34]) );
  FADDX1 intadd_0_U13 ( .A(b[35]), .B(a[35]), .CI(intadd_0_n13), .CO(
        intadd_0_n12), .S(out[35]) );
  FADDX1 intadd_0_U12 ( .A(b[36]), .B(a[36]), .CI(intadd_0_n12), .CO(
        intadd_0_n11), .S(out[36]) );
  FADDX1 intadd_0_U11 ( .A(b[37]), .B(a[37]), .CI(intadd_0_n11), .CO(
        intadd_0_n10), .S(out[37]) );
  FADDX1 intadd_0_U10 ( .A(b[38]), .B(a[38]), .CI(intadd_0_n10), .CO(
        intadd_0_n9), .S(out[38]) );
  FADDX1 intadd_0_U9 ( .A(b[39]), .B(a[39]), .CI(intadd_0_n9), .CO(intadd_0_n8), .S(out[39]) );
  FADDX1 intadd_0_U8 ( .A(b[40]), .B(a[40]), .CI(intadd_0_n8), .CO(intadd_0_n7), .S(out[40]) );
  FADDX1 intadd_0_U7 ( .A(b[41]), .B(a[41]), .CI(intadd_0_n7), .CO(intadd_0_n6), .S(out[41]) );
  FADDX1 intadd_0_U6 ( .A(b[42]), .B(a[42]), .CI(intadd_0_n6), .CO(intadd_0_n5), .S(out[42]) );
  FADDX1 intadd_0_U5 ( .A(b[43]), .B(a[43]), .CI(intadd_0_n5), .CO(intadd_0_n4), .S(out[43]) );
  FADDX1 intadd_0_U4 ( .A(b[44]), .B(a[44]), .CI(intadd_0_n4), .CO(intadd_0_n3), .S(out[44]) );
  FADDX1 intadd_0_U3 ( .A(b[45]), .B(a[45]), .CI(intadd_0_n3), .CO(intadd_0_n2), .S(out[45]) );
  FADDX1 intadd_0_U2 ( .A(b[46]), .B(a[46]), .CI(intadd_0_n2), .CO(intadd_0_n1), .S(out[46]) );
  OA21X1 U2 ( .IN1(b[9]), .IN2(a[9]), .IN3(a[8]), .Q(n1) );
  AO22X1 U3 ( .IN1(b[9]), .IN2(a[9]), .IN3(b[8]), .IN4(n1), .Q(n2) );
  AO222X1 U4 ( .IN1(b[10]), .IN2(a[10]), .IN3(b[10]), .IN4(n2), .IN5(a[10]), 
        .IN6(n2), .Q(n3) );
  AO222X1 U5 ( .IN1(b[11]), .IN2(a[11]), .IN3(b[11]), .IN4(n3), .IN5(a[11]), 
        .IN6(n3), .Q(n4) );
  AO222X1 U6 ( .IN1(b[12]), .IN2(a[12]), .IN3(b[12]), .IN4(n4), .IN5(a[12]), 
        .IN6(n4), .Q(n5) );
  AO222X1 U7 ( .IN1(b[13]), .IN2(a[13]), .IN3(b[13]), .IN4(n5), .IN5(a[13]), 
        .IN6(n5), .Q(n6) );
  AO222X1 U8 ( .IN1(b[14]), .IN2(a[14]), .IN3(b[14]), .IN4(n6), .IN5(a[14]), 
        .IN6(n6), .Q(n7) );
  AO222X1 U9 ( .IN1(b[15]), .IN2(a[15]), .IN3(b[15]), .IN4(n7), .IN5(a[15]), 
        .IN6(n7), .Q(n8) );
  AO222X1 U10 ( .IN1(b[16]), .IN2(a[16]), .IN3(b[16]), .IN4(n8), .IN5(a[16]), 
        .IN6(n8), .Q(n9) );
  AO222X1 U11 ( .IN1(b[17]), .IN2(a[17]), .IN3(b[17]), .IN4(n9), .IN5(a[17]), 
        .IN6(n9), .Q(n10) );
  AO222X1 U12 ( .IN1(b[18]), .IN2(a[18]), .IN3(b[18]), .IN4(n10), .IN5(a[18]), 
        .IN6(n10), .Q(n11) );
  AO222X1 U13 ( .IN1(b[19]), .IN2(a[19]), .IN3(b[19]), .IN4(n11), .IN5(a[19]), 
        .IN6(n11), .Q(n12) );
  AO222X1 U14 ( .IN1(b[20]), .IN2(a[20]), .IN3(b[20]), .IN4(n12), .IN5(a[20]), 
        .IN6(n12), .Q(n13) );
  AO222X1 U15 ( .IN1(b[21]), .IN2(a[21]), .IN3(b[21]), .IN4(n13), .IN5(a[21]), 
        .IN6(n13), .Q(n14) );
  AO222X1 U16 ( .IN1(b[22]), .IN2(a[22]), .IN3(b[22]), .IN4(n14), .IN5(a[22]), 
        .IN6(n14), .Q(intadd_0_CI) );
  XOR3X1 U17 ( .IN1(intadd_0_n1), .IN2(a[47]), .IN3(b[47]), .Q(out[47]) );
endmodule


module csa51squ_73 ( sumout, in1, in2, in3, cout_50_, cout_49_, cout_48_, 
        cout_47_, cout_46_, cout_44_, cout_42_, cout_40_, cout_38_, cout_36_, 
        cout_34_, cout_32_, cout_30_, cout_28_, cout_27_, cout_7__BAR, cout_6_, 
        cout_5_, cout_4_, cout_3_, cout_2_, cout_1_, cout_0_, cout_8__BAR, 
        cout_9__BAR, cout_10__BAR, cout_11__BAR, cout_12__BAR, cout_13__BAR, 
        cout_14__BAR, cout_15__BAR, cout_16__BAR, cout_17__BAR, cout_18__BAR, 
        cout_19__BAR, cout_20__BAR, cout_21__BAR, cout_22__BAR, cout_23__BAR, 
        cout_24__BAR, cout_25__BAR, cout_26__BAR, cout_29__BAR, cout_31__BAR, 
        cout_33__BAR, cout_35__BAR, cout_37__BAR, cout_39__BAR, cout_41__BAR, 
        cout_43__BAR, cout_45__BAR );
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  output cout_50_, cout_49_, cout_48_, cout_47_, cout_46_, cout_44_, cout_42_,
         cout_40_, cout_38_, cout_36_, cout_34_, cout_32_, cout_30_, cout_28_,
         cout_27_, cout_7__BAR, cout_6_, cout_5_, cout_4_, cout_3_, cout_2_,
         cout_1_, cout_0_, cout_8__BAR, cout_9__BAR, cout_10__BAR,
         cout_11__BAR, cout_12__BAR, cout_13__BAR, cout_14__BAR, cout_15__BAR,
         cout_16__BAR, cout_17__BAR, cout_18__BAR, cout_19__BAR, cout_20__BAR,
         cout_21__BAR, cout_22__BAR, cout_23__BAR, cout_24__BAR, cout_25__BAR,
         cout_26__BAR, cout_29__BAR, cout_31__BAR, cout_33__BAR, cout_35__BAR,
         cout_37__BAR, cout_39__BAR, cout_41__BAR, cout_43__BAR, cout_45__BAR;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11;

  NAND2X0 U1 ( .IN1(in2[8]), .IN2(in1[8]), .QN(cout_8__BAR) );
  NAND2X0 U2 ( .IN1(in2[9]), .IN2(in1[9]), .QN(cout_9__BAR) );
  NAND2X0 U3 ( .IN1(in2[10]), .IN2(in1[10]), .QN(cout_10__BAR) );
  NAND2X0 U4 ( .IN1(in2[11]), .IN2(in1[11]), .QN(cout_11__BAR) );
  NAND2X0 U5 ( .IN1(in2[12]), .IN2(in1[12]), .QN(cout_12__BAR) );
  NAND2X0 U6 ( .IN1(in2[13]), .IN2(in1[13]), .QN(cout_13__BAR) );
  NAND2X0 U7 ( .IN1(in2[14]), .IN2(in1[14]), .QN(cout_14__BAR) );
  NAND2X0 U8 ( .IN1(in2[15]), .IN2(in1[15]), .QN(cout_15__BAR) );
  NAND2X0 U9 ( .IN1(in2[16]), .IN2(in1[16]), .QN(cout_16__BAR) );
  NAND2X0 U10 ( .IN1(in2[17]), .IN2(in1[17]), .QN(cout_17__BAR) );
  NAND2X0 U11 ( .IN1(in2[18]), .IN2(in1[18]), .QN(cout_18__BAR) );
  NAND2X0 U12 ( .IN1(in2[19]), .IN2(in1[19]), .QN(cout_19__BAR) );
  NAND2X0 U13 ( .IN1(in2[20]), .IN2(in1[20]), .QN(cout_20__BAR) );
  NAND2X0 U14 ( .IN1(in2[21]), .IN2(in1[21]), .QN(cout_21__BAR) );
  NAND2X0 U15 ( .IN1(in2[22]), .IN2(in1[22]), .QN(cout_22__BAR) );
  NAND2X0 U16 ( .IN1(in2[23]), .IN2(in1[23]), .QN(cout_23__BAR) );
  NAND2X0 U17 ( .IN1(in2[24]), .IN2(in1[24]), .QN(cout_24__BAR) );
  NAND2X0 U18 ( .IN1(in2[25]), .IN2(in1[25]), .QN(cout_25__BAR) );
  NAND2X0 U19 ( .IN1(in2[26]), .IN2(in1[26]), .QN(cout_26__BAR) );
  NAND2X0 U20 ( .IN1(in2[29]), .IN2(in1[29]), .QN(cout_29__BAR) );
  NAND2X0 U21 ( .IN1(in2[31]), .IN2(in1[31]), .QN(cout_31__BAR) );
  NAND2X0 U22 ( .IN1(in2[33]), .IN2(in1[33]), .QN(cout_33__BAR) );
  NAND2X0 U23 ( .IN1(in2[35]), .IN2(in1[35]), .QN(cout_35__BAR) );
  NAND2X0 U24 ( .IN1(in2[37]), .IN2(in1[37]), .QN(cout_37__BAR) );
  NAND2X0 U25 ( .IN1(in2[39]), .IN2(in1[39]), .QN(cout_39__BAR) );
  NAND2X0 U26 ( .IN1(in2[41]), .IN2(in1[41]), .QN(cout_41__BAR) );
  NAND2X0 U27 ( .IN1(in2[43]), .IN2(in1[43]), .QN(cout_43__BAR) );
  NAND2X0 U28 ( .IN1(in2[45]), .IN2(in1[45]), .QN(cout_45__BAR) );
  NAND2X0 U29 ( .IN1(in2[7]), .IN2(in1[7]), .QN(cout_7__BAR) );
  NAND2X0 U30 ( .IN1(n1), .IN2(cout_27_), .QN(sumout[27]) );
  NAND2X0 U31 ( .IN1(in1[27]), .IN2(in2[27]), .QN(n1) );
  NAND2X0 U32 ( .IN1(n2), .IN2(cout_28_), .QN(sumout[28]) );
  NAND2X0 U33 ( .IN1(in1[28]), .IN2(in2[28]), .QN(n2) );
  NAND2X0 U34 ( .IN1(n3), .IN2(cout_30_), .QN(sumout[30]) );
  NAND2X0 U35 ( .IN1(in1[30]), .IN2(in2[30]), .QN(n3) );
  NAND2X0 U36 ( .IN1(n4), .IN2(cout_32_), .QN(sumout[32]) );
  NAND2X0 U37 ( .IN1(in1[32]), .IN2(in2[32]), .QN(n4) );
  NAND2X0 U38 ( .IN1(n5), .IN2(cout_34_), .QN(sumout[34]) );
  NAND2X0 U39 ( .IN1(in1[34]), .IN2(in2[34]), .QN(n5) );
  NAND2X0 U40 ( .IN1(n6), .IN2(cout_36_), .QN(sumout[36]) );
  NAND2X0 U41 ( .IN1(in1[36]), .IN2(in2[36]), .QN(n6) );
  NAND2X0 U42 ( .IN1(n7), .IN2(cout_38_), .QN(sumout[38]) );
  NAND2X0 U43 ( .IN1(in1[38]), .IN2(in2[38]), .QN(n7) );
  NAND2X0 U44 ( .IN1(n8), .IN2(cout_40_), .QN(sumout[40]) );
  NAND2X0 U45 ( .IN1(in1[40]), .IN2(in2[40]), .QN(n8) );
  NAND2X0 U46 ( .IN1(n9), .IN2(cout_42_), .QN(sumout[42]) );
  NAND2X0 U47 ( .IN1(in1[42]), .IN2(in2[42]), .QN(n9) );
  NAND2X0 U48 ( .IN1(n10), .IN2(cout_44_), .QN(sumout[44]) );
  NAND2X0 U49 ( .IN1(in1[44]), .IN2(in2[44]), .QN(n10) );
  NAND2X0 U50 ( .IN1(n11), .IN2(cout_46_), .QN(sumout[46]) );
  NAND2X0 U51 ( .IN1(in1[46]), .IN2(in2[46]), .QN(n11) );
  OR2X1 U52 ( .IN1(in2[27]), .IN2(in1[27]), .Q(cout_27_) );
  OR2X1 U53 ( .IN1(in2[28]), .IN2(in1[28]), .Q(cout_28_) );
  OR2X1 U54 ( .IN1(in2[30]), .IN2(in1[30]), .Q(cout_30_) );
  OR2X1 U55 ( .IN1(in2[32]), .IN2(in1[32]), .Q(cout_32_) );
  OR2X1 U56 ( .IN1(in2[34]), .IN2(in1[34]), .Q(cout_34_) );
  OR2X1 U57 ( .IN1(in2[36]), .IN2(in1[36]), .Q(cout_36_) );
  OR2X1 U58 ( .IN1(in2[38]), .IN2(in1[38]), .Q(cout_38_) );
  OR2X1 U59 ( .IN1(in2[40]), .IN2(in1[40]), .Q(cout_40_) );
  OR2X1 U60 ( .IN1(in2[42]), .IN2(in1[42]), .Q(cout_42_) );
  OR2X1 U61 ( .IN1(in2[44]), .IN2(in1[44]), .Q(cout_44_) );
  OR2X1 U62 ( .IN1(in2[46]), .IN2(in1[46]), .Q(cout_46_) );
  OA21X1 U63 ( .IN1(in2[8]), .IN2(in1[8]), .IN3(cout_8__BAR), .Q(sumout[8]) );
  OA21X1 U64 ( .IN1(in2[9]), .IN2(in1[9]), .IN3(cout_9__BAR), .Q(sumout[9]) );
  OA21X1 U65 ( .IN1(in2[10]), .IN2(in1[10]), .IN3(cout_10__BAR), .Q(sumout[10]) );
  OA21X1 U66 ( .IN1(in2[11]), .IN2(in1[11]), .IN3(cout_11__BAR), .Q(sumout[11]) );
  OA21X1 U67 ( .IN1(in2[12]), .IN2(in1[12]), .IN3(cout_12__BAR), .Q(sumout[12]) );
  OA21X1 U68 ( .IN1(in2[13]), .IN2(in1[13]), .IN3(cout_13__BAR), .Q(sumout[13]) );
  OA21X1 U69 ( .IN1(in2[14]), .IN2(in1[14]), .IN3(cout_14__BAR), .Q(sumout[14]) );
  OA21X1 U70 ( .IN1(in2[15]), .IN2(in1[15]), .IN3(cout_15__BAR), .Q(sumout[15]) );
  OA21X1 U71 ( .IN1(in2[16]), .IN2(in1[16]), .IN3(cout_16__BAR), .Q(sumout[16]) );
  OA21X1 U72 ( .IN1(in2[17]), .IN2(in1[17]), .IN3(cout_17__BAR), .Q(sumout[17]) );
  OA21X1 U73 ( .IN1(in2[18]), .IN2(in1[18]), .IN3(cout_18__BAR), .Q(sumout[18]) );
  OA21X1 U74 ( .IN1(in2[19]), .IN2(in1[19]), .IN3(cout_19__BAR), .Q(sumout[19]) );
  OA21X1 U75 ( .IN1(in2[20]), .IN2(in1[20]), .IN3(cout_20__BAR), .Q(sumout[20]) );
  OA21X1 U76 ( .IN1(in2[21]), .IN2(in1[21]), .IN3(cout_21__BAR), .Q(sumout[21]) );
  OA21X1 U77 ( .IN1(in2[22]), .IN2(in1[22]), .IN3(cout_22__BAR), .Q(sumout[22]) );
  OA21X1 U78 ( .IN1(in2[23]), .IN2(in1[23]), .IN3(cout_23__BAR), .Q(sumout[23]) );
  OA21X1 U79 ( .IN1(in2[24]), .IN2(in1[24]), .IN3(cout_24__BAR), .Q(sumout[24]) );
  OA21X1 U80 ( .IN1(in2[25]), .IN2(in1[25]), .IN3(cout_25__BAR), .Q(sumout[25]) );
  OA21X1 U81 ( .IN1(in2[26]), .IN2(in1[26]), .IN3(cout_26__BAR), .Q(sumout[26]) );
  OA21X1 U82 ( .IN1(in2[29]), .IN2(in1[29]), .IN3(cout_29__BAR), .Q(sumout[29]) );
  OA21X1 U83 ( .IN1(in2[31]), .IN2(in1[31]), .IN3(cout_31__BAR), .Q(sumout[31]) );
  OA21X1 U84 ( .IN1(in2[33]), .IN2(in1[33]), .IN3(cout_33__BAR), .Q(sumout[33]) );
  OA21X1 U85 ( .IN1(in2[35]), .IN2(in1[35]), .IN3(cout_35__BAR), .Q(sumout[35]) );
  OA21X1 U86 ( .IN1(in2[37]), .IN2(in1[37]), .IN3(cout_37__BAR), .Q(sumout[37]) );
  OA21X1 U87 ( .IN1(in2[39]), .IN2(in1[39]), .IN3(cout_39__BAR), .Q(sumout[39]) );
  OA21X1 U88 ( .IN1(in2[41]), .IN2(in1[41]), .IN3(cout_41__BAR), .Q(sumout[41]) );
  OA21X1 U89 ( .IN1(in2[43]), .IN2(in1[43]), .IN3(cout_43__BAR), .Q(sumout[43]) );
  OA21X1 U90 ( .IN1(in2[45]), .IN2(in1[45]), .IN3(cout_45__BAR), .Q(sumout[45]) );
  XOR2X1 U91 ( .IN1(in1[47]), .IN2(in2[47]), .Q(sumout[47]) );
endmodule


module csa51squ_74 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;


  AO222X1 U1 ( .IN1(in2[6]), .IN2(in3[6]), .IN3(in2[6]), .IN4(in1[6]), .IN5(
        in3[6]), .IN6(in1[6]), .Q(cout[6]) );
  FADDX1 U2 ( .A(in1[10]), .B(in2[10]), .CI(in3[10]), .CO(cout[10]), .S(
        sumout[10]) );
  FADDX1 U3 ( .A(in1[11]), .B(in2[11]), .CI(in3[11]), .CO(cout[11]), .S(
        sumout[11]) );
  FADDX1 U4 ( .A(in1[12]), .B(in2[12]), .CI(in3[12]), .CO(cout[12]), .S(
        sumout[12]) );
  FADDX1 U5 ( .A(in1[13]), .B(in2[13]), .CI(in3[13]), .CO(cout[13]), .S(
        sumout[13]) );
  FADDX1 U6 ( .A(in1[14]), .B(in2[14]), .CI(in3[14]), .CO(cout[14]), .S(
        sumout[14]) );
  FADDX1 U7 ( .A(in1[15]), .B(in2[15]), .CI(in3[15]), .CO(cout[15]), .S(
        sumout[15]) );
  FADDX1 U8 ( .A(in1[16]), .B(in2[16]), .CI(in3[16]), .CO(cout[16]), .S(
        sumout[16]) );
  FADDX1 U9 ( .A(in1[17]), .B(in2[17]), .CI(in3[17]), .CO(cout[17]), .S(
        sumout[17]) );
  FADDX1 U10 ( .A(in1[18]), .B(in2[18]), .CI(in3[18]), .CO(cout[18]), .S(
        sumout[18]) );
  FADDX1 U11 ( .A(in1[19]), .B(in2[19]), .CI(in3[19]), .CO(cout[19]), .S(
        sumout[19]) );
  FADDX1 U12 ( .A(in1[20]), .B(in2[20]), .CI(in3[20]), .CO(cout[20]), .S(
        sumout[20]) );
  FADDX1 U13 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U14 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U15 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U16 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U17 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U18 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U19 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U20 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U21 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U22 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U23 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U24 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
  FADDX1 U25 ( .A(in1[33]), .B(in2[33]), .CI(in3[33]), .CO(cout[33]), .S(
        sumout[33]) );
  FADDX1 U26 ( .A(in1[34]), .B(in2[34]), .CI(in3[34]), .CO(cout[34]), .S(
        sumout[34]) );
  FADDX1 U27 ( .A(in1[35]), .B(in2[35]), .CI(in3[35]), .CO(cout[35]), .S(
        sumout[35]) );
  FADDX1 U28 ( .A(in1[36]), .B(in2[36]), .CI(in3[36]), .CO(cout[36]), .S(
        sumout[36]) );
  FADDX1 U29 ( .A(in1[37]), .B(in2[37]), .CI(in3[37]), .CO(cout[37]), .S(
        sumout[37]) );
  FADDX1 U30 ( .A(in1[38]), .B(in2[38]), .CI(in3[38]), .CO(cout[38]), .S(
        sumout[38]) );
  FADDX1 U31 ( .A(in1[39]), .B(in2[39]), .CI(in3[39]), .CO(cout[39]), .S(
        sumout[39]) );
  FADDX1 U32 ( .A(in1[40]), .B(in2[40]), .CI(in3[40]), .CO(cout[40]), .S(
        sumout[40]) );
  FADDX1 U33 ( .A(in1[41]), .B(in2[41]), .CI(in3[41]), .CO(cout[41]), .S(
        sumout[41]) );
  FADDX1 U34 ( .A(in1[42]), .B(in2[42]), .CI(in3[42]), .CO(cout[42]), .S(
        sumout[42]) );
  FADDX1 U35 ( .A(in1[43]), .B(in2[43]), .CI(in3[43]), .CO(cout[43]), .S(
        sumout[43]) );
  FADDX1 U36 ( .A(in1[44]), .B(in2[44]), .CI(in3[44]), .CO(cout[44]), .S(
        sumout[44]) );
  FADDX1 U37 ( .A(in1[45]), .B(in2[45]), .CI(in3[45]), .CO(cout[45]), .S(
        sumout[45]) );
  FADDX1 U38 ( .A(in1[46]), .B(in2[46]), .CI(in3[46]), .CO(cout[46]), .S(
        sumout[46]) );
  XOR3X1 U39 ( .IN1(in2[47]), .IN2(in3[47]), .IN3(in1[47]), .Q(sumout[47]) );
  FADDX1 U40 ( .A(in1[7]), .B(in2[7]), .CI(in3[7]), .CO(cout[7]), .S(sumout[7]) );
  FADDX1 U41 ( .A(in1[8]), .B(in2[8]), .CI(in3[8]), .CO(cout[8]), .S(sumout[8]) );
  FADDX1 U42 ( .A(in1[9]), .B(in2[9]), .CI(in3[9]), .CO(cout[9]), .S(sumout[9]) );
endmodule


module csa51squ_75 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14;

  AND2X1 U1 ( .IN1(in2[7]), .IN2(in1[7]), .Q(cout[7]) );
  NOR2X0 U2 ( .IN1(in2[7]), .IN2(in1[7]), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(cout[7]), .QN(sumout[7]) );
  AND2X1 U4 ( .IN1(in2[8]), .IN2(in1[8]), .Q(cout[8]) );
  NOR2X0 U5 ( .IN1(in2[8]), .IN2(in1[8]), .QN(n2) );
  NOR2X0 U6 ( .IN1(n2), .IN2(cout[8]), .QN(sumout[8]) );
  AND2X1 U7 ( .IN1(in2[9]), .IN2(in1[9]), .Q(cout[9]) );
  NOR2X0 U8 ( .IN1(in2[9]), .IN2(in1[9]), .QN(n3) );
  NOR2X0 U9 ( .IN1(n3), .IN2(cout[9]), .QN(sumout[9]) );
  AND2X1 U10 ( .IN1(in2[10]), .IN2(in1[10]), .Q(cout[10]) );
  NOR2X0 U11 ( .IN1(in2[10]), .IN2(in1[10]), .QN(n4) );
  NOR2X0 U12 ( .IN1(n4), .IN2(cout[10]), .QN(sumout[10]) );
  AND2X1 U13 ( .IN1(in2[11]), .IN2(in1[11]), .Q(cout[11]) );
  NOR2X0 U14 ( .IN1(in2[11]), .IN2(in1[11]), .QN(n5) );
  NOR2X0 U15 ( .IN1(n5), .IN2(cout[11]), .QN(sumout[11]) );
  AND2X1 U16 ( .IN1(in2[12]), .IN2(in1[12]), .Q(cout[12]) );
  NOR2X0 U17 ( .IN1(in2[12]), .IN2(in1[12]), .QN(n6) );
  NOR2X0 U18 ( .IN1(n6), .IN2(cout[12]), .QN(sumout[12]) );
  AND2X1 U19 ( .IN1(in2[5]), .IN2(in1[5]), .Q(cout[5]) );
  AND2X1 U20 ( .IN1(in2[6]), .IN2(in1[6]), .Q(cout[6]) );
  NOR2X0 U21 ( .IN1(in2[6]), .IN2(in1[6]), .QN(n7) );
  NOR2X0 U22 ( .IN1(n7), .IN2(cout[6]), .QN(sumout[6]) );
  AND2X1 U23 ( .IN1(in3[40]), .IN2(in2[40]), .Q(cout[40]) );
  NOR2X0 U24 ( .IN1(in3[40]), .IN2(in2[40]), .QN(n8) );
  NOR2X0 U25 ( .IN1(n8), .IN2(cout[40]), .QN(sumout[40]) );
  AND2X1 U26 ( .IN1(in3[41]), .IN2(in2[41]), .Q(cout[41]) );
  NOR2X0 U27 ( .IN1(in3[41]), .IN2(in2[41]), .QN(n9) );
  NOR2X0 U28 ( .IN1(n9), .IN2(cout[41]), .QN(sumout[41]) );
  AND2X1 U29 ( .IN1(in3[42]), .IN2(in2[42]), .Q(cout[42]) );
  NOR2X0 U30 ( .IN1(in3[42]), .IN2(in2[42]), .QN(n10) );
  NOR2X0 U31 ( .IN1(n10), .IN2(cout[42]), .QN(sumout[42]) );
  AND2X1 U32 ( .IN1(in3[43]), .IN2(in2[43]), .Q(cout[43]) );
  NOR2X0 U33 ( .IN1(in3[43]), .IN2(in2[43]), .QN(n11) );
  NOR2X0 U34 ( .IN1(n11), .IN2(cout[43]), .QN(sumout[43]) );
  AND2X1 U35 ( .IN1(in3[44]), .IN2(in2[44]), .Q(cout[44]) );
  NOR2X0 U36 ( .IN1(in3[44]), .IN2(in2[44]), .QN(n12) );
  NOR2X0 U37 ( .IN1(n12), .IN2(cout[44]), .QN(sumout[44]) );
  AND2X1 U38 ( .IN1(in3[45]), .IN2(in2[45]), .Q(cout[45]) );
  NOR2X0 U39 ( .IN1(in3[45]), .IN2(in2[45]), .QN(n13) );
  NOR2X0 U40 ( .IN1(n13), .IN2(cout[45]), .QN(sumout[45]) );
  AND2X1 U41 ( .IN1(in3[46]), .IN2(in2[46]), .Q(cout[46]) );
  NOR2X0 U42 ( .IN1(in3[46]), .IN2(in2[46]), .QN(n14) );
  NOR2X0 U43 ( .IN1(n14), .IN2(cout[46]), .QN(sumout[46]) );
  INVX0 U44 ( .INP(in3[47]), .ZN(sumout[47]) );
  FADDX1 U45 ( .A(in1[13]), .B(in2[13]), .CI(in3[13]), .CO(cout[13]), .S(
        sumout[13]) );
  FADDX1 U46 ( .A(in1[14]), .B(in2[14]), .CI(in3[14]), .CO(cout[14]), .S(
        sumout[14]) );
  FADDX1 U47 ( .A(in1[15]), .B(in2[15]), .CI(in3[15]), .CO(cout[15]), .S(
        sumout[15]) );
  FADDX1 U48 ( .A(in1[16]), .B(in2[16]), .CI(in3[16]), .CO(cout[16]), .S(
        sumout[16]) );
  FADDX1 U49 ( .A(in1[17]), .B(in2[17]), .CI(in3[17]), .CO(cout[17]), .S(
        sumout[17]) );
  FADDX1 U50 ( .A(in1[18]), .B(in2[18]), .CI(in3[18]), .CO(cout[18]), .S(
        sumout[18]) );
  FADDX1 U51 ( .A(in1[19]), .B(in2[19]), .CI(in3[19]), .CO(cout[19]), .S(
        sumout[19]) );
  FADDX1 U52 ( .A(in1[20]), .B(in2[20]), .CI(in3[20]), .CO(cout[20]), .S(
        sumout[20]) );
  FADDX1 U53 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U54 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U55 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U56 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U57 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U58 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U59 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U60 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U61 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U62 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U63 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U64 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
  FADDX1 U65 ( .A(in1[33]), .B(in2[33]), .CI(in3[33]), .CO(cout[33]), .S(
        sumout[33]) );
  FADDX1 U66 ( .A(in1[34]), .B(in2[34]), .CI(in3[34]), .CO(cout[34]), .S(
        sumout[34]) );
  FADDX1 U67 ( .A(in1[35]), .B(in2[35]), .CI(in3[35]), .CO(cout[35]), .S(
        sumout[35]) );
  FADDX1 U68 ( .A(in1[36]), .B(in2[36]), .CI(in3[36]), .CO(cout[36]), .S(
        sumout[36]) );
  FADDX1 U69 ( .A(in1[37]), .B(in2[37]), .CI(in3[37]), .CO(cout[37]), .S(
        sumout[37]) );
  FADDX1 U70 ( .A(in1[38]), .B(in2[38]), .CI(in3[38]), .CO(cout[38]), .S(
        sumout[38]) );
  FADDX1 U71 ( .A(in1[39]), .B(in2[39]), .CI(in3[39]), .CO(cout[39]), .S(
        sumout[39]) );
endmodule


module csa51squ_76 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17;

  NBUFFX2 U1 ( .INP(in1[6]), .Z(sumout[6]) );
  NBUFFX2 U2 ( .INP(in1[7]), .Z(sumout[7]) );
  NBUFFX2 U3 ( .INP(in1[8]), .Z(sumout[8]) );
  NBUFFX2 U4 ( .INP(in1[9]), .Z(sumout[9]) );
  NBUFFX2 U5 ( .INP(in1[10]), .Z(sumout[10]) );
  NBUFFX2 U6 ( .INP(in1[11]), .Z(sumout[11]) );
  AND2X1 U7 ( .IN1(in3[13]), .IN2(in1[13]), .Q(cout[13]) );
  NOR2X0 U8 ( .IN1(in3[13]), .IN2(in1[13]), .QN(n7) );
  NOR2X0 U9 ( .IN1(n7), .IN2(cout[13]), .QN(sumout[13]) );
  AND2X1 U10 ( .IN1(in3[15]), .IN2(in1[15]), .Q(cout[15]) );
  NOR2X0 U11 ( .IN1(in3[15]), .IN2(in1[15]), .QN(n8) );
  NOR2X0 U12 ( .IN1(n8), .IN2(cout[15]), .QN(sumout[15]) );
  AND2X1 U13 ( .IN1(in3[17]), .IN2(in1[17]), .Q(cout[17]) );
  NOR2X0 U14 ( .IN1(in3[17]), .IN2(in1[17]), .QN(n9) );
  NOR2X0 U15 ( .IN1(n9), .IN2(cout[17]), .QN(sumout[17]) );
  AND2X1 U16 ( .IN1(in3[43]), .IN2(in2[43]), .Q(cout[43]) );
  NOR2X0 U17 ( .IN1(in3[43]), .IN2(in2[43]), .QN(n10) );
  NOR2X0 U18 ( .IN1(n10), .IN2(cout[43]), .QN(sumout[43]) );
  AND2X1 U19 ( .IN1(in3[44]), .IN2(in2[44]), .Q(cout[44]) );
  NOR2X0 U20 ( .IN1(in3[44]), .IN2(in2[44]), .QN(n11) );
  NOR2X0 U21 ( .IN1(n11), .IN2(cout[44]), .QN(sumout[44]) );
  AND2X1 U22 ( .IN1(in3[45]), .IN2(in2[45]), .Q(cout[45]) );
  NOR2X0 U23 ( .IN1(in3[45]), .IN2(in2[45]), .QN(n12) );
  NOR2X0 U24 ( .IN1(n12), .IN2(cout[45]), .QN(sumout[45]) );
  AND2X1 U25 ( .IN1(in3[46]), .IN2(in2[46]), .Q(cout[46]) );
  NOR2X0 U26 ( .IN1(in3[46]), .IN2(in2[46]), .QN(n13) );
  NOR2X0 U27 ( .IN1(n13), .IN2(cout[46]), .QN(sumout[46]) );
  XOR2X1 U28 ( .IN1(in3[47]), .IN2(in2[47]), .Q(sumout[47]) );
  AND2X1 U29 ( .IN1(in3[12]), .IN2(in1[12]), .Q(cout[12]) );
  NOR2X0 U30 ( .IN1(in3[12]), .IN2(in1[12]), .QN(n14) );
  NOR2X0 U31 ( .IN1(n14), .IN2(cout[12]), .QN(sumout[12]) );
  AND2X1 U32 ( .IN1(in3[14]), .IN2(in1[14]), .Q(cout[14]) );
  NOR2X0 U33 ( .IN1(in3[14]), .IN2(in1[14]), .QN(n15) );
  NOR2X0 U34 ( .IN1(n15), .IN2(cout[14]), .QN(sumout[14]) );
  AND2X1 U35 ( .IN1(in3[16]), .IN2(in1[16]), .Q(cout[16]) );
  NOR2X0 U36 ( .IN1(in3[16]), .IN2(in1[16]), .QN(n16) );
  NOR2X0 U37 ( .IN1(n16), .IN2(cout[16]), .QN(sumout[16]) );
  AND2X1 U38 ( .IN1(in3[18]), .IN2(in1[18]), .Q(cout[18]) );
  NOR2X0 U39 ( .IN1(in3[18]), .IN2(in1[18]), .QN(n17) );
  NOR2X0 U40 ( .IN1(n17), .IN2(cout[18]), .QN(sumout[18]) );
  FADDX1 U41 ( .A(in1[19]), .B(in2[19]), .CI(in3[19]), .CO(cout[19]), .S(
        sumout[19]) );
  FADDX1 U42 ( .A(in1[20]), .B(in2[20]), .CI(in3[20]), .CO(cout[20]), .S(
        sumout[20]) );
  FADDX1 U43 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U44 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U45 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U46 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U47 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U48 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U49 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U50 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U51 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U52 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U53 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U54 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
  FADDX1 U55 ( .A(in1[33]), .B(in2[33]), .CI(in3[33]), .CO(cout[33]), .S(
        sumout[33]) );
  FADDX1 U56 ( .A(in1[34]), .B(in2[34]), .CI(in3[34]), .CO(cout[34]), .S(
        sumout[34]) );
  FADDX1 U57 ( .A(in1[35]), .B(in2[35]), .CI(in3[35]), .CO(cout[35]), .S(
        sumout[35]) );
  FADDX1 U58 ( .A(in1[36]), .B(in2[36]), .CI(in3[36]), .CO(cout[36]), .S(
        sumout[36]) );
  FADDX1 U59 ( .A(in1[37]), .B(in2[37]), .CI(in3[37]), .CO(cout[37]), .S(
        sumout[37]) );
  FADDX1 U60 ( .A(in1[38]), .B(in2[38]), .CI(in3[38]), .CO(cout[38]), .S(
        sumout[38]) );
  FADDX1 U61 ( .A(in1[39]), .B(in2[39]), .CI(in3[39]), .CO(cout[39]), .S(
        sumout[39]) );
  FADDX1 U62 ( .A(in1[40]), .B(in2[40]), .CI(in3[40]), .CO(cout[40]), .S(
        sumout[40]) );
  FADDX1 U63 ( .A(in1[41]), .B(in2[41]), .CI(in3[41]), .CO(cout[41]), .S(
        sumout[41]) );
  FADDX1 U64 ( .A(in1[42]), .B(in2[42]), .CI(in3[42]), .CO(cout[42]), .S(
        sumout[42]) );
endmodule


module csa51squ_77 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19;

  NBUFFX2 U1 ( .INP(in2[46]), .Z(sumout[46]) );
  NBUFFX2 U2 ( .INP(in2[45]), .Z(sumout[45]) );
  NBUFFX2 U3 ( .INP(in2[44]), .Z(sumout[44]) );
  NBUFFX2 U4 ( .INP(in2[43]), .Z(sumout[43]) );
  NBUFFX2 U5 ( .INP(in2[42]), .Z(sumout[42]) );
  NBUFFX2 U6 ( .INP(in2[41]), .Z(sumout[41]) );
  NBUFFX2 U7 ( .INP(in2[40]), .Z(sumout[40]) );
  NBUFFX2 U8 ( .INP(in2[39]), .Z(sumout[39]) );
  AND2X1 U9 ( .IN1(in2[7]), .IN2(in1[7]), .Q(cout[7]) );
  NOR2X0 U10 ( .IN1(in2[7]), .IN2(in1[7]), .QN(n9) );
  NOR2X0 U11 ( .IN1(n9), .IN2(cout[7]), .QN(sumout[7]) );
  AND2X1 U12 ( .IN1(in2[8]), .IN2(in1[8]), .Q(cout[8]) );
  NOR2X0 U13 ( .IN1(in2[8]), .IN2(in1[8]), .QN(n10) );
  NOR2X0 U14 ( .IN1(n10), .IN2(cout[8]), .QN(sumout[8]) );
  AND2X1 U15 ( .IN1(in2[9]), .IN2(in1[9]), .Q(cout[9]) );
  NOR2X0 U16 ( .IN1(in2[9]), .IN2(in1[9]), .QN(n11) );
  NOR2X0 U17 ( .IN1(n11), .IN2(cout[9]), .QN(sumout[9]) );
  AND2X1 U18 ( .IN1(in2[4]), .IN2(in1[4]), .Q(cout[4]) );
  AND2X1 U19 ( .IN1(in2[5]), .IN2(in1[5]), .Q(cout[5]) );
  NOR2X0 U20 ( .IN1(in2[5]), .IN2(in1[5]), .QN(n12) );
  NOR2X0 U21 ( .IN1(n12), .IN2(cout[5]), .QN(sumout[5]) );
  AND2X1 U22 ( .IN1(in2[6]), .IN2(in1[6]), .Q(cout[6]) );
  NOR2X0 U23 ( .IN1(in2[6]), .IN2(in1[6]), .QN(n13) );
  NOR2X0 U24 ( .IN1(n13), .IN2(cout[6]), .QN(sumout[6]) );
  AND2X1 U25 ( .IN1(in3[33]), .IN2(in2[33]), .Q(cout[33]) );
  NOR2X0 U26 ( .IN1(in3[33]), .IN2(in2[33]), .QN(n14) );
  NOR2X0 U27 ( .IN1(n14), .IN2(cout[33]), .QN(sumout[33]) );
  AND2X1 U28 ( .IN1(in3[34]), .IN2(in2[34]), .Q(cout[34]) );
  NOR2X0 U29 ( .IN1(in3[34]), .IN2(in2[34]), .QN(n15) );
  NOR2X0 U30 ( .IN1(n15), .IN2(cout[34]), .QN(sumout[34]) );
  AND2X1 U31 ( .IN1(in3[35]), .IN2(in2[35]), .Q(cout[35]) );
  NOR2X0 U32 ( .IN1(in3[35]), .IN2(in2[35]), .QN(n16) );
  NOR2X0 U33 ( .IN1(n16), .IN2(cout[35]), .QN(sumout[35]) );
  AND2X1 U34 ( .IN1(in3[36]), .IN2(in2[36]), .Q(cout[36]) );
  NOR2X0 U35 ( .IN1(in3[36]), .IN2(in2[36]), .QN(n17) );
  NOR2X0 U36 ( .IN1(n17), .IN2(cout[36]), .QN(sumout[36]) );
  AND2X1 U37 ( .IN1(in3[37]), .IN2(in2[37]), .Q(cout[37]) );
  NOR2X0 U38 ( .IN1(in3[37]), .IN2(in2[37]), .QN(n18) );
  NOR2X0 U39 ( .IN1(n18), .IN2(cout[37]), .QN(sumout[37]) );
  AND2X1 U40 ( .IN1(in3[38]), .IN2(in2[38]), .Q(cout[38]) );
  NOR2X0 U41 ( .IN1(in3[38]), .IN2(in2[38]), .QN(n19) );
  NOR2X0 U42 ( .IN1(n19), .IN2(cout[38]), .QN(sumout[38]) );
  FADDX1 U43 ( .A(in1[10]), .B(in2[10]), .CI(in3[10]), .CO(cout[10]), .S(
        sumout[10]) );
  FADDX1 U44 ( .A(in1[11]), .B(in2[11]), .CI(in3[11]), .CO(cout[11]), .S(
        sumout[11]) );
  FADDX1 U45 ( .A(in1[12]), .B(in2[12]), .CI(in3[12]), .CO(cout[12]), .S(
        sumout[12]) );
  FADDX1 U46 ( .A(in1[13]), .B(in2[13]), .CI(in3[13]), .CO(cout[13]), .S(
        sumout[13]) );
  FADDX1 U47 ( .A(in1[14]), .B(in2[14]), .CI(in3[14]), .CO(cout[14]), .S(
        sumout[14]) );
  FADDX1 U48 ( .A(in1[15]), .B(in2[15]), .CI(in3[15]), .CO(cout[15]), .S(
        sumout[15]) );
  FADDX1 U49 ( .A(in1[16]), .B(in2[16]), .CI(in3[16]), .CO(cout[16]), .S(
        sumout[16]) );
  FADDX1 U50 ( .A(in1[17]), .B(in2[17]), .CI(in3[17]), .CO(cout[17]), .S(
        sumout[17]) );
  FADDX1 U51 ( .A(in1[18]), .B(in2[18]), .CI(in3[18]), .CO(cout[18]), .S(
        sumout[18]) );
  FADDX1 U52 ( .A(in1[19]), .B(in2[19]), .CI(in3[19]), .CO(cout[19]), .S(
        sumout[19]) );
  FADDX1 U53 ( .A(in1[20]), .B(in2[20]), .CI(in3[20]), .CO(cout[20]), .S(
        sumout[20]) );
  FADDX1 U54 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U55 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U56 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U57 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U58 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U59 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U60 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U61 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U62 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U63 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U64 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U65 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
endmodule


module csa51squ_78 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n7, n8, n9, n10, n11, n12, n13;

  NBUFFX2 U1 ( .INP(in1[12]), .Z(sumout[12]) );
  NBUFFX2 U2 ( .INP(in1[13]), .Z(sumout[13]) );
  NBUFFX2 U3 ( .INP(in1[14]), .Z(sumout[14]) );
  NBUFFX2 U4 ( .INP(in1[15]), .Z(sumout[15]) );
  NBUFFX2 U5 ( .INP(in1[16]), .Z(sumout[16]) );
  NBUFFX2 U6 ( .INP(in1[17]), .Z(sumout[17]) );
  AND2X1 U7 ( .IN1(in3[19]), .IN2(in1[19]), .Q(cout[19]) );
  NOR2X0 U8 ( .IN1(in3[19]), .IN2(in1[19]), .QN(n7) );
  NOR2X0 U9 ( .IN1(n7), .IN2(cout[19]), .QN(sumout[19]) );
  AND2X1 U10 ( .IN1(in3[44]), .IN2(in2[44]), .Q(cout[44]) );
  NOR2X0 U11 ( .IN1(in3[44]), .IN2(in2[44]), .QN(n8) );
  NOR2X0 U12 ( .IN1(n8), .IN2(cout[44]), .QN(sumout[44]) );
  AND2X1 U13 ( .IN1(in3[45]), .IN2(in2[45]), .Q(cout[45]) );
  NOR2X0 U14 ( .IN1(in3[45]), .IN2(in2[45]), .QN(n9) );
  NOR2X0 U15 ( .IN1(n9), .IN2(cout[45]), .QN(sumout[45]) );
  AND2X1 U16 ( .IN1(in3[46]), .IN2(in2[46]), .Q(cout[46]) );
  NOR2X0 U17 ( .IN1(in3[46]), .IN2(in2[46]), .QN(n10) );
  NOR2X0 U18 ( .IN1(n10), .IN2(cout[46]), .QN(sumout[46]) );
  XOR2X1 U19 ( .IN1(in3[47]), .IN2(in2[47]), .Q(sumout[47]) );
  AND2X1 U20 ( .IN1(in3[18]), .IN2(in1[18]), .Q(cout[18]) );
  NOR2X0 U21 ( .IN1(in3[18]), .IN2(in1[18]), .QN(n11) );
  NOR2X0 U22 ( .IN1(n11), .IN2(cout[18]), .QN(sumout[18]) );
  AND2X1 U23 ( .IN1(in3[20]), .IN2(in1[20]), .Q(cout[20]) );
  NOR2X0 U24 ( .IN1(in3[20]), .IN2(in1[20]), .QN(n12) );
  NOR2X0 U25 ( .IN1(n12), .IN2(cout[20]), .QN(sumout[20]) );
  INVX0 U26 ( .INP(in1[42]), .ZN(n13) );
  FADDX1 U27 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U28 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U29 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U30 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U31 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U32 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U33 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U34 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U35 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U36 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U37 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U38 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
  FADDX1 U39 ( .A(in1[33]), .B(in2[33]), .CI(in3[33]), .CO(cout[33]), .S(
        sumout[33]) );
  FADDX1 U40 ( .A(in1[34]), .B(in2[34]), .CI(in3[34]), .CO(cout[34]), .S(
        sumout[34]) );
  FADDX1 U41 ( .A(in1[35]), .B(in2[35]), .CI(in3[35]), .CO(cout[35]), .S(
        sumout[35]) );
  FADDX1 U42 ( .A(in1[36]), .B(in2[36]), .CI(in3[36]), .CO(cout[36]), .S(
        sumout[36]) );
  FADDX1 U43 ( .A(in1[37]), .B(in2[37]), .CI(in3[37]), .CO(cout[37]), .S(
        sumout[37]) );
  FADDX1 U44 ( .A(in1[38]), .B(in2[38]), .CI(in3[38]), .CO(cout[38]), .S(
        sumout[38]) );
  FADDX1 U45 ( .A(in1[39]), .B(in2[39]), .CI(in3[39]), .CO(cout[39]), .S(
        sumout[39]) );
  FADDX1 U46 ( .A(in1[40]), .B(in2[40]), .CI(in3[40]), .CO(cout[40]), .S(
        sumout[40]) );
  FADDX1 U47 ( .A(in1[41]), .B(in2[41]), .CI(in3[41]), .CO(cout[41]), .S(
        sumout[41]) );
  FADDX1 U48 ( .A(in1[42]), .B(in2[42]), .CI(in3[42]), .CO(cout[42]), .S(
        sumout[42]) );
  FADDX1 U49 ( .A(in2[43]), .B(in3[43]), .CI(n13), .CO(cout[43]), .S(
        sumout[43]) );
endmodule


module csa51squ_79 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n9, n10, n11, n12, n13, n14, n15;

  NBUFFX2 U1 ( .INP(in2[6]), .Z(sumout[6]) );
  NBUFFX2 U2 ( .INP(in2[7]), .Z(sumout[7]) );
  NBUFFX2 U3 ( .INP(in2[8]), .Z(sumout[8]) );
  NBUFFX2 U4 ( .INP(in3[42]), .Z(sumout[42]) );
  NBUFFX2 U5 ( .INP(in3[41]), .Z(sumout[41]) );
  NBUFFX2 U6 ( .INP(in3[39]), .Z(sumout[39]) );
  NBUFFX2 U7 ( .INP(in3[38]), .Z(sumout[38]) );
  NBUFFX2 U8 ( .INP(in3[40]), .Z(sumout[40]) );
  AND2X1 U9 ( .IN1(in2[13]), .IN2(in1[13]), .Q(cout[13]) );
  NOR2X0 U10 ( .IN1(in2[13]), .IN2(in1[13]), .QN(n9) );
  NOR2X0 U11 ( .IN1(n9), .IN2(cout[13]), .QN(sumout[13]) );
  AND2X1 U12 ( .IN1(in2[37]), .IN2(in3[37]), .Q(cout[37]) );
  INVX0 U13 ( .INP(in2[37]), .ZN(n15) );
  MUX21X1 U14 ( .IN1(in2[37]), .IN2(n15), .S(in3[37]), .Q(sumout[37]) );
  AND2X1 U15 ( .IN1(in2[9]), .IN2(in1[9]), .Q(cout[9]) );
  NOR2X0 U16 ( .IN1(in2[9]), .IN2(in1[9]), .QN(n10) );
  NOR2X0 U17 ( .IN1(n10), .IN2(cout[9]), .QN(sumout[9]) );
  AND2X1 U18 ( .IN1(in2[10]), .IN2(in1[10]), .Q(cout[10]) );
  NOR2X0 U19 ( .IN1(in2[10]), .IN2(in1[10]), .QN(n11) );
  NOR2X0 U20 ( .IN1(n11), .IN2(cout[10]), .QN(sumout[10]) );
  AND2X1 U21 ( .IN1(in2[11]), .IN2(in1[11]), .Q(cout[11]) );
  NOR2X0 U22 ( .IN1(in2[11]), .IN2(in1[11]), .QN(n12) );
  NOR2X0 U23 ( .IN1(n12), .IN2(cout[11]), .QN(sumout[11]) );
  AND2X1 U24 ( .IN1(in2[12]), .IN2(in1[12]), .Q(cout[12]) );
  NOR2X0 U25 ( .IN1(in2[12]), .IN2(in1[12]), .QN(n13) );
  NOR2X0 U26 ( .IN1(n13), .IN2(cout[12]), .QN(sumout[12]) );
  AND2X1 U27 ( .IN1(in2[14]), .IN2(in1[14]), .Q(cout[14]) );
  NOR2X0 U28 ( .IN1(in2[14]), .IN2(in1[14]), .QN(n14) );
  NOR2X0 U29 ( .IN1(n14), .IN2(cout[14]), .QN(sumout[14]) );
  FADDX1 U30 ( .A(in1[15]), .B(in2[15]), .CI(in3[15]), .CO(cout[15]), .S(
        sumout[15]) );
  FADDX1 U31 ( .A(in1[16]), .B(in2[16]), .CI(in3[16]), .CO(cout[16]), .S(
        sumout[16]) );
  FADDX1 U32 ( .A(in1[17]), .B(in2[17]), .CI(in3[17]), .CO(cout[17]), .S(
        sumout[17]) );
  FADDX1 U33 ( .A(in1[18]), .B(in2[18]), .CI(in3[18]), .CO(cout[18]), .S(
        sumout[18]) );
  FADDX1 U34 ( .A(in1[19]), .B(in2[19]), .CI(in3[19]), .CO(cout[19]), .S(
        sumout[19]) );
  FADDX1 U35 ( .A(in1[20]), .B(in2[20]), .CI(in3[20]), .CO(cout[20]), .S(
        sumout[20]) );
  FADDX1 U36 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U37 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U38 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U39 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U40 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U41 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U42 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U43 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U44 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U45 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U46 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U47 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
  FADDX1 U48 ( .A(in1[33]), .B(in2[33]), .CI(in3[33]), .CO(cout[33]), .S(
        sumout[33]) );
  FADDX1 U49 ( .A(in1[34]), .B(in2[34]), .CI(in3[34]), .CO(cout[34]), .S(
        sumout[34]) );
  FADDX1 U50 ( .A(in1[35]), .B(in2[35]), .CI(in3[35]), .CO(cout[35]), .S(
        sumout[35]) );
  FADDX1 U51 ( .A(in1[36]), .B(in3[36]), .CI(n15), .CO(cout[36]), .S(
        sumout[36]) );
endmodule


module csa51squ_80 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36;

  NBUFFX2 U1 ( .INP(in3[46]), .Z(sumout[46]) );
  NBUFFX2 U2 ( .INP(in3[45]), .Z(sumout[45]) );
  NBUFFX2 U3 ( .INP(in3[44]), .Z(sumout[44]) );
  NBUFFX2 U4 ( .INP(in3[43]), .Z(sumout[43]) );
  NBUFFX2 U5 ( .INP(in3[42]), .Z(sumout[42]) );
  NBUFFX2 U6 ( .INP(in3[37]), .Z(sumout[37]) );
  NBUFFX2 U7 ( .INP(in3[35]), .Z(sumout[35]) );
  NBUFFX2 U8 ( .INP(in3[33]), .Z(sumout[33]) );
  NBUFFX2 U9 ( .INP(in3[41]), .Z(sumout[41]) );
  NBUFFX2 U10 ( .INP(in3[40]), .Z(sumout[40]) );
  NBUFFX2 U11 ( .INP(in3[39]), .Z(sumout[39]) );
  NBUFFX2 U12 ( .INP(in3[38]), .Z(sumout[38]) );
  NBUFFX2 U13 ( .INP(in3[36]), .Z(sumout[36]) );
  NBUFFX2 U14 ( .INP(in3[34]), .Z(sumout[34]) );
  NBUFFX2 U15 ( .INP(in3[32]), .Z(sumout[32]) );
  AND2X1 U16 ( .IN1(in2[3]), .IN2(in1[3]), .Q(cout[3]) );
  AND2X1 U17 ( .IN1(in2[4]), .IN2(in1[4]), .Q(cout[4]) );
  NOR2X0 U18 ( .IN1(in2[4]), .IN2(in1[4]), .QN(n16) );
  NOR2X0 U19 ( .IN1(n16), .IN2(cout[4]), .QN(sumout[4]) );
  AND2X1 U20 ( .IN1(in2[5]), .IN2(in1[5]), .Q(cout[5]) );
  NOR2X0 U21 ( .IN1(in2[5]), .IN2(in1[5]), .QN(n17) );
  NOR2X0 U22 ( .IN1(n17), .IN2(cout[5]), .QN(sumout[5]) );
  AND2X1 U23 ( .IN1(in2[6]), .IN2(in1[6]), .Q(cout[6]) );
  NOR2X0 U24 ( .IN1(in2[6]), .IN2(in1[6]), .QN(n18) );
  NOR2X0 U25 ( .IN1(n18), .IN2(cout[6]), .QN(sumout[6]) );
  AND2X1 U26 ( .IN1(in2[7]), .IN2(in1[7]), .Q(cout[7]) );
  NOR2X0 U27 ( .IN1(in2[7]), .IN2(in1[7]), .QN(n19) );
  NOR2X0 U28 ( .IN1(n19), .IN2(cout[7]), .QN(sumout[7]) );
  AND2X1 U29 ( .IN1(in2[8]), .IN2(in1[8]), .Q(cout[8]) );
  NOR2X0 U30 ( .IN1(in2[8]), .IN2(in1[8]), .QN(n20) );
  NOR2X0 U31 ( .IN1(n20), .IN2(cout[8]), .QN(sumout[8]) );
  AND2X1 U32 ( .IN1(in2[9]), .IN2(in1[9]), .Q(cout[9]) );
  NOR2X0 U33 ( .IN1(in2[9]), .IN2(in1[9]), .QN(n21) );
  NOR2X0 U34 ( .IN1(n21), .IN2(cout[9]), .QN(sumout[9]) );
  AND2X1 U35 ( .IN1(in2[10]), .IN2(in1[10]), .Q(cout[10]) );
  NOR2X0 U36 ( .IN1(in2[10]), .IN2(in1[10]), .QN(n22) );
  NOR2X0 U37 ( .IN1(n22), .IN2(cout[10]), .QN(sumout[10]) );
  AND2X1 U38 ( .IN1(in2[11]), .IN2(in1[11]), .Q(cout[11]) );
  NOR2X0 U39 ( .IN1(in2[11]), .IN2(in1[11]), .QN(n23) );
  NOR2X0 U40 ( .IN1(n23), .IN2(cout[11]), .QN(sumout[11]) );
  AND2X1 U41 ( .IN1(in2[12]), .IN2(in1[12]), .Q(cout[12]) );
  NOR2X0 U42 ( .IN1(in2[12]), .IN2(in1[12]), .QN(n24) );
  NOR2X0 U43 ( .IN1(n24), .IN2(cout[12]), .QN(sumout[12]) );
  AND2X1 U44 ( .IN1(in2[13]), .IN2(in1[13]), .Q(cout[13]) );
  NOR2X0 U45 ( .IN1(in2[13]), .IN2(in1[13]), .QN(n25) );
  NOR2X0 U46 ( .IN1(n25), .IN2(cout[13]), .QN(sumout[13]) );
  AND2X1 U47 ( .IN1(in2[14]), .IN2(in1[14]), .Q(cout[14]) );
  NOR2X0 U48 ( .IN1(in2[14]), .IN2(in1[14]), .QN(n26) );
  NOR2X0 U49 ( .IN1(n26), .IN2(cout[14]), .QN(sumout[14]) );
  AND2X1 U50 ( .IN1(in2[15]), .IN2(in1[15]), .Q(cout[15]) );
  NOR2X0 U51 ( .IN1(in2[15]), .IN2(in1[15]), .QN(n27) );
  NOR2X0 U52 ( .IN1(n27), .IN2(cout[15]), .QN(sumout[15]) );
  AND2X1 U53 ( .IN1(in2[16]), .IN2(in1[16]), .Q(cout[16]) );
  NOR2X0 U54 ( .IN1(in2[16]), .IN2(in1[16]), .QN(n28) );
  NOR2X0 U55 ( .IN1(n28), .IN2(cout[16]), .QN(sumout[16]) );
  AND2X1 U56 ( .IN1(in2[17]), .IN2(in1[17]), .Q(cout[17]) );
  NOR2X0 U57 ( .IN1(in2[17]), .IN2(in1[17]), .QN(n29) );
  NOR2X0 U58 ( .IN1(n29), .IN2(cout[17]), .QN(sumout[17]) );
  AND2X1 U59 ( .IN1(in2[18]), .IN2(in1[18]), .Q(cout[18]) );
  NOR2X0 U60 ( .IN1(in2[18]), .IN2(in1[18]), .QN(n30) );
  NOR2X0 U61 ( .IN1(n30), .IN2(cout[18]), .QN(sumout[18]) );
  AND2X1 U62 ( .IN1(in2[19]), .IN2(in1[19]), .Q(cout[19]) );
  NOR2X0 U63 ( .IN1(in2[19]), .IN2(in1[19]), .QN(n31) );
  NOR2X0 U64 ( .IN1(n31), .IN2(cout[19]), .QN(sumout[19]) );
  AND2X1 U65 ( .IN1(in2[20]), .IN2(in1[20]), .Q(cout[20]) );
  NOR2X0 U66 ( .IN1(in2[20]), .IN2(in1[20]), .QN(n32) );
  NOR2X0 U67 ( .IN1(n32), .IN2(cout[20]), .QN(sumout[20]) );
  AND2X1 U68 ( .IN1(in2[21]), .IN2(in1[21]), .Q(cout[21]) );
  NOR2X0 U69 ( .IN1(in2[21]), .IN2(in1[21]), .QN(n33) );
  NOR2X0 U70 ( .IN1(n33), .IN2(cout[21]), .QN(sumout[21]) );
  AND2X1 U71 ( .IN1(in2[22]), .IN2(in1[22]), .Q(cout[22]) );
  NOR2X0 U72 ( .IN1(in2[22]), .IN2(in1[22]), .QN(n34) );
  NOR2X0 U73 ( .IN1(n34), .IN2(cout[22]), .QN(sumout[22]) );
  AND2X1 U74 ( .IN1(in2[23]), .IN2(in1[23]), .Q(cout[23]) );
  NOR2X0 U75 ( .IN1(in2[23]), .IN2(in1[23]), .QN(n35) );
  NOR2X0 U76 ( .IN1(n35), .IN2(cout[23]), .QN(sumout[23]) );
  AND2X1 U77 ( .IN1(in2[31]), .IN2(in3[31]), .Q(cout[31]) );
  INVX0 U78 ( .INP(in2[31]), .ZN(n36) );
  MUX21X1 U79 ( .IN1(in2[31]), .IN2(n36), .S(in3[31]), .Q(sumout[31]) );
  FADDX1 U80 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U81 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U82 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U83 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U84 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U85 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U86 ( .A(in1[30]), .B(in3[30]), .CI(n36), .CO(cout[30]), .S(
        sumout[30]) );
endmodule


module csa51squ_81 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n3, n4, n5, n6, n7;

  NBUFFX2 U1 ( .INP(in1[18]), .Z(sumout[18]) );
  NBUFFX2 U2 ( .INP(in1[19]), .Z(sumout[19]) );
  AND2X1 U3 ( .IN1(in2[20]), .IN2(in1[20]), .Q(cout[20]) );
  NOR2X0 U4 ( .IN1(in2[20]), .IN2(in1[20]), .QN(n3) );
  NOR2X0 U5 ( .IN1(n3), .IN2(cout[20]), .QN(sumout[20]) );
  AND2X1 U6 ( .IN1(in2[21]), .IN2(in1[21]), .Q(cout[21]) );
  NOR2X0 U7 ( .IN1(in2[21]), .IN2(in1[21]), .QN(n4) );
  NOR2X0 U8 ( .IN1(n4), .IN2(cout[21]), .QN(sumout[21]) );
  AND2X1 U9 ( .IN1(in2[46]), .IN2(in3[46]), .Q(cout[46]) );
  NOR2X0 U10 ( .IN1(in2[46]), .IN2(in3[46]), .QN(n5) );
  NOR2X0 U11 ( .IN1(n5), .IN2(cout[46]), .QN(sumout[46]) );
  INVX0 U12 ( .INP(in2[46]), .ZN(n6) );
  MUX21X1 U13 ( .IN1(n6), .IN2(in2[46]), .S(in3[47]), .Q(sumout[47]) );
  INVX0 U14 ( .INP(in1[44]), .ZN(n7) );
  FADDX1 U15 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U16 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U17 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U18 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U19 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U20 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U21 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U22 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U23 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U24 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U25 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
  FADDX1 U26 ( .A(in1[33]), .B(in2[33]), .CI(in3[33]), .CO(cout[33]), .S(
        sumout[33]) );
  FADDX1 U27 ( .A(in1[34]), .B(in2[34]), .CI(in3[34]), .CO(cout[34]), .S(
        sumout[34]) );
  FADDX1 U28 ( .A(in1[35]), .B(in2[35]), .CI(in3[35]), .CO(cout[35]), .S(
        sumout[35]) );
  FADDX1 U29 ( .A(in1[36]), .B(in2[36]), .CI(in3[36]), .CO(cout[36]), .S(
        sumout[36]) );
  FADDX1 U30 ( .A(in1[37]), .B(in2[37]), .CI(in3[37]), .CO(cout[37]), .S(
        sumout[37]) );
  FADDX1 U31 ( .A(in1[38]), .B(in2[38]), .CI(in3[38]), .CO(cout[38]), .S(
        sumout[38]) );
  FADDX1 U32 ( .A(in1[39]), .B(in2[39]), .CI(in3[39]), .CO(cout[39]), .S(
        sumout[39]) );
  FADDX1 U33 ( .A(in1[40]), .B(in2[40]), .CI(in3[40]), .CO(cout[40]), .S(
        sumout[40]) );
  FADDX1 U34 ( .A(in1[41]), .B(in2[41]), .CI(in3[41]), .CO(cout[41]), .S(
        sumout[41]) );
  FADDX1 U35 ( .A(in1[42]), .B(in2[42]), .CI(in3[42]), .CO(cout[42]), .S(
        sumout[42]) );
  FADDX1 U36 ( .A(in1[43]), .B(in2[43]), .CI(in3[43]), .CO(cout[43]), .S(
        sumout[43]) );
  FADDX1 U37 ( .A(in1[44]), .B(in2[44]), .CI(in3[44]), .CO(cout[44]), .S(
        sumout[44]) );
  FADDX1 U38 ( .A(in2[45]), .B(in3[45]), .CI(n7), .CO(cout[45]), .S(sumout[45]) );
endmodule


module csa51squ_82 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n4, n5, n6, n7, n8;

  NBUFFX2 U1 ( .INP(in1[12]), .Z(sumout[12]) );
  NBUFFX2 U2 ( .INP(in1[13]), .Z(sumout[13]) );
  NBUFFX2 U3 ( .INP(in3[42]), .Z(sumout[42]) );
  AND2X1 U4 ( .IN1(in2[14]), .IN2(in1[14]), .Q(cout[14]) );
  NOR2X0 U5 ( .IN1(in2[14]), .IN2(in1[14]), .QN(n4) );
  NOR2X0 U6 ( .IN1(n4), .IN2(cout[14]), .QN(sumout[14]) );
  AND2X1 U7 ( .IN1(in2[15]), .IN2(in1[15]), .Q(cout[15]) );
  NOR2X0 U8 ( .IN1(in2[15]), .IN2(in1[15]), .QN(n5) );
  NOR2X0 U9 ( .IN1(n5), .IN2(cout[15]), .QN(sumout[15]) );
  AND2X1 U10 ( .IN1(in2[40]), .IN2(in3[40]), .Q(cout[40]) );
  NOR2X0 U11 ( .IN1(in2[40]), .IN2(in3[40]), .QN(n6) );
  NOR2X0 U12 ( .IN1(n6), .IN2(cout[40]), .QN(sumout[40]) );
  INVX0 U13 ( .INP(in3[41]), .ZN(n7) );
  NOR2X0 U14 ( .IN1(in2[40]), .IN2(n7), .QN(cout[41]) );
  MUX21X1 U15 ( .IN1(n7), .IN2(in3[41]), .S(in2[40]), .Q(sumout[41]) );
  INVX0 U16 ( .INP(in1[38]), .ZN(n8) );
  FADDX1 U17 ( .A(in1[16]), .B(in2[16]), .CI(in3[16]), .CO(cout[16]), .S(
        sumout[16]) );
  FADDX1 U18 ( .A(in1[17]), .B(in2[17]), .CI(in3[17]), .CO(cout[17]), .S(
        sumout[17]) );
  FADDX1 U19 ( .A(in1[18]), .B(in2[18]), .CI(in3[18]), .CO(cout[18]), .S(
        sumout[18]) );
  FADDX1 U20 ( .A(in1[19]), .B(in2[19]), .CI(in3[19]), .CO(cout[19]), .S(
        sumout[19]) );
  FADDX1 U21 ( .A(in1[20]), .B(in2[20]), .CI(in3[20]), .CO(cout[20]), .S(
        sumout[20]) );
  FADDX1 U22 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U23 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U24 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U25 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U26 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U27 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U28 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U29 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U30 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U31 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U32 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U33 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
  FADDX1 U34 ( .A(in1[33]), .B(in2[33]), .CI(in3[33]), .CO(cout[33]), .S(
        sumout[33]) );
  FADDX1 U35 ( .A(in1[34]), .B(in2[34]), .CI(in3[34]), .CO(cout[34]), .S(
        sumout[34]) );
  FADDX1 U36 ( .A(in1[35]), .B(in2[35]), .CI(in3[35]), .CO(cout[35]), .S(
        sumout[35]) );
  FADDX1 U37 ( .A(in1[36]), .B(in2[36]), .CI(in3[36]), .CO(cout[36]), .S(
        sumout[36]) );
  FADDX1 U38 ( .A(in1[37]), .B(in2[37]), .CI(in3[37]), .CO(cout[37]), .S(
        sumout[37]) );
  FADDX1 U39 ( .A(in1[38]), .B(in2[38]), .CI(in3[38]), .CO(cout[38]), .S(
        sumout[38]) );
  FADDX1 U40 ( .A(in2[39]), .B(in3[39]), .CI(n8), .CO(cout[39]), .S(sumout[39]) );
endmodule


module csa51squ_83 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n4, n5, n6, n7, n8;

  NBUFFX2 U1 ( .INP(in1[6]), .Z(sumout[6]) );
  NBUFFX2 U2 ( .INP(in1[7]), .Z(sumout[7]) );
  NBUFFX2 U3 ( .INP(in3[37]), .Z(sumout[37]) );
  AND2X1 U4 ( .IN1(in2[8]), .IN2(in1[8]), .Q(cout[8]) );
  NOR2X0 U5 ( .IN1(in2[8]), .IN2(in1[8]), .QN(n4) );
  NOR2X0 U6 ( .IN1(n4), .IN2(cout[8]), .QN(sumout[8]) );
  AND2X1 U7 ( .IN1(in2[9]), .IN2(in1[9]), .Q(cout[9]) );
  NOR2X0 U8 ( .IN1(in2[9]), .IN2(in1[9]), .QN(n5) );
  NOR2X0 U9 ( .IN1(n5), .IN2(cout[9]), .QN(sumout[9]) );
  AND2X1 U10 ( .IN1(in2[34]), .IN2(in3[34]), .Q(cout[34]) );
  NOR2X0 U11 ( .IN1(in2[34]), .IN2(in3[34]), .QN(n6) );
  NOR2X0 U12 ( .IN1(n6), .IN2(cout[34]), .QN(sumout[34]) );
  INVX0 U13 ( .INP(in3[35]), .ZN(n7) );
  NOR2X0 U14 ( .IN1(in2[34]), .IN2(n7), .QN(cout[35]) );
  MUX21X1 U15 ( .IN1(n7), .IN2(in3[35]), .S(in2[34]), .Q(sumout[35]) );
  INVX0 U16 ( .INP(in1[32]), .ZN(n8) );
  FADDX1 U17 ( .A(in1[10]), .B(in2[10]), .CI(in3[10]), .CO(cout[10]), .S(
        sumout[10]) );
  FADDX1 U18 ( .A(in1[11]), .B(in2[11]), .CI(in3[11]), .CO(cout[11]), .S(
        sumout[11]) );
  FADDX1 U19 ( .A(in1[12]), .B(in2[12]), .CI(in3[12]), .CO(cout[12]), .S(
        sumout[12]) );
  FADDX1 U20 ( .A(in1[13]), .B(in2[13]), .CI(in3[13]), .CO(cout[13]), .S(
        sumout[13]) );
  FADDX1 U21 ( .A(in1[14]), .B(in2[14]), .CI(in3[14]), .CO(cout[14]), .S(
        sumout[14]) );
  FADDX1 U22 ( .A(in1[15]), .B(in2[15]), .CI(in3[15]), .CO(cout[15]), .S(
        sumout[15]) );
  FADDX1 U23 ( .A(in1[16]), .B(in2[16]), .CI(in3[16]), .CO(cout[16]), .S(
        sumout[16]) );
  FADDX1 U24 ( .A(in1[17]), .B(in2[17]), .CI(in3[17]), .CO(cout[17]), .S(
        sumout[17]) );
  FADDX1 U25 ( .A(in1[18]), .B(in2[18]), .CI(in3[18]), .CO(cout[18]), .S(
        sumout[18]) );
  FADDX1 U26 ( .A(in1[19]), .B(in2[19]), .CI(in3[19]), .CO(cout[19]), .S(
        sumout[19]) );
  FADDX1 U27 ( .A(in1[20]), .B(in2[20]), .CI(in3[20]), .CO(cout[20]), .S(
        sumout[20]) );
  FADDX1 U28 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U29 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U30 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U31 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U32 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U33 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U34 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U35 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U36 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U37 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U38 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U39 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
  FADDX1 U40 ( .A(in2[33]), .B(in3[33]), .CI(n8), .CO(cout[33]), .S(sumout[33]) );
endmodule


module booth27_79 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;


  NBUFFX2 U3 ( .INP(in2[22]), .Z(out1[22]) );
  NBUFFX2 U4 ( .INP(in2[21]), .Z(out1[21]) );
  NBUFFX2 U5 ( .INP(in2[20]), .Z(out1[20]) );
  NBUFFX2 U6 ( .INP(in2[0]), .Z(out1[0]) );
  NBUFFX2 U7 ( .INP(in2[19]), .Z(out1[19]) );
  NBUFFX2 U8 ( .INP(in2[18]), .Z(out1[18]) );
  NBUFFX2 U9 ( .INP(in2[1]), .Z(out1[1]) );
  NBUFFX2 U10 ( .INP(in2[5]), .Z(out1[5]) );
  NBUFFX2 U11 ( .INP(in2[3]), .Z(out1[3]) );
  NBUFFX2 U12 ( .INP(in2[13]), .Z(out1[13]) );
  NBUFFX2 U13 ( .INP(in2[11]), .Z(out1[11]) );
  NBUFFX2 U14 ( .INP(in2[9]), .Z(out1[9]) );
  NBUFFX2 U15 ( .INP(in2[7]), .Z(out1[7]) );
  NBUFFX2 U16 ( .INP(in2[17]), .Z(out1[17]) );
  NBUFFX2 U17 ( .INP(in2[16]), .Z(out1[16]) );
  NBUFFX2 U18 ( .INP(in2[15]), .Z(out1[15]) );
  NBUFFX2 U19 ( .INP(in2[14]), .Z(out1[14]) );
  NBUFFX2 U20 ( .INP(in2[12]), .Z(out1[12]) );
  NBUFFX2 U21 ( .INP(in2[10]), .Z(out1[10]) );
  NBUFFX2 U22 ( .INP(in2[8]), .Z(out1[8]) );
  NBUFFX2 U23 ( .INP(in2[6]), .Z(out1[6]) );
  NBUFFX2 U24 ( .INP(in2[4]), .Z(out1[4]) );
  NBUFFX2 U25 ( .INP(in2[2]), .Z(out1[2]) );
endmodule


module booth27_80 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76;

  NAND2X0 U3 ( .IN1(n1), .IN2(n2), .QN(n8) );
  NAND2X0 U4 ( .IN1(n16), .IN2(in2[4]), .QN(n17) );
  NAND2X0 U5 ( .IN1(n19), .IN2(in2[5]), .QN(n20) );
  NAND2X0 U6 ( .IN1(n22), .IN2(in2[6]), .QN(n23) );
  NAND2X0 U7 ( .IN1(n25), .IN2(in2[7]), .QN(n26) );
  NAND2X0 U8 ( .IN1(n28), .IN2(in2[8]), .QN(n29) );
  NAND2X0 U9 ( .IN1(n31), .IN2(in2[9]), .QN(n32) );
  NAND2X0 U10 ( .IN1(n34), .IN2(in2[10]), .QN(n35) );
  NAND2X0 U11 ( .IN1(n37), .IN2(in2[11]), .QN(n38) );
  NAND2X0 U12 ( .IN1(n40), .IN2(in2[12]), .QN(n41) );
  NAND2X0 U13 ( .IN1(n43), .IN2(in2[13]), .QN(n44) );
  NAND2X0 U14 ( .IN1(n46), .IN2(in2[14]), .QN(n47) );
  NAND2X0 U15 ( .IN1(n49), .IN2(in2[15]), .QN(n50) );
  NAND2X0 U16 ( .IN1(n52), .IN2(in2[16]), .QN(n53) );
  NAND2X0 U17 ( .IN1(n55), .IN2(in2[17]), .QN(n56) );
  NAND2X0 U18 ( .IN1(n7), .IN2(n15), .QN(out1[1]) );
  NAND2X0 U19 ( .IN1(n10), .IN2(n9), .QN(out1[2]) );
  NAND2X0 U20 ( .IN1(n58), .IN2(in2[18]), .QN(n59) );
  NAND2X0 U21 ( .IN1(n61), .IN2(in2[19]), .QN(n62) );
  NOR2X0 U22 ( .IN1(in1[1]), .IN2(in1[0]), .QN(n71) );
  INVX0 U23 ( .INP(in2[1]), .ZN(n2) );
  INVX0 U24 ( .INP(in2[0]), .ZN(n1) );
  INVX0 U25 ( .INP(in2[3]), .ZN(n3) );
  INVX0 U26 ( .INP(in2[21]), .ZN(n4) );
  INVX0 U27 ( .INP(in2[22]), .ZN(n5) );
  INVX0 U28 ( .INP(in1[1]), .ZN(n6) );
  MUX21X1 U29 ( .IN1(in1[1]), .IN2(n6), .S(in1[0]), .Q(n74) );
  INVX0 U30 ( .INP(n74), .ZN(n76) );
  AO221X1 U31 ( .IN1(in2[0]), .IN2(in2[1]), .IN3(n1), .IN4(n2), .IN5(n76), .Q(
        n7) );
  NAND2X0 U32 ( .IN1(n71), .IN2(in2[0]), .QN(n15) );
  MUX21X1 U33 ( .IN1(n2), .IN2(n8), .S(in2[2]), .Q(n12) );
  AO221X1 U34 ( .IN1(n12), .IN2(in2[2]), .IN3(n12), .IN4(n1), .IN5(n76), .Q(
        n10) );
  INVX0 U35 ( .INP(n71), .ZN(n13) );
  AO221X1 U36 ( .IN1(in2[0]), .IN2(in2[1]), .IN3(n1), .IN4(n2), .IN5(n13), .Q(
        n9) );
  NOR3X0 U37 ( .IN1(in2[0]), .IN2(in2[2]), .IN3(in2[1]), .QN(n11) );
  OR4X1 U38 ( .IN1(in2[3]), .IN2(in2[0]), .IN3(in2[2]), .IN4(in2[1]), .Q(n16)
         );
  OA21X1 U39 ( .IN1(n11), .IN2(n3), .IN3(n16), .Q(n18) );
  INVX0 U40 ( .INP(n18), .ZN(n14) );
  OAI222X1 U41 ( .IN1(n15), .IN2(in2[2]), .IN3(n14), .IN4(n76), .IN5(n13), 
        .IN6(n12), .QN(out1[3]) );
  OR2X1 U42 ( .IN1(in2[4]), .IN2(n16), .Q(n19) );
  AND2X1 U43 ( .IN1(n19), .IN2(n17), .Q(n21) );
  AO22X1 U44 ( .IN1(n71), .IN2(n18), .IN3(n21), .IN4(n74), .Q(out1[4]) );
  OR2X1 U45 ( .IN1(in2[5]), .IN2(n19), .Q(n22) );
  AND2X1 U46 ( .IN1(n22), .IN2(n20), .Q(n24) );
  AO22X1 U47 ( .IN1(n71), .IN2(n21), .IN3(n24), .IN4(n74), .Q(out1[5]) );
  OR2X1 U48 ( .IN1(in2[6]), .IN2(n22), .Q(n25) );
  AND2X1 U49 ( .IN1(n25), .IN2(n23), .Q(n27) );
  AO22X1 U50 ( .IN1(n71), .IN2(n24), .IN3(n27), .IN4(n74), .Q(out1[6]) );
  OR2X1 U51 ( .IN1(in2[7]), .IN2(n25), .Q(n28) );
  AND2X1 U52 ( .IN1(n28), .IN2(n26), .Q(n30) );
  AO22X1 U53 ( .IN1(n71), .IN2(n27), .IN3(n30), .IN4(n74), .Q(out1[7]) );
  OR2X1 U54 ( .IN1(in2[8]), .IN2(n28), .Q(n31) );
  AND2X1 U55 ( .IN1(n31), .IN2(n29), .Q(n33) );
  AO22X1 U56 ( .IN1(n71), .IN2(n30), .IN3(n33), .IN4(n74), .Q(out1[8]) );
  OR2X1 U57 ( .IN1(in2[9]), .IN2(n31), .Q(n34) );
  AND2X1 U58 ( .IN1(n34), .IN2(n32), .Q(n36) );
  AO22X1 U59 ( .IN1(n71), .IN2(n33), .IN3(n36), .IN4(n74), .Q(out1[9]) );
  OR2X1 U60 ( .IN1(in2[10]), .IN2(n34), .Q(n37) );
  AND2X1 U61 ( .IN1(n37), .IN2(n35), .Q(n39) );
  AO22X1 U62 ( .IN1(n71), .IN2(n36), .IN3(n39), .IN4(n74), .Q(out1[10]) );
  OR2X1 U63 ( .IN1(in2[11]), .IN2(n37), .Q(n40) );
  AND2X1 U64 ( .IN1(n40), .IN2(n38), .Q(n42) );
  AO22X1 U65 ( .IN1(n71), .IN2(n39), .IN3(n42), .IN4(n74), .Q(out1[11]) );
  OR2X1 U66 ( .IN1(in2[12]), .IN2(n40), .Q(n43) );
  AND2X1 U67 ( .IN1(n43), .IN2(n41), .Q(n45) );
  AO22X1 U68 ( .IN1(n71), .IN2(n42), .IN3(n45), .IN4(n74), .Q(out1[12]) );
  OR2X1 U69 ( .IN1(in2[13]), .IN2(n43), .Q(n46) );
  AND2X1 U70 ( .IN1(n46), .IN2(n44), .Q(n48) );
  AO22X1 U71 ( .IN1(n71), .IN2(n45), .IN3(n48), .IN4(n74), .Q(out1[13]) );
  OR2X1 U72 ( .IN1(in2[14]), .IN2(n46), .Q(n49) );
  AND2X1 U73 ( .IN1(n49), .IN2(n47), .Q(n51) );
  AO22X1 U74 ( .IN1(n71), .IN2(n48), .IN3(n51), .IN4(n74), .Q(out1[14]) );
  OR2X1 U75 ( .IN1(in2[15]), .IN2(n49), .Q(n52) );
  AND2X1 U76 ( .IN1(n52), .IN2(n50), .Q(n54) );
  AO22X1 U77 ( .IN1(n71), .IN2(n51), .IN3(n54), .IN4(n74), .Q(out1[15]) );
  OR2X1 U78 ( .IN1(in2[16]), .IN2(n52), .Q(n55) );
  AND2X1 U79 ( .IN1(n55), .IN2(n53), .Q(n57) );
  AO22X1 U80 ( .IN1(n71), .IN2(n54), .IN3(n57), .IN4(n74), .Q(out1[16]) );
  OR2X1 U81 ( .IN1(in2[17]), .IN2(n55), .Q(n58) );
  AND2X1 U82 ( .IN1(n58), .IN2(n56), .Q(n60) );
  AO22X1 U83 ( .IN1(n71), .IN2(n57), .IN3(n60), .IN4(n74), .Q(out1[17]) );
  OR2X1 U84 ( .IN1(in2[18]), .IN2(n58), .Q(n61) );
  AND2X1 U85 ( .IN1(n61), .IN2(n59), .Q(n63) );
  AO22X1 U86 ( .IN1(n71), .IN2(n60), .IN3(n63), .IN4(n74), .Q(out1[18]) );
  OR2X1 U87 ( .IN1(in2[19]), .IN2(n61), .Q(n64) );
  AND2X1 U88 ( .IN1(n64), .IN2(n62), .Q(n65) );
  AO22X1 U89 ( .IN1(n71), .IN2(n63), .IN3(n65), .IN4(n74), .Q(out1[19]) );
  NOR2X0 U90 ( .IN1(in2[20]), .IN2(n64), .QN(n72) );
  AOI21X1 U91 ( .IN1(in2[20]), .IN2(n64), .IN3(n72), .QN(n66) );
  AO22X1 U92 ( .IN1(n71), .IN2(n65), .IN3(n66), .IN4(n74), .Q(out1[20]) );
  MUX21X1 U93 ( .IN1(n4), .IN2(in2[21]), .S(n72), .Q(n69) );
  AO22X1 U94 ( .IN1(n71), .IN2(n66), .IN3(n69), .IN4(n74), .Q(out1[21]) );
  INVX0 U95 ( .INP(n72), .ZN(n67) );
  NOR2X0 U96 ( .IN1(in2[21]), .IN2(n67), .QN(n70) );
  MUX21X1 U97 ( .IN1(n5), .IN2(in2[22]), .S(n70), .Q(n68) );
  AO22X1 U98 ( .IN1(n71), .IN2(n69), .IN3(n68), .IN4(n74), .Q(out1[22]) );
  MUX21X1 U99 ( .IN1(n71), .IN2(n74), .S(n70), .Q(n73) );
  AND3X1 U100 ( .IN1(n72), .IN2(n71), .IN3(n4), .Q(n75) );
  MUX21X1 U101 ( .IN1(n73), .IN2(n75), .S(in2[22]), .Q(out1[23]) );
  AO21X1 U102 ( .IN1(n75), .IN2(n5), .IN3(n74), .Q(out1[24]) );
  NAND2X0 U103 ( .IN1(in1[1]), .IN2(in1[0]), .QN(out1[25]) );
  NOR2X0 U104 ( .IN1(n76), .IN2(n1), .QN(out1[0]) );
endmodule


module booth27_81 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n19), .IN2(n25), .QN(n24) );
  NAND2X0 U4 ( .IN1(n28), .IN2(n33), .QN(n32) );
  NAND2X0 U5 ( .IN1(n37), .IN2(n42), .QN(n41) );
  NAND2X0 U6 ( .IN1(n46), .IN2(n51), .QN(n50) );
  NAND2X0 U7 ( .IN1(n55), .IN2(n60), .QN(n59) );
  NAND2X0 U8 ( .IN1(n64), .IN2(n71), .QN(n77) );
  NAND2X0 U9 ( .IN1(n81), .IN2(n7), .QN(n89) );
  NAND2X0 U10 ( .IN1(n93), .IN2(n9), .QN(n101) );
  NAND2X0 U11 ( .IN1(n105), .IN2(n11), .QN(n114) );
  NAND2X0 U12 ( .IN1(n21), .IN2(n132), .QN(n4) );
  NAND2X0 U13 ( .IN1(in1[2]), .IN2(n77), .QN(n70) );
  NAND2X0 U14 ( .IN1(n69), .IN2(n132), .QN(n74) );
  NAND2X0 U15 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U16 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U17 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U18 ( .IN1(n118), .IN2(n13), .QN(n125) );
  NAND2X0 U19 ( .IN1(n141), .IN2(n130), .QN(n18) );
  NAND2X0 U20 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NAND2X0 U21 ( .IN1(n27), .IN2(n26), .QN(out1[3]) );
  NAND2X0 U22 ( .IN1(n31), .IN2(n30), .QN(out1[4]) );
  NAND2X0 U23 ( .IN1(n36), .IN2(n35), .QN(out1[5]) );
  NAND2X0 U24 ( .IN1(n40), .IN2(n39), .QN(out1[6]) );
  NAND2X0 U25 ( .IN1(n45), .IN2(n44), .QN(out1[7]) );
  NAND2X0 U26 ( .IN1(n49), .IN2(n48), .QN(out1[8]) );
  NAND2X0 U27 ( .IN1(n54), .IN2(n53), .QN(out1[9]) );
  NAND2X0 U28 ( .IN1(n58), .IN2(n57), .QN(out1[10]) );
  NAND2X0 U29 ( .IN1(n63), .IN2(n62), .QN(out1[11]) );
  NAND2X0 U30 ( .IN1(n68), .IN2(n67), .QN(out1[12]) );
  NAND2X0 U31 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U32 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U33 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U34 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U35 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U36 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U37 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U38 ( .IN1(n17), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U39 ( .IN1(in1[2]), .IN2(n16), .QN(n17) );
  NOR2X0 U40 ( .IN1(n22), .IN2(n20), .QN(n3) );
  NOR2X0 U41 ( .IN1(n142), .IN2(n15), .QN(n1) );
  NOR2X0 U42 ( .IN1(n142), .IN2(n111), .QN(n138) );
  INVX0 U43 ( .INP(n130), .ZN(n137) );
  INVX0 U44 ( .INP(n132), .ZN(n141) );
  NOR3X0 U45 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  NAND3X0 U46 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  MUX21X1 U47 ( .IN1(n16), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  INVX0 U48 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U49 ( .INP(in2[13]), .ZN(n6) );
  INVX0 U50 ( .INP(in2[14]), .ZN(n7) );
  INVX0 U51 ( .INP(in2[15]), .ZN(n8) );
  INVX0 U52 ( .INP(in2[16]), .ZN(n9) );
  INVX0 U53 ( .INP(in2[17]), .ZN(n10) );
  INVX0 U54 ( .INP(in2[18]), .ZN(n11) );
  INVX0 U55 ( .INP(in2[19]), .ZN(n12) );
  INVX0 U56 ( .INP(in2[20]), .ZN(n13) );
  INVX0 U57 ( .INP(in2[21]), .ZN(n14) );
  INVX0 U58 ( .INP(in2[22]), .ZN(n15) );
  INVX0 U59 ( .INP(in1[1]), .ZN(n16) );
  INVX0 U60 ( .INP(in1[2]), .ZN(n111) );
  INVX0 U61 ( .INP(n138), .ZN(n140) );
  NOR2X0 U62 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n19) );
  AOI21X1 U63 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n19), .QN(n21) );
  NOR2X0 U64 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U65 ( .IN1(n18), .IN2(in2[0]), .IN3(n138), .IN4(n21), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U66 ( .INP(n133), .ZN(n66) );
  INVX0 U67 ( .INP(in2[2]), .ZN(n25) );
  NOR2X0 U68 ( .IN1(n66), .IN2(n25), .QN(n22) );
  OA21X1 U69 ( .IN1(n19), .IN2(n25), .IN3(n24), .Q(n23) );
  AO22X1 U70 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n23), .Q(n20) );
  AOI22X1 U71 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n23), .QN(n27) );
  NOR2X0 U72 ( .IN1(in2[3]), .IN2(n24), .QN(n28) );
  AO21X1 U73 ( .IN1(in2[3]), .IN2(n24), .IN3(n28), .Q(n29) );
  OA22X1 U74 ( .IN1(n25), .IN2(n130), .IN3(n140), .IN4(n29), .Q(n26) );
  INVX0 U75 ( .INP(in2[4]), .ZN(n33) );
  OA21X1 U76 ( .IN1(n28), .IN2(n33), .IN3(n32), .Q(n34) );
  AOI22X1 U77 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n34), .QN(n31) );
  OA22X1 U78 ( .IN1(n66), .IN2(n33), .IN3(n141), .IN4(n29), .Q(n30) );
  NOR2X0 U79 ( .IN1(in2[5]), .IN2(n32), .QN(n37) );
  AO21X1 U80 ( .IN1(in2[5]), .IN2(n32), .IN3(n37), .Q(n38) );
  OA22X1 U81 ( .IN1(n33), .IN2(n130), .IN3(n140), .IN4(n38), .Q(n36) );
  AOI22X1 U82 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n34), .QN(n35) );
  INVX0 U83 ( .INP(in2[6]), .ZN(n42) );
  OA21X1 U84 ( .IN1(n37), .IN2(n42), .IN3(n41), .Q(n43) );
  AOI22X1 U85 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n43), .QN(n40) );
  OA22X1 U86 ( .IN1(n66), .IN2(n42), .IN3(n141), .IN4(n38), .Q(n39) );
  NOR2X0 U87 ( .IN1(in2[7]), .IN2(n41), .QN(n46) );
  AO21X1 U88 ( .IN1(in2[7]), .IN2(n41), .IN3(n46), .Q(n47) );
  OA22X1 U89 ( .IN1(n42), .IN2(n130), .IN3(n140), .IN4(n47), .Q(n45) );
  AOI22X1 U90 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n43), .QN(n44) );
  INVX0 U91 ( .INP(in2[8]), .ZN(n51) );
  OA21X1 U92 ( .IN1(n46), .IN2(n51), .IN3(n50), .Q(n52) );
  AOI22X1 U93 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n52), .QN(n49) );
  OA22X1 U94 ( .IN1(n66), .IN2(n51), .IN3(n141), .IN4(n47), .Q(n48) );
  NOR2X0 U95 ( .IN1(in2[9]), .IN2(n50), .QN(n55) );
  AO21X1 U96 ( .IN1(in2[9]), .IN2(n50), .IN3(n55), .Q(n56) );
  OA22X1 U97 ( .IN1(n51), .IN2(n130), .IN3(n140), .IN4(n56), .Q(n54) );
  AOI22X1 U98 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n52), .QN(n53) );
  INVX0 U99 ( .INP(in2[10]), .ZN(n60) );
  OA21X1 U100 ( .IN1(n55), .IN2(n60), .IN3(n59), .Q(n61) );
  AOI22X1 U101 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n61), .QN(n58) );
  OA22X1 U102 ( .IN1(n66), .IN2(n60), .IN3(n141), .IN4(n56), .Q(n57) );
  NOR2X0 U103 ( .IN1(in2[11]), .IN2(n59), .QN(n64) );
  AO21X1 U104 ( .IN1(in2[11]), .IN2(n59), .IN3(n64), .Q(n65) );
  OA22X1 U105 ( .IN1(n60), .IN2(n130), .IN3(n140), .IN4(n65), .Q(n63) );
  AOI22X1 U106 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n61), .QN(n62) );
  INVX0 U107 ( .INP(in2[12]), .ZN(n71) );
  OA21X1 U108 ( .IN1(n64), .IN2(n71), .IN3(n77), .Q(n69) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n69), .QN(n68) );
  OA22X1 U110 ( .IN1(n66), .IN2(n71), .IN3(n141), .IN4(n65), .Q(n67) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n6), .S(n70), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n71), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n7), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n6), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n6), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n8), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n7), .IN4(n85), .IN5(n84), .Q(
        out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n9), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n8), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n8), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n10), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n9), .IN4(n97), .IN5(n96), .Q(
        out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n11), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n10), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n10), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n12), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n11), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n13), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n12), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n12), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n14), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n13), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n15), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n14), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n14), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n15), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_82 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n28), .IN2(n33), .QN(n32) );
  NAND2X0 U4 ( .IN1(n37), .IN2(n42), .QN(n41) );
  NAND2X0 U5 ( .IN1(n46), .IN2(n51), .QN(n50) );
  NAND2X0 U6 ( .IN1(n55), .IN2(n60), .QN(n59) );
  NAND2X0 U7 ( .IN1(n19), .IN2(n25), .QN(n24) );
  NAND2X0 U8 ( .IN1(n64), .IN2(n71), .QN(n77) );
  NAND2X0 U9 ( .IN1(n81), .IN2(n7), .QN(n89) );
  NAND2X0 U10 ( .IN1(n93), .IN2(n9), .QN(n101) );
  NAND2X0 U11 ( .IN1(n105), .IN2(n11), .QN(n114) );
  NAND2X0 U12 ( .IN1(n118), .IN2(n13), .QN(n125) );
  NAND2X0 U13 ( .IN1(in1[2]), .IN2(n77), .QN(n70) );
  NAND2X0 U14 ( .IN1(n69), .IN2(n132), .QN(n74) );
  NAND2X0 U15 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U16 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U17 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U18 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U19 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U20 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U21 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U22 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NAND2X0 U23 ( .IN1(n21), .IN2(n132), .QN(n4) );
  NAND2X0 U24 ( .IN1(n27), .IN2(n26), .QN(out1[3]) );
  NAND2X0 U25 ( .IN1(n31), .IN2(n30), .QN(out1[4]) );
  NAND2X0 U26 ( .IN1(n36), .IN2(n35), .QN(out1[5]) );
  NAND2X0 U27 ( .IN1(n40), .IN2(n39), .QN(out1[6]) );
  NAND2X0 U28 ( .IN1(n45), .IN2(n44), .QN(out1[7]) );
  NAND2X0 U29 ( .IN1(n49), .IN2(n48), .QN(out1[8]) );
  NAND2X0 U30 ( .IN1(n54), .IN2(n53), .QN(out1[9]) );
  NAND2X0 U31 ( .IN1(n58), .IN2(n57), .QN(out1[10]) );
  NAND2X0 U32 ( .IN1(n63), .IN2(n62), .QN(out1[11]) );
  NAND2X0 U33 ( .IN1(n68), .IN2(n67), .QN(out1[12]) );
  NAND2X0 U34 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U35 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U36 ( .IN1(n141), .IN2(n130), .QN(n18) );
  NAND2X0 U37 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U38 ( .IN1(n17), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U39 ( .IN1(in1[2]), .IN2(n16), .QN(n17) );
  NOR2X0 U40 ( .IN1(n22), .IN2(n20), .QN(n3) );
  NOR2X0 U41 ( .IN1(n142), .IN2(n111), .QN(n138) );
  NOR2X0 U42 ( .IN1(n142), .IN2(n15), .QN(n1) );
  INVX0 U43 ( .INP(n130), .ZN(n137) );
  INVX0 U44 ( .INP(n132), .ZN(n141) );
  NOR3X0 U45 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  NAND3X0 U46 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  MUX21X1 U47 ( .IN1(n16), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  INVX0 U48 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U49 ( .INP(in2[13]), .ZN(n6) );
  INVX0 U50 ( .INP(in2[14]), .ZN(n7) );
  INVX0 U51 ( .INP(in2[15]), .ZN(n8) );
  INVX0 U52 ( .INP(in2[16]), .ZN(n9) );
  INVX0 U53 ( .INP(in2[17]), .ZN(n10) );
  INVX0 U54 ( .INP(in2[18]), .ZN(n11) );
  INVX0 U55 ( .INP(in2[19]), .ZN(n12) );
  INVX0 U56 ( .INP(in2[20]), .ZN(n13) );
  INVX0 U57 ( .INP(in2[21]), .ZN(n14) );
  INVX0 U58 ( .INP(in2[22]), .ZN(n15) );
  INVX0 U59 ( .INP(in1[1]), .ZN(n16) );
  INVX0 U60 ( .INP(in1[2]), .ZN(n111) );
  INVX0 U61 ( .INP(n138), .ZN(n140) );
  NOR2X0 U62 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n19) );
  AOI21X1 U63 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n19), .QN(n21) );
  NOR2X0 U64 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U65 ( .IN1(n18), .IN2(in2[0]), .IN3(n138), .IN4(n21), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U66 ( .INP(n133), .ZN(n66) );
  INVX0 U67 ( .INP(in2[2]), .ZN(n25) );
  NOR2X0 U68 ( .IN1(n66), .IN2(n25), .QN(n22) );
  OA21X1 U69 ( .IN1(n19), .IN2(n25), .IN3(n24), .Q(n23) );
  AO22X1 U70 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n23), .Q(n20) );
  AOI22X1 U71 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n23), .QN(n27) );
  NOR2X0 U72 ( .IN1(in2[3]), .IN2(n24), .QN(n28) );
  AO21X1 U73 ( .IN1(in2[3]), .IN2(n24), .IN3(n28), .Q(n29) );
  OA22X1 U74 ( .IN1(n25), .IN2(n130), .IN3(n140), .IN4(n29), .Q(n26) );
  INVX0 U75 ( .INP(in2[4]), .ZN(n33) );
  OA21X1 U76 ( .IN1(n28), .IN2(n33), .IN3(n32), .Q(n34) );
  AOI22X1 U77 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n34), .QN(n31) );
  OA22X1 U78 ( .IN1(n66), .IN2(n33), .IN3(n141), .IN4(n29), .Q(n30) );
  NOR2X0 U79 ( .IN1(in2[5]), .IN2(n32), .QN(n37) );
  AO21X1 U80 ( .IN1(in2[5]), .IN2(n32), .IN3(n37), .Q(n38) );
  OA22X1 U81 ( .IN1(n33), .IN2(n130), .IN3(n140), .IN4(n38), .Q(n36) );
  AOI22X1 U82 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n34), .QN(n35) );
  INVX0 U83 ( .INP(in2[6]), .ZN(n42) );
  OA21X1 U84 ( .IN1(n37), .IN2(n42), .IN3(n41), .Q(n43) );
  AOI22X1 U85 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n43), .QN(n40) );
  OA22X1 U86 ( .IN1(n66), .IN2(n42), .IN3(n141), .IN4(n38), .Q(n39) );
  NOR2X0 U87 ( .IN1(in2[7]), .IN2(n41), .QN(n46) );
  AO21X1 U88 ( .IN1(in2[7]), .IN2(n41), .IN3(n46), .Q(n47) );
  OA22X1 U89 ( .IN1(n42), .IN2(n130), .IN3(n140), .IN4(n47), .Q(n45) );
  AOI22X1 U90 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n43), .QN(n44) );
  INVX0 U91 ( .INP(in2[8]), .ZN(n51) );
  OA21X1 U92 ( .IN1(n46), .IN2(n51), .IN3(n50), .Q(n52) );
  AOI22X1 U93 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n52), .QN(n49) );
  OA22X1 U94 ( .IN1(n66), .IN2(n51), .IN3(n141), .IN4(n47), .Q(n48) );
  NOR2X0 U95 ( .IN1(in2[9]), .IN2(n50), .QN(n55) );
  AO21X1 U96 ( .IN1(in2[9]), .IN2(n50), .IN3(n55), .Q(n56) );
  OA22X1 U97 ( .IN1(n51), .IN2(n130), .IN3(n140), .IN4(n56), .Q(n54) );
  AOI22X1 U98 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n52), .QN(n53) );
  INVX0 U99 ( .INP(in2[10]), .ZN(n60) );
  OA21X1 U100 ( .IN1(n55), .IN2(n60), .IN3(n59), .Q(n61) );
  AOI22X1 U101 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n61), .QN(n58) );
  OA22X1 U102 ( .IN1(n66), .IN2(n60), .IN3(n141), .IN4(n56), .Q(n57) );
  NOR2X0 U103 ( .IN1(in2[11]), .IN2(n59), .QN(n64) );
  AO21X1 U104 ( .IN1(in2[11]), .IN2(n59), .IN3(n64), .Q(n65) );
  OA22X1 U105 ( .IN1(n60), .IN2(n130), .IN3(n140), .IN4(n65), .Q(n63) );
  AOI22X1 U106 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n61), .QN(n62) );
  INVX0 U107 ( .INP(in2[12]), .ZN(n71) );
  OA21X1 U108 ( .IN1(n64), .IN2(n71), .IN3(n77), .Q(n69) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n69), .QN(n68) );
  OA22X1 U110 ( .IN1(n66), .IN2(n71), .IN3(n141), .IN4(n65), .Q(n67) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n6), .S(n70), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n71), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n7), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n6), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n6), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n8), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n7), .IN4(n85), .IN5(n84), .Q(
        out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n9), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n8), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n8), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n10), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n9), .IN4(n97), .IN5(n96), .Q(
        out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n11), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n10), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n10), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n12), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n11), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n13), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n12), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n12), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n14), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n13), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n15), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n14), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n14), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n15), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_83 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n37), .IN2(n42), .QN(n41) );
  NAND2X0 U4 ( .IN1(n46), .IN2(n51), .QN(n50) );
  NAND2X0 U5 ( .IN1(n55), .IN2(n60), .QN(n59) );
  NAND2X0 U6 ( .IN1(n19), .IN2(n25), .QN(n24) );
  NAND2X0 U7 ( .IN1(n28), .IN2(n33), .QN(n32) );
  NAND2X0 U8 ( .IN1(n64), .IN2(n71), .QN(n77) );
  NAND2X0 U9 ( .IN1(n81), .IN2(n7), .QN(n89) );
  NAND2X0 U10 ( .IN1(n93), .IN2(n9), .QN(n101) );
  NAND2X0 U11 ( .IN1(in1[2]), .IN2(n77), .QN(n70) );
  NAND2X0 U12 ( .IN1(n69), .IN2(n132), .QN(n74) );
  NAND2X0 U13 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U14 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U15 ( .IN1(n105), .IN2(n11), .QN(n114) );
  NAND2X0 U16 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U17 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U18 ( .IN1(n21), .IN2(n132), .QN(n4) );
  NAND2X0 U19 ( .IN1(n141), .IN2(n130), .QN(n18) );
  NAND2X0 U20 ( .IN1(n36), .IN2(n35), .QN(out1[5]) );
  NAND2X0 U21 ( .IN1(n40), .IN2(n39), .QN(out1[6]) );
  NAND2X0 U22 ( .IN1(n45), .IN2(n44), .QN(out1[7]) );
  NAND2X0 U23 ( .IN1(n49), .IN2(n48), .QN(out1[8]) );
  NAND2X0 U24 ( .IN1(n54), .IN2(n53), .QN(out1[9]) );
  NAND2X0 U25 ( .IN1(n58), .IN2(n57), .QN(out1[10]) );
  NAND2X0 U26 ( .IN1(n63), .IN2(n62), .QN(out1[11]) );
  NAND2X0 U27 ( .IN1(n68), .IN2(n67), .QN(out1[12]) );
  NAND2X0 U28 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U29 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U30 ( .IN1(n118), .IN2(n13), .QN(n125) );
  NAND2X0 U31 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U32 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U33 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U34 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U35 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NAND2X0 U36 ( .IN1(n27), .IN2(n26), .QN(out1[3]) );
  NAND2X0 U37 ( .IN1(n31), .IN2(n30), .QN(out1[4]) );
  NAND2X0 U38 ( .IN1(n17), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U39 ( .IN1(in1[2]), .IN2(n16), .QN(n17) );
  NOR2X0 U40 ( .IN1(n22), .IN2(n20), .QN(n3) );
  NOR2X0 U41 ( .IN1(n142), .IN2(n15), .QN(n1) );
  INVX0 U42 ( .INP(n132), .ZN(n141) );
  INVX0 U43 ( .INP(n130), .ZN(n137) );
  NOR2X0 U44 ( .IN1(n142), .IN2(n111), .QN(n138) );
  MUX21X1 U45 ( .IN1(n16), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  NAND3X0 U46 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  NOR3X0 U47 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  INVX0 U48 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U49 ( .INP(in2[13]), .ZN(n6) );
  INVX0 U50 ( .INP(in2[14]), .ZN(n7) );
  INVX0 U51 ( .INP(in2[15]), .ZN(n8) );
  INVX0 U52 ( .INP(in2[16]), .ZN(n9) );
  INVX0 U53 ( .INP(in2[17]), .ZN(n10) );
  INVX0 U54 ( .INP(in2[18]), .ZN(n11) );
  INVX0 U55 ( .INP(in2[19]), .ZN(n12) );
  INVX0 U56 ( .INP(in2[20]), .ZN(n13) );
  INVX0 U57 ( .INP(in2[21]), .ZN(n14) );
  INVX0 U58 ( .INP(in2[22]), .ZN(n15) );
  INVX0 U59 ( .INP(in1[1]), .ZN(n16) );
  INVX0 U60 ( .INP(in1[2]), .ZN(n111) );
  INVX0 U61 ( .INP(n138), .ZN(n140) );
  NOR2X0 U62 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n19) );
  AOI21X1 U63 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n19), .QN(n21) );
  NOR2X0 U64 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U65 ( .IN1(n18), .IN2(in2[0]), .IN3(n138), .IN4(n21), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U66 ( .INP(n133), .ZN(n66) );
  INVX0 U67 ( .INP(in2[2]), .ZN(n25) );
  NOR2X0 U68 ( .IN1(n66), .IN2(n25), .QN(n22) );
  OA21X1 U69 ( .IN1(n19), .IN2(n25), .IN3(n24), .Q(n23) );
  AO22X1 U70 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n23), .Q(n20) );
  AOI22X1 U71 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n23), .QN(n27) );
  NOR2X0 U72 ( .IN1(in2[3]), .IN2(n24), .QN(n28) );
  AO21X1 U73 ( .IN1(in2[3]), .IN2(n24), .IN3(n28), .Q(n29) );
  OA22X1 U74 ( .IN1(n25), .IN2(n130), .IN3(n140), .IN4(n29), .Q(n26) );
  INVX0 U75 ( .INP(in2[4]), .ZN(n33) );
  OA21X1 U76 ( .IN1(n28), .IN2(n33), .IN3(n32), .Q(n34) );
  AOI22X1 U77 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n34), .QN(n31) );
  OA22X1 U78 ( .IN1(n66), .IN2(n33), .IN3(n141), .IN4(n29), .Q(n30) );
  NOR2X0 U79 ( .IN1(in2[5]), .IN2(n32), .QN(n37) );
  AO21X1 U80 ( .IN1(in2[5]), .IN2(n32), .IN3(n37), .Q(n38) );
  OA22X1 U81 ( .IN1(n33), .IN2(n130), .IN3(n140), .IN4(n38), .Q(n36) );
  AOI22X1 U82 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n34), .QN(n35) );
  INVX0 U83 ( .INP(in2[6]), .ZN(n42) );
  OA21X1 U84 ( .IN1(n37), .IN2(n42), .IN3(n41), .Q(n43) );
  AOI22X1 U85 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n43), .QN(n40) );
  OA22X1 U86 ( .IN1(n66), .IN2(n42), .IN3(n141), .IN4(n38), .Q(n39) );
  NOR2X0 U87 ( .IN1(in2[7]), .IN2(n41), .QN(n46) );
  AO21X1 U88 ( .IN1(in2[7]), .IN2(n41), .IN3(n46), .Q(n47) );
  OA22X1 U89 ( .IN1(n42), .IN2(n130), .IN3(n140), .IN4(n47), .Q(n45) );
  AOI22X1 U90 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n43), .QN(n44) );
  INVX0 U91 ( .INP(in2[8]), .ZN(n51) );
  OA21X1 U92 ( .IN1(n46), .IN2(n51), .IN3(n50), .Q(n52) );
  AOI22X1 U93 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n52), .QN(n49) );
  OA22X1 U94 ( .IN1(n66), .IN2(n51), .IN3(n141), .IN4(n47), .Q(n48) );
  NOR2X0 U95 ( .IN1(in2[9]), .IN2(n50), .QN(n55) );
  AO21X1 U96 ( .IN1(in2[9]), .IN2(n50), .IN3(n55), .Q(n56) );
  OA22X1 U97 ( .IN1(n51), .IN2(n130), .IN3(n140), .IN4(n56), .Q(n54) );
  AOI22X1 U98 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n52), .QN(n53) );
  INVX0 U99 ( .INP(in2[10]), .ZN(n60) );
  OA21X1 U100 ( .IN1(n55), .IN2(n60), .IN3(n59), .Q(n61) );
  AOI22X1 U101 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n61), .QN(n58) );
  OA22X1 U102 ( .IN1(n66), .IN2(n60), .IN3(n141), .IN4(n56), .Q(n57) );
  NOR2X0 U103 ( .IN1(in2[11]), .IN2(n59), .QN(n64) );
  AO21X1 U104 ( .IN1(in2[11]), .IN2(n59), .IN3(n64), .Q(n65) );
  OA22X1 U105 ( .IN1(n60), .IN2(n130), .IN3(n140), .IN4(n65), .Q(n63) );
  AOI22X1 U106 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n61), .QN(n62) );
  INVX0 U107 ( .INP(in2[12]), .ZN(n71) );
  OA21X1 U108 ( .IN1(n64), .IN2(n71), .IN3(n77), .Q(n69) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n69), .QN(n68) );
  OA22X1 U110 ( .IN1(n66), .IN2(n71), .IN3(n141), .IN4(n65), .Q(n67) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n6), .S(n70), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n71), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n7), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n6), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n6), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n8), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n7), .IN4(n85), .IN5(n84), .Q(
        out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n9), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n8), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n8), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n10), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n9), .IN4(n97), .IN5(n96), .Q(
        out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n11), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n10), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n10), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n12), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n11), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n13), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n12), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n12), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n14), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n13), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n15), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n14), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n14), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n15), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_84 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n46), .IN2(n51), .QN(n50) );
  NAND2X0 U4 ( .IN1(n55), .IN2(n60), .QN(n59) );
  NAND2X0 U5 ( .IN1(n19), .IN2(n25), .QN(n24) );
  NAND2X0 U6 ( .IN1(n28), .IN2(n33), .QN(n32) );
  NAND2X0 U7 ( .IN1(n37), .IN2(n42), .QN(n41) );
  NAND2X0 U8 ( .IN1(n64), .IN2(n71), .QN(n77) );
  NAND2X0 U9 ( .IN1(n81), .IN2(n7), .QN(n89) );
  NAND2X0 U10 ( .IN1(n93), .IN2(n9), .QN(n101) );
  NAND2X0 U11 ( .IN1(n105), .IN2(n11), .QN(n114) );
  NAND2X0 U12 ( .IN1(in1[2]), .IN2(n77), .QN(n70) );
  NAND2X0 U13 ( .IN1(n69), .IN2(n132), .QN(n74) );
  NAND2X0 U14 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U15 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U16 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U17 ( .IN1(n118), .IN2(n13), .QN(n125) );
  NAND2X0 U18 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U19 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U20 ( .IN1(n21), .IN2(n132), .QN(n4) );
  NAND2X0 U21 ( .IN1(n45), .IN2(n44), .QN(out1[7]) );
  NAND2X0 U22 ( .IN1(n49), .IN2(n48), .QN(out1[8]) );
  NAND2X0 U23 ( .IN1(n54), .IN2(n53), .QN(out1[9]) );
  NAND2X0 U24 ( .IN1(n58), .IN2(n57), .QN(out1[10]) );
  NAND2X0 U25 ( .IN1(n63), .IN2(n62), .QN(out1[11]) );
  NAND2X0 U26 ( .IN1(n68), .IN2(n67), .QN(out1[12]) );
  NAND2X0 U27 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U28 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U29 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U30 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U31 ( .IN1(n141), .IN2(n130), .QN(n18) );
  NAND2X0 U32 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NAND2X0 U33 ( .IN1(n31), .IN2(n30), .QN(out1[4]) );
  NAND2X0 U34 ( .IN1(n27), .IN2(n26), .QN(out1[3]) );
  NAND2X0 U35 ( .IN1(n36), .IN2(n35), .QN(out1[5]) );
  NAND2X0 U36 ( .IN1(n40), .IN2(n39), .QN(out1[6]) );
  NAND2X0 U37 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U38 ( .IN1(n17), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U39 ( .IN1(in1[2]), .IN2(n16), .QN(n17) );
  NOR2X0 U40 ( .IN1(n22), .IN2(n20), .QN(n3) );
  INVX0 U41 ( .INP(n130), .ZN(n137) );
  NAND3X0 U42 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  NOR2X0 U43 ( .IN1(n142), .IN2(n15), .QN(n1) );
  NOR2X0 U44 ( .IN1(n142), .IN2(n111), .QN(n138) );
  MUX21X1 U45 ( .IN1(n16), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  INVX0 U46 ( .INP(n132), .ZN(n141) );
  NOR3X0 U47 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  INVX0 U48 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U49 ( .INP(in2[13]), .ZN(n6) );
  INVX0 U50 ( .INP(in2[14]), .ZN(n7) );
  INVX0 U51 ( .INP(in2[15]), .ZN(n8) );
  INVX0 U52 ( .INP(in2[16]), .ZN(n9) );
  INVX0 U53 ( .INP(in2[17]), .ZN(n10) );
  INVX0 U54 ( .INP(in2[18]), .ZN(n11) );
  INVX0 U55 ( .INP(in2[19]), .ZN(n12) );
  INVX0 U56 ( .INP(in2[20]), .ZN(n13) );
  INVX0 U57 ( .INP(in2[21]), .ZN(n14) );
  INVX0 U58 ( .INP(in2[22]), .ZN(n15) );
  INVX0 U59 ( .INP(in1[1]), .ZN(n16) );
  INVX0 U60 ( .INP(in1[2]), .ZN(n111) );
  INVX0 U61 ( .INP(n138), .ZN(n140) );
  NOR2X0 U62 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n19) );
  AOI21X1 U63 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n19), .QN(n21) );
  NOR2X0 U64 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U65 ( .IN1(n18), .IN2(in2[0]), .IN3(n138), .IN4(n21), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U66 ( .INP(n133), .ZN(n66) );
  INVX0 U67 ( .INP(in2[2]), .ZN(n25) );
  NOR2X0 U68 ( .IN1(n66), .IN2(n25), .QN(n22) );
  OA21X1 U69 ( .IN1(n19), .IN2(n25), .IN3(n24), .Q(n23) );
  AO22X1 U70 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n23), .Q(n20) );
  AOI22X1 U71 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n23), .QN(n27) );
  NOR2X0 U72 ( .IN1(in2[3]), .IN2(n24), .QN(n28) );
  AO21X1 U73 ( .IN1(in2[3]), .IN2(n24), .IN3(n28), .Q(n29) );
  OA22X1 U74 ( .IN1(n25), .IN2(n130), .IN3(n140), .IN4(n29), .Q(n26) );
  INVX0 U75 ( .INP(in2[4]), .ZN(n33) );
  OA21X1 U76 ( .IN1(n28), .IN2(n33), .IN3(n32), .Q(n34) );
  AOI22X1 U77 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n34), .QN(n31) );
  OA22X1 U78 ( .IN1(n66), .IN2(n33), .IN3(n141), .IN4(n29), .Q(n30) );
  NOR2X0 U79 ( .IN1(in2[5]), .IN2(n32), .QN(n37) );
  AO21X1 U80 ( .IN1(in2[5]), .IN2(n32), .IN3(n37), .Q(n38) );
  OA22X1 U81 ( .IN1(n33), .IN2(n130), .IN3(n140), .IN4(n38), .Q(n36) );
  AOI22X1 U82 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n34), .QN(n35) );
  INVX0 U83 ( .INP(in2[6]), .ZN(n42) );
  OA21X1 U84 ( .IN1(n37), .IN2(n42), .IN3(n41), .Q(n43) );
  AOI22X1 U85 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n43), .QN(n40) );
  OA22X1 U86 ( .IN1(n66), .IN2(n42), .IN3(n141), .IN4(n38), .Q(n39) );
  NOR2X0 U87 ( .IN1(in2[7]), .IN2(n41), .QN(n46) );
  AO21X1 U88 ( .IN1(in2[7]), .IN2(n41), .IN3(n46), .Q(n47) );
  OA22X1 U89 ( .IN1(n42), .IN2(n130), .IN3(n140), .IN4(n47), .Q(n45) );
  AOI22X1 U90 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n43), .QN(n44) );
  INVX0 U91 ( .INP(in2[8]), .ZN(n51) );
  OA21X1 U92 ( .IN1(n46), .IN2(n51), .IN3(n50), .Q(n52) );
  AOI22X1 U93 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n52), .QN(n49) );
  OA22X1 U94 ( .IN1(n66), .IN2(n51), .IN3(n141), .IN4(n47), .Q(n48) );
  NOR2X0 U95 ( .IN1(in2[9]), .IN2(n50), .QN(n55) );
  AO21X1 U96 ( .IN1(in2[9]), .IN2(n50), .IN3(n55), .Q(n56) );
  OA22X1 U97 ( .IN1(n51), .IN2(n130), .IN3(n140), .IN4(n56), .Q(n54) );
  AOI22X1 U98 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n52), .QN(n53) );
  INVX0 U99 ( .INP(in2[10]), .ZN(n60) );
  OA21X1 U100 ( .IN1(n55), .IN2(n60), .IN3(n59), .Q(n61) );
  AOI22X1 U101 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n61), .QN(n58) );
  OA22X1 U102 ( .IN1(n66), .IN2(n60), .IN3(n141), .IN4(n56), .Q(n57) );
  NOR2X0 U103 ( .IN1(in2[11]), .IN2(n59), .QN(n64) );
  AO21X1 U104 ( .IN1(in2[11]), .IN2(n59), .IN3(n64), .Q(n65) );
  OA22X1 U105 ( .IN1(n60), .IN2(n130), .IN3(n140), .IN4(n65), .Q(n63) );
  AOI22X1 U106 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n61), .QN(n62) );
  INVX0 U107 ( .INP(in2[12]), .ZN(n71) );
  OA21X1 U108 ( .IN1(n64), .IN2(n71), .IN3(n77), .Q(n69) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n69), .QN(n68) );
  OA22X1 U110 ( .IN1(n66), .IN2(n71), .IN3(n141), .IN4(n65), .Q(n67) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n6), .S(n70), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n71), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n7), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n6), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n6), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n8), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n7), .IN4(n85), .IN5(n84), .Q(
        out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n9), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n8), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n8), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n10), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n9), .IN4(n97), .IN5(n96), .Q(
        out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n11), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n10), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n10), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n12), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n11), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n13), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n12), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n12), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n14), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n13), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n15), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n14), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n14), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n15), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_85 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n55), .IN2(n60), .QN(n59) );
  NAND2X0 U4 ( .IN1(n28), .IN2(n33), .QN(n32) );
  NAND2X0 U5 ( .IN1(n46), .IN2(n51), .QN(n50) );
  NAND2X0 U6 ( .IN1(n37), .IN2(n42), .QN(n41) );
  NAND2X0 U7 ( .IN1(n64), .IN2(n71), .QN(n77) );
  NAND2X0 U8 ( .IN1(n81), .IN2(n7), .QN(n89) );
  NAND2X0 U9 ( .IN1(n93), .IN2(n9), .QN(n101) );
  NAND2X0 U10 ( .IN1(n105), .IN2(n11), .QN(n114) );
  NAND2X0 U11 ( .IN1(n118), .IN2(n13), .QN(n125) );
  NAND2X0 U12 ( .IN1(n19), .IN2(n25), .QN(n24) );
  NAND2X0 U13 ( .IN1(in1[2]), .IN2(n77), .QN(n70) );
  NAND2X0 U14 ( .IN1(n69), .IN2(n132), .QN(n74) );
  NAND2X0 U15 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U16 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U17 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U18 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U19 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U20 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U21 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U22 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U23 ( .IN1(n54), .IN2(n53), .QN(out1[9]) );
  NAND2X0 U24 ( .IN1(n58), .IN2(n57), .QN(out1[10]) );
  NAND2X0 U25 ( .IN1(n63), .IN2(n62), .QN(out1[11]) );
  NAND2X0 U26 ( .IN1(n68), .IN2(n67), .QN(out1[12]) );
  NAND2X0 U27 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U28 ( .IN1(n17), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U29 ( .IN1(in1[2]), .IN2(n16), .QN(n17) );
  NAND2X0 U30 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NAND2X0 U31 ( .IN1(n21), .IN2(n132), .QN(n4) );
  NAND2X0 U32 ( .IN1(n27), .IN2(n26), .QN(out1[3]) );
  NAND2X0 U33 ( .IN1(n31), .IN2(n30), .QN(out1[4]) );
  NAND2X0 U34 ( .IN1(n40), .IN2(n39), .QN(out1[6]) );
  NAND2X0 U35 ( .IN1(n36), .IN2(n35), .QN(out1[5]) );
  NAND2X0 U36 ( .IN1(n45), .IN2(n44), .QN(out1[7]) );
  NAND2X0 U37 ( .IN1(n49), .IN2(n48), .QN(out1[8]) );
  NAND2X0 U38 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U39 ( .IN1(n141), .IN2(n130), .QN(n18) );
  NOR2X0 U40 ( .IN1(n22), .IN2(n20), .QN(n3) );
  NOR2X0 U41 ( .IN1(n142), .IN2(n15), .QN(n1) );
  INVX0 U42 ( .INP(n132), .ZN(n141) );
  INVX0 U43 ( .INP(n130), .ZN(n137) );
  NAND3X0 U44 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  NOR3X0 U45 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  NOR2X0 U46 ( .IN1(n142), .IN2(n111), .QN(n138) );
  MUX21X1 U47 ( .IN1(n16), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  INVX0 U48 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U49 ( .INP(in2[13]), .ZN(n6) );
  INVX0 U50 ( .INP(in2[14]), .ZN(n7) );
  INVX0 U51 ( .INP(in2[15]), .ZN(n8) );
  INVX0 U52 ( .INP(in2[16]), .ZN(n9) );
  INVX0 U53 ( .INP(in2[17]), .ZN(n10) );
  INVX0 U54 ( .INP(in2[18]), .ZN(n11) );
  INVX0 U55 ( .INP(in2[19]), .ZN(n12) );
  INVX0 U56 ( .INP(in2[20]), .ZN(n13) );
  INVX0 U57 ( .INP(in2[21]), .ZN(n14) );
  INVX0 U58 ( .INP(in2[22]), .ZN(n15) );
  INVX0 U59 ( .INP(in1[1]), .ZN(n16) );
  INVX0 U60 ( .INP(in1[2]), .ZN(n111) );
  INVX0 U61 ( .INP(n138), .ZN(n140) );
  NOR2X0 U62 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n19) );
  AOI21X1 U63 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n19), .QN(n21) );
  NOR2X0 U64 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U65 ( .IN1(n18), .IN2(in2[0]), .IN3(n138), .IN4(n21), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U66 ( .INP(n133), .ZN(n66) );
  INVX0 U67 ( .INP(in2[2]), .ZN(n25) );
  NOR2X0 U68 ( .IN1(n66), .IN2(n25), .QN(n22) );
  OA21X1 U69 ( .IN1(n19), .IN2(n25), .IN3(n24), .Q(n23) );
  AO22X1 U70 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n23), .Q(n20) );
  AOI22X1 U71 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n23), .QN(n27) );
  NOR2X0 U72 ( .IN1(in2[3]), .IN2(n24), .QN(n28) );
  AO21X1 U73 ( .IN1(in2[3]), .IN2(n24), .IN3(n28), .Q(n29) );
  OA22X1 U74 ( .IN1(n25), .IN2(n130), .IN3(n140), .IN4(n29), .Q(n26) );
  INVX0 U75 ( .INP(in2[4]), .ZN(n33) );
  OA21X1 U76 ( .IN1(n28), .IN2(n33), .IN3(n32), .Q(n34) );
  AOI22X1 U77 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n34), .QN(n31) );
  OA22X1 U78 ( .IN1(n66), .IN2(n33), .IN3(n141), .IN4(n29), .Q(n30) );
  NOR2X0 U79 ( .IN1(in2[5]), .IN2(n32), .QN(n37) );
  AO21X1 U80 ( .IN1(in2[5]), .IN2(n32), .IN3(n37), .Q(n38) );
  OA22X1 U81 ( .IN1(n33), .IN2(n130), .IN3(n140), .IN4(n38), .Q(n36) );
  AOI22X1 U82 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n34), .QN(n35) );
  INVX0 U83 ( .INP(in2[6]), .ZN(n42) );
  OA21X1 U84 ( .IN1(n37), .IN2(n42), .IN3(n41), .Q(n43) );
  AOI22X1 U85 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n43), .QN(n40) );
  OA22X1 U86 ( .IN1(n66), .IN2(n42), .IN3(n141), .IN4(n38), .Q(n39) );
  NOR2X0 U87 ( .IN1(in2[7]), .IN2(n41), .QN(n46) );
  AO21X1 U88 ( .IN1(in2[7]), .IN2(n41), .IN3(n46), .Q(n47) );
  OA22X1 U89 ( .IN1(n42), .IN2(n130), .IN3(n140), .IN4(n47), .Q(n45) );
  AOI22X1 U90 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n43), .QN(n44) );
  INVX0 U91 ( .INP(in2[8]), .ZN(n51) );
  OA21X1 U92 ( .IN1(n46), .IN2(n51), .IN3(n50), .Q(n52) );
  AOI22X1 U93 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n52), .QN(n49) );
  OA22X1 U94 ( .IN1(n66), .IN2(n51), .IN3(n141), .IN4(n47), .Q(n48) );
  NOR2X0 U95 ( .IN1(in2[9]), .IN2(n50), .QN(n55) );
  AO21X1 U96 ( .IN1(in2[9]), .IN2(n50), .IN3(n55), .Q(n56) );
  OA22X1 U97 ( .IN1(n51), .IN2(n130), .IN3(n140), .IN4(n56), .Q(n54) );
  AOI22X1 U98 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n52), .QN(n53) );
  INVX0 U99 ( .INP(in2[10]), .ZN(n60) );
  OA21X1 U100 ( .IN1(n55), .IN2(n60), .IN3(n59), .Q(n61) );
  AOI22X1 U101 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n61), .QN(n58) );
  OA22X1 U102 ( .IN1(n66), .IN2(n60), .IN3(n141), .IN4(n56), .Q(n57) );
  NOR2X0 U103 ( .IN1(in2[11]), .IN2(n59), .QN(n64) );
  AO21X1 U104 ( .IN1(in2[11]), .IN2(n59), .IN3(n64), .Q(n65) );
  OA22X1 U105 ( .IN1(n60), .IN2(n130), .IN3(n140), .IN4(n65), .Q(n63) );
  AOI22X1 U106 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n61), .QN(n62) );
  INVX0 U107 ( .INP(in2[12]), .ZN(n71) );
  OA21X1 U108 ( .IN1(n64), .IN2(n71), .IN3(n77), .Q(n69) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n69), .QN(n68) );
  OA22X1 U110 ( .IN1(n66), .IN2(n71), .IN3(n141), .IN4(n65), .Q(n67) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n6), .S(n70), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n71), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n7), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n6), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n6), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n8), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n7), .IN4(n85), .IN5(n84), .Q(
        out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n9), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n8), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n8), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n10), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n9), .IN4(n97), .IN5(n96), .Q(
        out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n11), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n10), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n10), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n12), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n11), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n13), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n12), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n12), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n14), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n13), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n15), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n14), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n14), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n15), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_86 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n55), .IN2(n60), .QN(n59) );
  NAND2X0 U4 ( .IN1(n19), .IN2(n25), .QN(n24) );
  NAND2X0 U5 ( .IN1(n28), .IN2(n33), .QN(n32) );
  NAND2X0 U6 ( .IN1(n46), .IN2(n51), .QN(n50) );
  NAND2X0 U7 ( .IN1(n37), .IN2(n42), .QN(n41) );
  NAND2X0 U8 ( .IN1(n64), .IN2(n71), .QN(n77) );
  NAND2X0 U9 ( .IN1(n81), .IN2(n7), .QN(n89) );
  NAND2X0 U10 ( .IN1(n93), .IN2(n9), .QN(n101) );
  NAND2X0 U11 ( .IN1(n105), .IN2(n11), .QN(n114) );
  NAND2X0 U12 ( .IN1(in1[2]), .IN2(n77), .QN(n70) );
  NAND2X0 U13 ( .IN1(n69), .IN2(n132), .QN(n74) );
  NAND2X0 U14 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U15 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U16 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U17 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U18 ( .IN1(n118), .IN2(n13), .QN(n125) );
  NAND2X0 U19 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U20 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U21 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U22 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U23 ( .IN1(n141), .IN2(n130), .QN(n18) );
  NAND2X0 U24 ( .IN1(n21), .IN2(n132), .QN(n4) );
  NAND2X0 U25 ( .IN1(n54), .IN2(n53), .QN(out1[9]) );
  NAND2X0 U26 ( .IN1(n58), .IN2(n57), .QN(out1[10]) );
  NAND2X0 U27 ( .IN1(n63), .IN2(n62), .QN(out1[11]) );
  NAND2X0 U28 ( .IN1(n68), .IN2(n67), .QN(out1[12]) );
  NAND2X0 U29 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U30 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U31 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NAND2X0 U32 ( .IN1(n27), .IN2(n26), .QN(out1[3]) );
  NAND2X0 U33 ( .IN1(n31), .IN2(n30), .QN(out1[4]) );
  NAND2X0 U34 ( .IN1(n36), .IN2(n35), .QN(out1[5]) );
  NAND2X0 U35 ( .IN1(n40), .IN2(n39), .QN(out1[6]) );
  NAND2X0 U36 ( .IN1(n45), .IN2(n44), .QN(out1[7]) );
  NAND2X0 U37 ( .IN1(n49), .IN2(n48), .QN(out1[8]) );
  NAND2X0 U38 ( .IN1(n17), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U39 ( .IN1(in1[2]), .IN2(n16), .QN(n17) );
  NOR2X0 U40 ( .IN1(n22), .IN2(n20), .QN(n3) );
  NOR2X0 U41 ( .IN1(n142), .IN2(n15), .QN(n1) );
  INVX0 U42 ( .INP(n132), .ZN(n141) );
  INVX0 U43 ( .INP(n130), .ZN(n137) );
  NAND3X0 U44 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  NOR3X0 U45 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  NOR2X0 U46 ( .IN1(n142), .IN2(n111), .QN(n138) );
  MUX21X1 U47 ( .IN1(n16), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  INVX0 U48 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U49 ( .INP(in2[13]), .ZN(n6) );
  INVX0 U50 ( .INP(in2[14]), .ZN(n7) );
  INVX0 U51 ( .INP(in2[15]), .ZN(n8) );
  INVX0 U52 ( .INP(in2[16]), .ZN(n9) );
  INVX0 U53 ( .INP(in2[17]), .ZN(n10) );
  INVX0 U54 ( .INP(in2[18]), .ZN(n11) );
  INVX0 U55 ( .INP(in2[19]), .ZN(n12) );
  INVX0 U56 ( .INP(in2[20]), .ZN(n13) );
  INVX0 U57 ( .INP(in2[21]), .ZN(n14) );
  INVX0 U58 ( .INP(in2[22]), .ZN(n15) );
  INVX0 U59 ( .INP(in1[1]), .ZN(n16) );
  INVX0 U60 ( .INP(in1[2]), .ZN(n111) );
  INVX0 U61 ( .INP(n138), .ZN(n140) );
  NOR2X0 U62 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n19) );
  AOI21X1 U63 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n19), .QN(n21) );
  NOR2X0 U64 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U65 ( .IN1(n18), .IN2(in2[0]), .IN3(n138), .IN4(n21), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U66 ( .INP(n133), .ZN(n66) );
  INVX0 U67 ( .INP(in2[2]), .ZN(n25) );
  NOR2X0 U68 ( .IN1(n66), .IN2(n25), .QN(n22) );
  OA21X1 U69 ( .IN1(n19), .IN2(n25), .IN3(n24), .Q(n23) );
  AO22X1 U70 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n23), .Q(n20) );
  AOI22X1 U71 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n23), .QN(n27) );
  NOR2X0 U72 ( .IN1(in2[3]), .IN2(n24), .QN(n28) );
  AO21X1 U73 ( .IN1(in2[3]), .IN2(n24), .IN3(n28), .Q(n29) );
  OA22X1 U74 ( .IN1(n25), .IN2(n130), .IN3(n140), .IN4(n29), .Q(n26) );
  INVX0 U75 ( .INP(in2[4]), .ZN(n33) );
  OA21X1 U76 ( .IN1(n28), .IN2(n33), .IN3(n32), .Q(n34) );
  AOI22X1 U77 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n34), .QN(n31) );
  OA22X1 U78 ( .IN1(n66), .IN2(n33), .IN3(n141), .IN4(n29), .Q(n30) );
  NOR2X0 U79 ( .IN1(in2[5]), .IN2(n32), .QN(n37) );
  AO21X1 U80 ( .IN1(in2[5]), .IN2(n32), .IN3(n37), .Q(n38) );
  OA22X1 U81 ( .IN1(n33), .IN2(n130), .IN3(n140), .IN4(n38), .Q(n36) );
  AOI22X1 U82 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n34), .QN(n35) );
  INVX0 U83 ( .INP(in2[6]), .ZN(n42) );
  OA21X1 U84 ( .IN1(n37), .IN2(n42), .IN3(n41), .Q(n43) );
  AOI22X1 U85 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n43), .QN(n40) );
  OA22X1 U86 ( .IN1(n66), .IN2(n42), .IN3(n141), .IN4(n38), .Q(n39) );
  NOR2X0 U87 ( .IN1(in2[7]), .IN2(n41), .QN(n46) );
  AO21X1 U88 ( .IN1(in2[7]), .IN2(n41), .IN3(n46), .Q(n47) );
  OA22X1 U89 ( .IN1(n42), .IN2(n130), .IN3(n140), .IN4(n47), .Q(n45) );
  AOI22X1 U90 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n43), .QN(n44) );
  INVX0 U91 ( .INP(in2[8]), .ZN(n51) );
  OA21X1 U92 ( .IN1(n46), .IN2(n51), .IN3(n50), .Q(n52) );
  AOI22X1 U93 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n52), .QN(n49) );
  OA22X1 U94 ( .IN1(n66), .IN2(n51), .IN3(n141), .IN4(n47), .Q(n48) );
  NOR2X0 U95 ( .IN1(in2[9]), .IN2(n50), .QN(n55) );
  AO21X1 U96 ( .IN1(in2[9]), .IN2(n50), .IN3(n55), .Q(n56) );
  OA22X1 U97 ( .IN1(n51), .IN2(n130), .IN3(n140), .IN4(n56), .Q(n54) );
  AOI22X1 U98 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n52), .QN(n53) );
  INVX0 U99 ( .INP(in2[10]), .ZN(n60) );
  OA21X1 U100 ( .IN1(n55), .IN2(n60), .IN3(n59), .Q(n61) );
  AOI22X1 U101 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n61), .QN(n58) );
  OA22X1 U102 ( .IN1(n66), .IN2(n60), .IN3(n141), .IN4(n56), .Q(n57) );
  NOR2X0 U103 ( .IN1(in2[11]), .IN2(n59), .QN(n64) );
  AO21X1 U104 ( .IN1(in2[11]), .IN2(n59), .IN3(n64), .Q(n65) );
  OA22X1 U105 ( .IN1(n60), .IN2(n130), .IN3(n140), .IN4(n65), .Q(n63) );
  AOI22X1 U106 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n61), .QN(n62) );
  INVX0 U107 ( .INP(in2[12]), .ZN(n71) );
  OA21X1 U108 ( .IN1(n64), .IN2(n71), .IN3(n77), .Q(n69) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n69), .QN(n68) );
  OA22X1 U110 ( .IN1(n66), .IN2(n71), .IN3(n141), .IN4(n65), .Q(n67) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n6), .S(n70), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n71), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n7), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n6), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n6), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n8), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n7), .IN4(n85), .IN5(n84), .Q(
        out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n9), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n8), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n8), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n10), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n9), .IN4(n97), .IN5(n96), .Q(
        out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n11), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n10), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n10), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n12), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n11), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n13), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n12), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n12), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n14), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n13), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n15), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n14), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n14), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n15), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_87 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n19), .IN2(n25), .QN(n24) );
  NAND2X0 U4 ( .IN1(n28), .IN2(n33), .QN(n32) );
  NAND2X0 U5 ( .IN1(n37), .IN2(n42), .QN(n41) );
  NAND2X0 U6 ( .IN1(n55), .IN2(n60), .QN(n59) );
  NAND2X0 U7 ( .IN1(n46), .IN2(n51), .QN(n50) );
  NAND2X0 U8 ( .IN1(n64), .IN2(n71), .QN(n77) );
  NAND2X0 U9 ( .IN1(n81), .IN2(n7), .QN(n89) );
  NAND2X0 U10 ( .IN1(n93), .IN2(n9), .QN(n101) );
  NAND2X0 U11 ( .IN1(n105), .IN2(n11), .QN(n114) );
  NAND2X0 U12 ( .IN1(n118), .IN2(n13), .QN(n125) );
  NAND2X0 U13 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U14 ( .IN1(in1[2]), .IN2(n77), .QN(n70) );
  NAND2X0 U15 ( .IN1(n69), .IN2(n132), .QN(n74) );
  NAND2X0 U16 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U17 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U18 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U19 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U20 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U21 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U22 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U23 ( .IN1(n141), .IN2(n130), .QN(n18) );
  NAND2X0 U24 ( .IN1(n21), .IN2(n132), .QN(n4) );
  NAND2X0 U25 ( .IN1(n63), .IN2(n62), .QN(out1[11]) );
  NAND2X0 U26 ( .IN1(n68), .IN2(n67), .QN(out1[12]) );
  NAND2X0 U27 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U28 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U29 ( .IN1(n17), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U30 ( .IN1(in1[2]), .IN2(n16), .QN(n17) );
  NAND2X0 U31 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NAND2X0 U32 ( .IN1(n27), .IN2(n26), .QN(out1[3]) );
  NAND2X0 U33 ( .IN1(n31), .IN2(n30), .QN(out1[4]) );
  NAND2X0 U34 ( .IN1(n36), .IN2(n35), .QN(out1[5]) );
  NAND2X0 U35 ( .IN1(n40), .IN2(n39), .QN(out1[6]) );
  NAND2X0 U36 ( .IN1(n45), .IN2(n44), .QN(out1[7]) );
  NAND2X0 U37 ( .IN1(n49), .IN2(n48), .QN(out1[8]) );
  NAND2X0 U38 ( .IN1(n54), .IN2(n53), .QN(out1[9]) );
  NAND2X0 U39 ( .IN1(n58), .IN2(n57), .QN(out1[10]) );
  NOR2X0 U40 ( .IN1(n22), .IN2(n20), .QN(n3) );
  INVX0 U41 ( .INP(n130), .ZN(n137) );
  NAND3X0 U42 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  NOR2X0 U43 ( .IN1(n142), .IN2(n15), .QN(n1) );
  NOR2X0 U44 ( .IN1(n142), .IN2(n111), .QN(n138) );
  MUX21X1 U45 ( .IN1(n16), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  INVX0 U46 ( .INP(n132), .ZN(n141) );
  NOR3X0 U47 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  INVX0 U48 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U49 ( .INP(in2[13]), .ZN(n6) );
  INVX0 U50 ( .INP(in2[14]), .ZN(n7) );
  INVX0 U51 ( .INP(in2[15]), .ZN(n8) );
  INVX0 U52 ( .INP(in2[16]), .ZN(n9) );
  INVX0 U53 ( .INP(in2[17]), .ZN(n10) );
  INVX0 U54 ( .INP(in2[18]), .ZN(n11) );
  INVX0 U55 ( .INP(in2[19]), .ZN(n12) );
  INVX0 U56 ( .INP(in2[20]), .ZN(n13) );
  INVX0 U57 ( .INP(in2[21]), .ZN(n14) );
  INVX0 U58 ( .INP(in2[22]), .ZN(n15) );
  INVX0 U59 ( .INP(in1[1]), .ZN(n16) );
  INVX0 U60 ( .INP(in1[2]), .ZN(n111) );
  INVX0 U61 ( .INP(n138), .ZN(n140) );
  NOR2X0 U62 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n19) );
  AOI21X1 U63 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n19), .QN(n21) );
  NOR2X0 U64 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U65 ( .IN1(n18), .IN2(in2[0]), .IN3(n138), .IN4(n21), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U66 ( .INP(n133), .ZN(n66) );
  INVX0 U67 ( .INP(in2[2]), .ZN(n25) );
  NOR2X0 U68 ( .IN1(n66), .IN2(n25), .QN(n22) );
  OA21X1 U69 ( .IN1(n19), .IN2(n25), .IN3(n24), .Q(n23) );
  AO22X1 U70 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n23), .Q(n20) );
  AOI22X1 U71 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n23), .QN(n27) );
  NOR2X0 U72 ( .IN1(in2[3]), .IN2(n24), .QN(n28) );
  AO21X1 U73 ( .IN1(in2[3]), .IN2(n24), .IN3(n28), .Q(n29) );
  OA22X1 U74 ( .IN1(n25), .IN2(n130), .IN3(n140), .IN4(n29), .Q(n26) );
  INVX0 U75 ( .INP(in2[4]), .ZN(n33) );
  OA21X1 U76 ( .IN1(n28), .IN2(n33), .IN3(n32), .Q(n34) );
  AOI22X1 U77 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n34), .QN(n31) );
  OA22X1 U78 ( .IN1(n66), .IN2(n33), .IN3(n141), .IN4(n29), .Q(n30) );
  NOR2X0 U79 ( .IN1(in2[5]), .IN2(n32), .QN(n37) );
  AO21X1 U80 ( .IN1(in2[5]), .IN2(n32), .IN3(n37), .Q(n38) );
  OA22X1 U81 ( .IN1(n33), .IN2(n130), .IN3(n140), .IN4(n38), .Q(n36) );
  AOI22X1 U82 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n34), .QN(n35) );
  INVX0 U83 ( .INP(in2[6]), .ZN(n42) );
  OA21X1 U84 ( .IN1(n37), .IN2(n42), .IN3(n41), .Q(n43) );
  AOI22X1 U85 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n43), .QN(n40) );
  OA22X1 U86 ( .IN1(n66), .IN2(n42), .IN3(n141), .IN4(n38), .Q(n39) );
  NOR2X0 U87 ( .IN1(in2[7]), .IN2(n41), .QN(n46) );
  AO21X1 U88 ( .IN1(in2[7]), .IN2(n41), .IN3(n46), .Q(n47) );
  OA22X1 U89 ( .IN1(n42), .IN2(n130), .IN3(n140), .IN4(n47), .Q(n45) );
  AOI22X1 U90 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n43), .QN(n44) );
  INVX0 U91 ( .INP(in2[8]), .ZN(n51) );
  OA21X1 U92 ( .IN1(n46), .IN2(n51), .IN3(n50), .Q(n52) );
  AOI22X1 U93 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n52), .QN(n49) );
  OA22X1 U94 ( .IN1(n66), .IN2(n51), .IN3(n141), .IN4(n47), .Q(n48) );
  NOR2X0 U95 ( .IN1(in2[9]), .IN2(n50), .QN(n55) );
  AO21X1 U96 ( .IN1(in2[9]), .IN2(n50), .IN3(n55), .Q(n56) );
  OA22X1 U97 ( .IN1(n51), .IN2(n130), .IN3(n140), .IN4(n56), .Q(n54) );
  AOI22X1 U98 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n52), .QN(n53) );
  INVX0 U99 ( .INP(in2[10]), .ZN(n60) );
  OA21X1 U100 ( .IN1(n55), .IN2(n60), .IN3(n59), .Q(n61) );
  AOI22X1 U101 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n61), .QN(n58) );
  OA22X1 U102 ( .IN1(n66), .IN2(n60), .IN3(n141), .IN4(n56), .Q(n57) );
  NOR2X0 U103 ( .IN1(in2[11]), .IN2(n59), .QN(n64) );
  AO21X1 U104 ( .IN1(in2[11]), .IN2(n59), .IN3(n64), .Q(n65) );
  OA22X1 U105 ( .IN1(n60), .IN2(n130), .IN3(n140), .IN4(n65), .Q(n63) );
  AOI22X1 U106 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n61), .QN(n62) );
  INVX0 U107 ( .INP(in2[12]), .ZN(n71) );
  OA21X1 U108 ( .IN1(n64), .IN2(n71), .IN3(n77), .Q(n69) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n69), .QN(n68) );
  OA22X1 U110 ( .IN1(n66), .IN2(n71), .IN3(n141), .IN4(n65), .Q(n67) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n6), .S(n70), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n71), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n7), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n6), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n6), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n8), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n7), .IN4(n85), .IN5(n84), .Q(
        out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n9), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n8), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n8), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n10), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n9), .IN4(n97), .IN5(n96), .Q(
        out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n11), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n10), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n10), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n12), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n11), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n13), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n12), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n12), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n14), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n13), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n15), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n14), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n14), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n15), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_88 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n19), .IN2(n25), .QN(n24) );
  NAND2X0 U4 ( .IN1(n28), .IN2(n33), .QN(n32) );
  NAND2X0 U5 ( .IN1(n37), .IN2(n42), .QN(n41) );
  NAND2X0 U6 ( .IN1(n46), .IN2(n51), .QN(n50) );
  NAND2X0 U7 ( .IN1(n55), .IN2(n60), .QN(n59) );
  NAND2X0 U8 ( .IN1(n64), .IN2(n71), .QN(n77) );
  NAND2X0 U9 ( .IN1(n81), .IN2(n7), .QN(n89) );
  NAND2X0 U10 ( .IN1(n93), .IN2(n9), .QN(n101) );
  NAND2X0 U11 ( .IN1(n105), .IN2(n11), .QN(n114) );
  NAND2X0 U12 ( .IN1(n118), .IN2(n13), .QN(n125) );
  NAND2X0 U13 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U14 ( .IN1(in1[2]), .IN2(n77), .QN(n70) );
  NAND2X0 U15 ( .IN1(n69), .IN2(n132), .QN(n74) );
  NAND2X0 U16 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U17 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U18 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U19 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U20 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U21 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U22 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U23 ( .IN1(n17), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U24 ( .IN1(in1[2]), .IN2(n16), .QN(n17) );
  NAND2X0 U25 ( .IN1(n27), .IN2(n26), .QN(out1[3]) );
  NAND2X0 U26 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U27 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U28 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NAND2X0 U29 ( .IN1(n21), .IN2(n132), .QN(n4) );
  NAND2X0 U30 ( .IN1(n31), .IN2(n30), .QN(out1[4]) );
  NAND2X0 U31 ( .IN1(n36), .IN2(n35), .QN(out1[5]) );
  NAND2X0 U32 ( .IN1(n40), .IN2(n39), .QN(out1[6]) );
  NAND2X0 U33 ( .IN1(n45), .IN2(n44), .QN(out1[7]) );
  NAND2X0 U34 ( .IN1(n49), .IN2(n48), .QN(out1[8]) );
  NAND2X0 U35 ( .IN1(n54), .IN2(n53), .QN(out1[9]) );
  NAND2X0 U36 ( .IN1(n58), .IN2(n57), .QN(out1[10]) );
  NAND2X0 U37 ( .IN1(n63), .IN2(n62), .QN(out1[11]) );
  NAND2X0 U38 ( .IN1(n68), .IN2(n67), .QN(out1[12]) );
  NAND2X0 U39 ( .IN1(n141), .IN2(n130), .QN(n18) );
  NOR2X0 U40 ( .IN1(n22), .IN2(n20), .QN(n3) );
  NOR2X0 U41 ( .IN1(n142), .IN2(n15), .QN(n1) );
  INVX0 U42 ( .INP(n132), .ZN(n141) );
  INVX0 U43 ( .INP(n130), .ZN(n137) );
  NAND3X0 U44 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  NOR3X0 U45 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  NOR2X0 U46 ( .IN1(n142), .IN2(n111), .QN(n138) );
  MUX21X1 U47 ( .IN1(n16), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  INVX0 U48 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U49 ( .INP(in2[13]), .ZN(n6) );
  INVX0 U50 ( .INP(in2[14]), .ZN(n7) );
  INVX0 U51 ( .INP(in2[15]), .ZN(n8) );
  INVX0 U52 ( .INP(in2[16]), .ZN(n9) );
  INVX0 U53 ( .INP(in2[17]), .ZN(n10) );
  INVX0 U54 ( .INP(in2[18]), .ZN(n11) );
  INVX0 U55 ( .INP(in2[19]), .ZN(n12) );
  INVX0 U56 ( .INP(in2[20]), .ZN(n13) );
  INVX0 U57 ( .INP(in2[21]), .ZN(n14) );
  INVX0 U58 ( .INP(in2[22]), .ZN(n15) );
  INVX0 U59 ( .INP(in1[1]), .ZN(n16) );
  INVX0 U60 ( .INP(in1[2]), .ZN(n111) );
  INVX0 U61 ( .INP(n138), .ZN(n140) );
  NOR2X0 U62 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n19) );
  AOI21X1 U63 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n19), .QN(n21) );
  NOR2X0 U64 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U65 ( .IN1(n18), .IN2(in2[0]), .IN3(n138), .IN4(n21), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U66 ( .INP(n133), .ZN(n66) );
  INVX0 U67 ( .INP(in2[2]), .ZN(n25) );
  NOR2X0 U68 ( .IN1(n66), .IN2(n25), .QN(n22) );
  OA21X1 U69 ( .IN1(n19), .IN2(n25), .IN3(n24), .Q(n23) );
  AO22X1 U70 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n23), .Q(n20) );
  AOI22X1 U71 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n23), .QN(n27) );
  NOR2X0 U72 ( .IN1(in2[3]), .IN2(n24), .QN(n28) );
  AO21X1 U73 ( .IN1(in2[3]), .IN2(n24), .IN3(n28), .Q(n29) );
  OA22X1 U74 ( .IN1(n25), .IN2(n130), .IN3(n140), .IN4(n29), .Q(n26) );
  INVX0 U75 ( .INP(in2[4]), .ZN(n33) );
  OA21X1 U76 ( .IN1(n28), .IN2(n33), .IN3(n32), .Q(n34) );
  AOI22X1 U77 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n34), .QN(n31) );
  OA22X1 U78 ( .IN1(n66), .IN2(n33), .IN3(n141), .IN4(n29), .Q(n30) );
  NOR2X0 U79 ( .IN1(in2[5]), .IN2(n32), .QN(n37) );
  AO21X1 U80 ( .IN1(in2[5]), .IN2(n32), .IN3(n37), .Q(n38) );
  OA22X1 U81 ( .IN1(n33), .IN2(n130), .IN3(n140), .IN4(n38), .Q(n36) );
  AOI22X1 U82 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n34), .QN(n35) );
  INVX0 U83 ( .INP(in2[6]), .ZN(n42) );
  OA21X1 U84 ( .IN1(n37), .IN2(n42), .IN3(n41), .Q(n43) );
  AOI22X1 U85 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n43), .QN(n40) );
  OA22X1 U86 ( .IN1(n66), .IN2(n42), .IN3(n141), .IN4(n38), .Q(n39) );
  NOR2X0 U87 ( .IN1(in2[7]), .IN2(n41), .QN(n46) );
  AO21X1 U88 ( .IN1(in2[7]), .IN2(n41), .IN3(n46), .Q(n47) );
  OA22X1 U89 ( .IN1(n42), .IN2(n130), .IN3(n140), .IN4(n47), .Q(n45) );
  AOI22X1 U90 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n43), .QN(n44) );
  INVX0 U91 ( .INP(in2[8]), .ZN(n51) );
  OA21X1 U92 ( .IN1(n46), .IN2(n51), .IN3(n50), .Q(n52) );
  AOI22X1 U93 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n52), .QN(n49) );
  OA22X1 U94 ( .IN1(n66), .IN2(n51), .IN3(n141), .IN4(n47), .Q(n48) );
  NOR2X0 U95 ( .IN1(in2[9]), .IN2(n50), .QN(n55) );
  AO21X1 U96 ( .IN1(in2[9]), .IN2(n50), .IN3(n55), .Q(n56) );
  OA22X1 U97 ( .IN1(n51), .IN2(n130), .IN3(n140), .IN4(n56), .Q(n54) );
  AOI22X1 U98 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n52), .QN(n53) );
  INVX0 U99 ( .INP(in2[10]), .ZN(n60) );
  OA21X1 U100 ( .IN1(n55), .IN2(n60), .IN3(n59), .Q(n61) );
  AOI22X1 U101 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n61), .QN(n58) );
  OA22X1 U102 ( .IN1(n66), .IN2(n60), .IN3(n141), .IN4(n56), .Q(n57) );
  NOR2X0 U103 ( .IN1(in2[11]), .IN2(n59), .QN(n64) );
  AO21X1 U104 ( .IN1(in2[11]), .IN2(n59), .IN3(n64), .Q(n65) );
  OA22X1 U105 ( .IN1(n60), .IN2(n130), .IN3(n140), .IN4(n65), .Q(n63) );
  AOI22X1 U106 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n61), .QN(n62) );
  INVX0 U107 ( .INP(in2[12]), .ZN(n71) );
  OA21X1 U108 ( .IN1(n64), .IN2(n71), .IN3(n77), .Q(n69) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n69), .QN(n68) );
  OA22X1 U110 ( .IN1(n66), .IN2(n71), .IN3(n141), .IN4(n65), .Q(n67) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n6), .S(n70), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n71), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n7), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n6), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n6), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n8), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n7), .IN4(n85), .IN5(n84), .Q(
        out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n9), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n8), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n8), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n10), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n9), .IN4(n97), .IN5(n96), .Q(
        out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n11), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n10), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n10), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n12), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n11), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n13), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n12), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n12), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n14), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n13), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n15), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n14), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n14), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n15), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_89 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n19), .IN2(n25), .QN(n24) );
  NAND2X0 U4 ( .IN1(n28), .IN2(n33), .QN(n32) );
  NAND2X0 U5 ( .IN1(n37), .IN2(n42), .QN(n41) );
  NAND2X0 U6 ( .IN1(n46), .IN2(n51), .QN(n50) );
  NAND2X0 U7 ( .IN1(n55), .IN2(n60), .QN(n59) );
  NAND2X0 U8 ( .IN1(n64), .IN2(n71), .QN(n77) );
  NAND2X0 U9 ( .IN1(n81), .IN2(n7), .QN(n89) );
  NAND2X0 U10 ( .IN1(n105), .IN2(n11), .QN(n114) );
  NAND2X0 U11 ( .IN1(n93), .IN2(n9), .QN(n101) );
  NAND2X0 U12 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U13 ( .IN1(n118), .IN2(n13), .QN(n125) );
  NAND2X0 U14 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U15 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U16 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U17 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U18 ( .IN1(n21), .IN2(n132), .QN(n4) );
  NAND2X0 U19 ( .IN1(n141), .IN2(n130), .QN(n18) );
  NAND2X0 U20 ( .IN1(n27), .IN2(n26), .QN(out1[3]) );
  NAND2X0 U21 ( .IN1(n31), .IN2(n30), .QN(out1[4]) );
  NAND2X0 U22 ( .IN1(in1[2]), .IN2(n77), .QN(n70) );
  NAND2X0 U23 ( .IN1(n69), .IN2(n132), .QN(n74) );
  NAND2X0 U24 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U25 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U26 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U27 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U28 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NAND2X0 U29 ( .IN1(n36), .IN2(n35), .QN(out1[5]) );
  NAND2X0 U30 ( .IN1(n40), .IN2(n39), .QN(out1[6]) );
  NAND2X0 U31 ( .IN1(n45), .IN2(n44), .QN(out1[7]) );
  NAND2X0 U32 ( .IN1(n49), .IN2(n48), .QN(out1[8]) );
  NAND2X0 U33 ( .IN1(n54), .IN2(n53), .QN(out1[9]) );
  NAND2X0 U34 ( .IN1(n58), .IN2(n57), .QN(out1[10]) );
  NAND2X0 U35 ( .IN1(n63), .IN2(n62), .QN(out1[11]) );
  NAND2X0 U36 ( .IN1(n68), .IN2(n67), .QN(out1[12]) );
  NAND2X0 U37 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U38 ( .IN1(n17), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U39 ( .IN1(in1[2]), .IN2(n16), .QN(n17) );
  NOR2X0 U40 ( .IN1(n22), .IN2(n20), .QN(n3) );
  INVX0 U41 ( .INP(n130), .ZN(n137) );
  INVX0 U42 ( .INP(n132), .ZN(n141) );
  NOR3X0 U43 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  NAND3X0 U44 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  NOR2X0 U45 ( .IN1(n142), .IN2(n15), .QN(n1) );
  NOR2X0 U46 ( .IN1(n142), .IN2(n111), .QN(n138) );
  MUX21X1 U47 ( .IN1(n16), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  INVX0 U48 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U49 ( .INP(in2[13]), .ZN(n6) );
  INVX0 U50 ( .INP(in2[14]), .ZN(n7) );
  INVX0 U51 ( .INP(in2[15]), .ZN(n8) );
  INVX0 U52 ( .INP(in2[16]), .ZN(n9) );
  INVX0 U53 ( .INP(in2[17]), .ZN(n10) );
  INVX0 U54 ( .INP(in2[18]), .ZN(n11) );
  INVX0 U55 ( .INP(in2[19]), .ZN(n12) );
  INVX0 U56 ( .INP(in2[20]), .ZN(n13) );
  INVX0 U57 ( .INP(in2[21]), .ZN(n14) );
  INVX0 U58 ( .INP(in2[22]), .ZN(n15) );
  INVX0 U59 ( .INP(in1[1]), .ZN(n16) );
  INVX0 U60 ( .INP(in1[2]), .ZN(n111) );
  INVX0 U61 ( .INP(n138), .ZN(n140) );
  NOR2X0 U62 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n19) );
  AOI21X1 U63 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n19), .QN(n21) );
  NOR2X0 U64 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U65 ( .IN1(n18), .IN2(in2[0]), .IN3(n138), .IN4(n21), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U66 ( .INP(n133), .ZN(n66) );
  INVX0 U67 ( .INP(in2[2]), .ZN(n25) );
  NOR2X0 U68 ( .IN1(n66), .IN2(n25), .QN(n22) );
  OA21X1 U69 ( .IN1(n19), .IN2(n25), .IN3(n24), .Q(n23) );
  AO22X1 U70 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n23), .Q(n20) );
  AOI22X1 U71 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n23), .QN(n27) );
  NOR2X0 U72 ( .IN1(in2[3]), .IN2(n24), .QN(n28) );
  AO21X1 U73 ( .IN1(in2[3]), .IN2(n24), .IN3(n28), .Q(n29) );
  OA22X1 U74 ( .IN1(n25), .IN2(n130), .IN3(n140), .IN4(n29), .Q(n26) );
  INVX0 U75 ( .INP(in2[4]), .ZN(n33) );
  OA21X1 U76 ( .IN1(n28), .IN2(n33), .IN3(n32), .Q(n34) );
  AOI22X1 U77 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n34), .QN(n31) );
  OA22X1 U78 ( .IN1(n66), .IN2(n33), .IN3(n141), .IN4(n29), .Q(n30) );
  NOR2X0 U79 ( .IN1(in2[5]), .IN2(n32), .QN(n37) );
  AO21X1 U80 ( .IN1(in2[5]), .IN2(n32), .IN3(n37), .Q(n38) );
  OA22X1 U81 ( .IN1(n33), .IN2(n130), .IN3(n140), .IN4(n38), .Q(n36) );
  AOI22X1 U82 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n34), .QN(n35) );
  INVX0 U83 ( .INP(in2[6]), .ZN(n42) );
  OA21X1 U84 ( .IN1(n37), .IN2(n42), .IN3(n41), .Q(n43) );
  AOI22X1 U85 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n43), .QN(n40) );
  OA22X1 U86 ( .IN1(n66), .IN2(n42), .IN3(n141), .IN4(n38), .Q(n39) );
  NOR2X0 U87 ( .IN1(in2[7]), .IN2(n41), .QN(n46) );
  AO21X1 U88 ( .IN1(in2[7]), .IN2(n41), .IN3(n46), .Q(n47) );
  OA22X1 U89 ( .IN1(n42), .IN2(n130), .IN3(n140), .IN4(n47), .Q(n45) );
  AOI22X1 U90 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n43), .QN(n44) );
  INVX0 U91 ( .INP(in2[8]), .ZN(n51) );
  OA21X1 U92 ( .IN1(n46), .IN2(n51), .IN3(n50), .Q(n52) );
  AOI22X1 U93 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n52), .QN(n49) );
  OA22X1 U94 ( .IN1(n66), .IN2(n51), .IN3(n141), .IN4(n47), .Q(n48) );
  NOR2X0 U95 ( .IN1(in2[9]), .IN2(n50), .QN(n55) );
  AO21X1 U96 ( .IN1(in2[9]), .IN2(n50), .IN3(n55), .Q(n56) );
  OA22X1 U97 ( .IN1(n51), .IN2(n130), .IN3(n140), .IN4(n56), .Q(n54) );
  AOI22X1 U98 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n52), .QN(n53) );
  INVX0 U99 ( .INP(in2[10]), .ZN(n60) );
  OA21X1 U100 ( .IN1(n55), .IN2(n60), .IN3(n59), .Q(n61) );
  AOI22X1 U101 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n61), .QN(n58) );
  OA22X1 U102 ( .IN1(n66), .IN2(n60), .IN3(n141), .IN4(n56), .Q(n57) );
  NOR2X0 U103 ( .IN1(in2[11]), .IN2(n59), .QN(n64) );
  AO21X1 U104 ( .IN1(in2[11]), .IN2(n59), .IN3(n64), .Q(n65) );
  OA22X1 U105 ( .IN1(n60), .IN2(n130), .IN3(n140), .IN4(n65), .Q(n63) );
  AOI22X1 U106 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n61), .QN(n62) );
  INVX0 U107 ( .INP(in2[12]), .ZN(n71) );
  OA21X1 U108 ( .IN1(n64), .IN2(n71), .IN3(n77), .Q(n69) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n69), .QN(n68) );
  OA22X1 U110 ( .IN1(n66), .IN2(n71), .IN3(n141), .IN4(n65), .Q(n67) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n6), .S(n70), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n71), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n7), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n6), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n6), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n8), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n7), .IN4(n85), .IN5(n84), .Q(
        out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n9), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n8), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n8), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n10), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n9), .IN4(n97), .IN5(n96), .Q(
        out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n11), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n10), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n10), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n12), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n11), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n13), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n12), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n12), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n14), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n13), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n15), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n14), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n14), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n15), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_90 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n28), .IN2(n33), .QN(n32) );
  NAND2X0 U4 ( .IN1(n37), .IN2(n42), .QN(n41) );
  NAND2X0 U5 ( .IN1(n46), .IN2(n51), .QN(n50) );
  NAND2X0 U6 ( .IN1(n55), .IN2(n60), .QN(n59) );
  NAND2X0 U7 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U8 ( .IN1(n19), .IN2(n25), .QN(n24) );
  NAND2X0 U9 ( .IN1(n64), .IN2(n71), .QN(n77) );
  NAND2X0 U10 ( .IN1(n81), .IN2(n7), .QN(n89) );
  NAND2X0 U11 ( .IN1(n93), .IN2(n9), .QN(n101) );
  NAND2X0 U12 ( .IN1(n118), .IN2(n13), .QN(n125) );
  NAND2X0 U13 ( .IN1(n105), .IN2(n11), .QN(n114) );
  NAND2X0 U14 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U15 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U16 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U17 ( .IN1(n36), .IN2(n35), .QN(out1[5]) );
  NAND2X0 U18 ( .IN1(n40), .IN2(n39), .QN(out1[6]) );
  NAND2X0 U19 ( .IN1(in1[2]), .IN2(n77), .QN(n70) );
  NAND2X0 U20 ( .IN1(n69), .IN2(n132), .QN(n74) );
  NAND2X0 U21 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U22 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U23 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U24 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U25 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U26 ( .IN1(n17), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U27 ( .IN1(in1[2]), .IN2(n16), .QN(n17) );
  NAND2X0 U28 ( .IN1(n31), .IN2(n30), .QN(out1[4]) );
  NAND2X0 U29 ( .IN1(n27), .IN2(n26), .QN(out1[3]) );
  NAND2X0 U30 ( .IN1(n21), .IN2(n132), .QN(n4) );
  NAND2X0 U31 ( .IN1(n45), .IN2(n44), .QN(out1[7]) );
  NAND2X0 U32 ( .IN1(n49), .IN2(n48), .QN(out1[8]) );
  NAND2X0 U33 ( .IN1(n54), .IN2(n53), .QN(out1[9]) );
  NAND2X0 U34 ( .IN1(n58), .IN2(n57), .QN(out1[10]) );
  NAND2X0 U35 ( .IN1(n63), .IN2(n62), .QN(out1[11]) );
  NAND2X0 U36 ( .IN1(n68), .IN2(n67), .QN(out1[12]) );
  NAND2X0 U37 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U38 ( .IN1(n141), .IN2(n130), .QN(n18) );
  NAND2X0 U39 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NOR2X0 U40 ( .IN1(n22), .IN2(n20), .QN(n3) );
  NOR2X0 U41 ( .IN1(n142), .IN2(n15), .QN(n1) );
  INVX0 U42 ( .INP(n132), .ZN(n141) );
  INVX0 U43 ( .INP(n130), .ZN(n137) );
  NAND3X0 U44 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  NOR2X0 U45 ( .IN1(n142), .IN2(n111), .QN(n138) );
  MUX21X1 U46 ( .IN1(n16), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  NOR3X0 U47 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  INVX0 U48 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U49 ( .INP(in2[13]), .ZN(n6) );
  INVX0 U50 ( .INP(in2[14]), .ZN(n7) );
  INVX0 U51 ( .INP(in2[15]), .ZN(n8) );
  INVX0 U52 ( .INP(in2[16]), .ZN(n9) );
  INVX0 U53 ( .INP(in2[17]), .ZN(n10) );
  INVX0 U54 ( .INP(in2[18]), .ZN(n11) );
  INVX0 U55 ( .INP(in2[19]), .ZN(n12) );
  INVX0 U56 ( .INP(in2[20]), .ZN(n13) );
  INVX0 U57 ( .INP(in2[21]), .ZN(n14) );
  INVX0 U58 ( .INP(in2[22]), .ZN(n15) );
  INVX0 U59 ( .INP(in1[1]), .ZN(n16) );
  INVX0 U60 ( .INP(in1[2]), .ZN(n111) );
  INVX0 U61 ( .INP(n138), .ZN(n140) );
  NOR2X0 U62 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n19) );
  AOI21X1 U63 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n19), .QN(n21) );
  NOR2X0 U64 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U65 ( .IN1(n18), .IN2(in2[0]), .IN3(n138), .IN4(n21), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U66 ( .INP(n133), .ZN(n66) );
  INVX0 U67 ( .INP(in2[2]), .ZN(n25) );
  NOR2X0 U68 ( .IN1(n66), .IN2(n25), .QN(n22) );
  OA21X1 U69 ( .IN1(n19), .IN2(n25), .IN3(n24), .Q(n23) );
  AO22X1 U70 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n23), .Q(n20) );
  AOI22X1 U71 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n23), .QN(n27) );
  NOR2X0 U72 ( .IN1(in2[3]), .IN2(n24), .QN(n28) );
  AO21X1 U73 ( .IN1(in2[3]), .IN2(n24), .IN3(n28), .Q(n29) );
  OA22X1 U74 ( .IN1(n25), .IN2(n130), .IN3(n140), .IN4(n29), .Q(n26) );
  INVX0 U75 ( .INP(in2[4]), .ZN(n33) );
  OA21X1 U76 ( .IN1(n28), .IN2(n33), .IN3(n32), .Q(n34) );
  AOI22X1 U77 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n34), .QN(n31) );
  OA22X1 U78 ( .IN1(n66), .IN2(n33), .IN3(n141), .IN4(n29), .Q(n30) );
  NOR2X0 U79 ( .IN1(in2[5]), .IN2(n32), .QN(n37) );
  AO21X1 U80 ( .IN1(in2[5]), .IN2(n32), .IN3(n37), .Q(n38) );
  OA22X1 U81 ( .IN1(n33), .IN2(n130), .IN3(n140), .IN4(n38), .Q(n36) );
  AOI22X1 U82 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n34), .QN(n35) );
  INVX0 U83 ( .INP(in2[6]), .ZN(n42) );
  OA21X1 U84 ( .IN1(n37), .IN2(n42), .IN3(n41), .Q(n43) );
  AOI22X1 U85 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n43), .QN(n40) );
  OA22X1 U86 ( .IN1(n66), .IN2(n42), .IN3(n141), .IN4(n38), .Q(n39) );
  NOR2X0 U87 ( .IN1(in2[7]), .IN2(n41), .QN(n46) );
  AO21X1 U88 ( .IN1(in2[7]), .IN2(n41), .IN3(n46), .Q(n47) );
  OA22X1 U89 ( .IN1(n42), .IN2(n130), .IN3(n140), .IN4(n47), .Q(n45) );
  AOI22X1 U90 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n43), .QN(n44) );
  INVX0 U91 ( .INP(in2[8]), .ZN(n51) );
  OA21X1 U92 ( .IN1(n46), .IN2(n51), .IN3(n50), .Q(n52) );
  AOI22X1 U93 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n52), .QN(n49) );
  OA22X1 U94 ( .IN1(n66), .IN2(n51), .IN3(n141), .IN4(n47), .Q(n48) );
  NOR2X0 U95 ( .IN1(in2[9]), .IN2(n50), .QN(n55) );
  AO21X1 U96 ( .IN1(in2[9]), .IN2(n50), .IN3(n55), .Q(n56) );
  OA22X1 U97 ( .IN1(n51), .IN2(n130), .IN3(n140), .IN4(n56), .Q(n54) );
  AOI22X1 U98 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n52), .QN(n53) );
  INVX0 U99 ( .INP(in2[10]), .ZN(n60) );
  OA21X1 U100 ( .IN1(n55), .IN2(n60), .IN3(n59), .Q(n61) );
  AOI22X1 U101 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n61), .QN(n58) );
  OA22X1 U102 ( .IN1(n66), .IN2(n60), .IN3(n141), .IN4(n56), .Q(n57) );
  NOR2X0 U103 ( .IN1(in2[11]), .IN2(n59), .QN(n64) );
  AO21X1 U104 ( .IN1(in2[11]), .IN2(n59), .IN3(n64), .Q(n65) );
  OA22X1 U105 ( .IN1(n60), .IN2(n130), .IN3(n140), .IN4(n65), .Q(n63) );
  AOI22X1 U106 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n61), .QN(n62) );
  INVX0 U107 ( .INP(in2[12]), .ZN(n71) );
  OA21X1 U108 ( .IN1(n64), .IN2(n71), .IN3(n77), .Q(n69) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n69), .QN(n68) );
  OA22X1 U110 ( .IN1(n66), .IN2(n71), .IN3(n141), .IN4(n65), .Q(n67) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n6), .S(n70), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n71), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n7), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n6), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n6), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n8), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n7), .IN4(n85), .IN5(n84), .Q(
        out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n9), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n8), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n8), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n10), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n9), .IN4(n97), .IN5(n96), .Q(
        out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n11), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n10), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n10), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n12), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n11), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n13), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n12), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n12), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n14), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n13), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n15), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n14), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n14), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n15), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module mul26_0 ( clk, rst_n, in1, in2, en, mulout );
  input [25:0] in1;
  input [25:0] in2;
  output [50:0] mulout;
  input clk, rst_n, en;
  wire   N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24,
         N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38,
         N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N62, N63,
         N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77,
         N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91,
         N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, n3, n6, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22,
         SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24,
         SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26,
         SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28,
         SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30,
         SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32,
         SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34,
         SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36,
         SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38,
         SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40,
         SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42,
         SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44,
         SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46,
         SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48,
         SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50,
         SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52,
         SYNOPSYS_UNCONNECTED_53, SYNOPSYS_UNCONNECTED_54,
         SYNOPSYS_UNCONNECTED_55, SYNOPSYS_UNCONNECTED_56,
         SYNOPSYS_UNCONNECTED_57, SYNOPSYS_UNCONNECTED_58,
         SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_60,
         SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_62,
         SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_64,
         SYNOPSYS_UNCONNECTED_65, SYNOPSYS_UNCONNECTED_66,
         SYNOPSYS_UNCONNECTED_67, SYNOPSYS_UNCONNECTED_68,
         SYNOPSYS_UNCONNECTED_69, SYNOPSYS_UNCONNECTED_70,
         SYNOPSYS_UNCONNECTED_71, SYNOPSYS_UNCONNECTED_72,
         SYNOPSYS_UNCONNECTED_73, SYNOPSYS_UNCONNECTED_74,
         SYNOPSYS_UNCONNECTED_75, SYNOPSYS_UNCONNECTED_76,
         SYNOPSYS_UNCONNECTED_77, SYNOPSYS_UNCONNECTED_78,
         SYNOPSYS_UNCONNECTED_79, SYNOPSYS_UNCONNECTED_80,
         SYNOPSYS_UNCONNECTED_81, SYNOPSYS_UNCONNECTED_82,
         SYNOPSYS_UNCONNECTED_83, SYNOPSYS_UNCONNECTED_84,
         SYNOPSYS_UNCONNECTED_85, SYNOPSYS_UNCONNECTED_86,
         SYNOPSYS_UNCONNECTED_87, SYNOPSYS_UNCONNECTED_88,
         SYNOPSYS_UNCONNECTED_89, SYNOPSYS_UNCONNECTED_90,
         SYNOPSYS_UNCONNECTED_91, SYNOPSYS_UNCONNECTED_92,
         SYNOPSYS_UNCONNECTED_93, SYNOPSYS_UNCONNECTED_94,
         SYNOPSYS_UNCONNECTED_95, SYNOPSYS_UNCONNECTED_96,
         SYNOPSYS_UNCONNECTED_97, SYNOPSYS_UNCONNECTED_98,
         SYNOPSYS_UNCONNECTED_99, SYNOPSYS_UNCONNECTED_100,
         SYNOPSYS_UNCONNECTED_101, SYNOPSYS_UNCONNECTED_102,
         SYNOPSYS_UNCONNECTED_103, SYNOPSYS_UNCONNECTED_104,
         SYNOPSYS_UNCONNECTED_105, SYNOPSYS_UNCONNECTED_106,
         SYNOPSYS_UNCONNECTED_107, SYNOPSYS_UNCONNECTED_108,
         SYNOPSYS_UNCONNECTED_109, SYNOPSYS_UNCONNECTED_110,
         SYNOPSYS_UNCONNECTED_111, SYNOPSYS_UNCONNECTED_112,
         SYNOPSYS_UNCONNECTED_113, SYNOPSYS_UNCONNECTED_114,
         SYNOPSYS_UNCONNECTED_115, SYNOPSYS_UNCONNECTED_116,
         SYNOPSYS_UNCONNECTED_117, SYNOPSYS_UNCONNECTED_118,
         SYNOPSYS_UNCONNECTED_119, SYNOPSYS_UNCONNECTED_120,
         SYNOPSYS_UNCONNECTED_121, SYNOPSYS_UNCONNECTED_122,
         SYNOPSYS_UNCONNECTED_123, SYNOPSYS_UNCONNECTED_124,
         SYNOPSYS_UNCONNECTED_125, SYNOPSYS_UNCONNECTED_126,
         SYNOPSYS_UNCONNECTED_127, SYNOPSYS_UNCONNECTED_128,
         SYNOPSYS_UNCONNECTED_129, SYNOPSYS_UNCONNECTED_130,
         SYNOPSYS_UNCONNECTED_131, SYNOPSYS_UNCONNECTED_132,
         SYNOPSYS_UNCONNECTED_133, SYNOPSYS_UNCONNECTED_134,
         SYNOPSYS_UNCONNECTED_135, SYNOPSYS_UNCONNECTED_136,
         SYNOPSYS_UNCONNECTED_137, SYNOPSYS_UNCONNECTED_138,
         SYNOPSYS_UNCONNECTED_139, SYNOPSYS_UNCONNECTED_140,
         SYNOPSYS_UNCONNECTED_141, SYNOPSYS_UNCONNECTED_142,
         SYNOPSYS_UNCONNECTED_143, SYNOPSYS_UNCONNECTED_144,
         SYNOPSYS_UNCONNECTED_145, SYNOPSYS_UNCONNECTED_146,
         SYNOPSYS_UNCONNECTED_147, SYNOPSYS_UNCONNECTED_148,
         SYNOPSYS_UNCONNECTED_149, SYNOPSYS_UNCONNECTED_150,
         SYNOPSYS_UNCONNECTED_151, SYNOPSYS_UNCONNECTED_152,
         SYNOPSYS_UNCONNECTED_153, SYNOPSYS_UNCONNECTED_154,
         SYNOPSYS_UNCONNECTED_155, SYNOPSYS_UNCONNECTED_156,
         SYNOPSYS_UNCONNECTED_157, SYNOPSYS_UNCONNECTED_158,
         SYNOPSYS_UNCONNECTED_159, SYNOPSYS_UNCONNECTED_160,
         SYNOPSYS_UNCONNECTED_161, SYNOPSYS_UNCONNECTED_162,
         SYNOPSYS_UNCONNECTED_163, SYNOPSYS_UNCONNECTED_164,
         SYNOPSYS_UNCONNECTED_165, SYNOPSYS_UNCONNECTED_166,
         SYNOPSYS_UNCONNECTED_167, SYNOPSYS_UNCONNECTED_168,
         SYNOPSYS_UNCONNECTED_169, SYNOPSYS_UNCONNECTED_170,
         SYNOPSYS_UNCONNECTED_171, SYNOPSYS_UNCONNECTED_172,
         SYNOPSYS_UNCONNECTED_173, SYNOPSYS_UNCONNECTED_174,
         SYNOPSYS_UNCONNECTED_175, SYNOPSYS_UNCONNECTED_176,
         SYNOPSYS_UNCONNECTED_177, SYNOPSYS_UNCONNECTED_178,
         SYNOPSYS_UNCONNECTED_179, SYNOPSYS_UNCONNECTED_180,
         SYNOPSYS_UNCONNECTED_181, SYNOPSYS_UNCONNECTED_182,
         SYNOPSYS_UNCONNECTED_183, SYNOPSYS_UNCONNECTED_184,
         SYNOPSYS_UNCONNECTED_185, SYNOPSYS_UNCONNECTED_186,
         SYNOPSYS_UNCONNECTED_187, SYNOPSYS_UNCONNECTED_188,
         SYNOPSYS_UNCONNECTED_189, SYNOPSYS_UNCONNECTED_190,
         SYNOPSYS_UNCONNECTED_191, SYNOPSYS_UNCONNECTED_192,
         SYNOPSYS_UNCONNECTED_193, SYNOPSYS_UNCONNECTED_194,
         SYNOPSYS_UNCONNECTED_195, SYNOPSYS_UNCONNECTED_196,
         SYNOPSYS_UNCONNECTED_197, SYNOPSYS_UNCONNECTED_198,
         SYNOPSYS_UNCONNECTED_199, SYNOPSYS_UNCONNECTED_200,
         SYNOPSYS_UNCONNECTED_201, SYNOPSYS_UNCONNECTED_202,
         SYNOPSYS_UNCONNECTED_203, SYNOPSYS_UNCONNECTED_204,
         SYNOPSYS_UNCONNECTED_205, SYNOPSYS_UNCONNECTED_206,
         SYNOPSYS_UNCONNECTED_207, SYNOPSYS_UNCONNECTED_208,
         SYNOPSYS_UNCONNECTED_209, SYNOPSYS_UNCONNECTED_210,
         SYNOPSYS_UNCONNECTED_211, SYNOPSYS_UNCONNECTED_212,
         SYNOPSYS_UNCONNECTED_213, SYNOPSYS_UNCONNECTED_214,
         SYNOPSYS_UNCONNECTED_215, SYNOPSYS_UNCONNECTED_216,
         SYNOPSYS_UNCONNECTED_217, SYNOPSYS_UNCONNECTED_218,
         SYNOPSYS_UNCONNECTED_219, SYNOPSYS_UNCONNECTED_220,
         SYNOPSYS_UNCONNECTED_221, SYNOPSYS_UNCONNECTED_222,
         SYNOPSYS_UNCONNECTED_223, SYNOPSYS_UNCONNECTED_224,
         SYNOPSYS_UNCONNECTED_225, SYNOPSYS_UNCONNECTED_226,
         SYNOPSYS_UNCONNECTED_227, SYNOPSYS_UNCONNECTED_228,
         SYNOPSYS_UNCONNECTED_229, SYNOPSYS_UNCONNECTED_230,
         SYNOPSYS_UNCONNECTED_231, SYNOPSYS_UNCONNECTED_232,
         SYNOPSYS_UNCONNECTED_233, SYNOPSYS_UNCONNECTED_234,
         SYNOPSYS_UNCONNECTED_235, SYNOPSYS_UNCONNECTED_236,
         SYNOPSYS_UNCONNECTED_237, SYNOPSYS_UNCONNECTED_238,
         SYNOPSYS_UNCONNECTED_239, SYNOPSYS_UNCONNECTED_240,
         SYNOPSYS_UNCONNECTED_241, SYNOPSYS_UNCONNECTED_242,
         SYNOPSYS_UNCONNECTED_243, SYNOPSYS_UNCONNECTED_244,
         SYNOPSYS_UNCONNECTED_245, SYNOPSYS_UNCONNECTED_246,
         SYNOPSYS_UNCONNECTED_247, SYNOPSYS_UNCONNECTED_248,
         SYNOPSYS_UNCONNECTED_249, SYNOPSYS_UNCONNECTED_250,
         SYNOPSYS_UNCONNECTED_251, SYNOPSYS_UNCONNECTED_252,
         SYNOPSYS_UNCONNECTED_253, SYNOPSYS_UNCONNECTED_254,
         SYNOPSYS_UNCONNECTED_255, SYNOPSYS_UNCONNECTED_256,
         SYNOPSYS_UNCONNECTED_257, SYNOPSYS_UNCONNECTED_258,
         SYNOPSYS_UNCONNECTED_259, SYNOPSYS_UNCONNECTED_260,
         SYNOPSYS_UNCONNECTED_261, SYNOPSYS_UNCONNECTED_262,
         SYNOPSYS_UNCONNECTED_263, SYNOPSYS_UNCONNECTED_264,
         SYNOPSYS_UNCONNECTED_265, SYNOPSYS_UNCONNECTED_266,
         SYNOPSYS_UNCONNECTED_267, SYNOPSYS_UNCONNECTED_268,
         SYNOPSYS_UNCONNECTED_269, SYNOPSYS_UNCONNECTED_270,
         SYNOPSYS_UNCONNECTED_271, SYNOPSYS_UNCONNECTED_272,
         SYNOPSYS_UNCONNECTED_273, SYNOPSYS_UNCONNECTED_274,
         SYNOPSYS_UNCONNECTED_275, SYNOPSYS_UNCONNECTED_276,
         SYNOPSYS_UNCONNECTED_277, SYNOPSYS_UNCONNECTED_278,
         SYNOPSYS_UNCONNECTED_279, SYNOPSYS_UNCONNECTED_280,
         SYNOPSYS_UNCONNECTED_281, SYNOPSYS_UNCONNECTED_282,
         SYNOPSYS_UNCONNECTED_283, SYNOPSYS_UNCONNECTED_284,
         SYNOPSYS_UNCONNECTED_285, SYNOPSYS_UNCONNECTED_286,
         SYNOPSYS_UNCONNECTED_287, SYNOPSYS_UNCONNECTED_288,
         SYNOPSYS_UNCONNECTED_289, SYNOPSYS_UNCONNECTED_290,
         SYNOPSYS_UNCONNECTED_291, SYNOPSYS_UNCONNECTED_292,
         SYNOPSYS_UNCONNECTED_293, SYNOPSYS_UNCONNECTED_294,
         SYNOPSYS_UNCONNECTED_295, SYNOPSYS_UNCONNECTED_296,
         SYNOPSYS_UNCONNECTED_297, SYNOPSYS_UNCONNECTED_298,
         SYNOPSYS_UNCONNECTED_299, SYNOPSYS_UNCONNECTED_300,
         SYNOPSYS_UNCONNECTED_301, SYNOPSYS_UNCONNECTED_302,
         SYNOPSYS_UNCONNECTED_303, SYNOPSYS_UNCONNECTED_304,
         SYNOPSYS_UNCONNECTED_305, SYNOPSYS_UNCONNECTED_306,
         SYNOPSYS_UNCONNECTED_307, SYNOPSYS_UNCONNECTED_308,
         SYNOPSYS_UNCONNECTED_309, SYNOPSYS_UNCONNECTED_310,
         SYNOPSYS_UNCONNECTED_311, SYNOPSYS_UNCONNECTED_312,
         SYNOPSYS_UNCONNECTED_313, SYNOPSYS_UNCONNECTED_314,
         SYNOPSYS_UNCONNECTED_315, SYNOPSYS_UNCONNECTED_316,
         SYNOPSYS_UNCONNECTED_317, SYNOPSYS_UNCONNECTED_318,
         SYNOPSYS_UNCONNECTED_319, SYNOPSYS_UNCONNECTED_320,
         SYNOPSYS_UNCONNECTED_321, SYNOPSYS_UNCONNECTED_322,
         SYNOPSYS_UNCONNECTED_323, SYNOPSYS_UNCONNECTED_324,
         SYNOPSYS_UNCONNECTED_325, SYNOPSYS_UNCONNECTED_326,
         SYNOPSYS_UNCONNECTED_327, SYNOPSYS_UNCONNECTED_328,
         SYNOPSYS_UNCONNECTED_329, SYNOPSYS_UNCONNECTED_330,
         SYNOPSYS_UNCONNECTED_331, SYNOPSYS_UNCONNECTED_332,
         SYNOPSYS_UNCONNECTED_333, SYNOPSYS_UNCONNECTED_334,
         SYNOPSYS_UNCONNECTED_335, SYNOPSYS_UNCONNECTED_336,
         SYNOPSYS_UNCONNECTED_337, SYNOPSYS_UNCONNECTED_338,
         SYNOPSYS_UNCONNECTED_339, SYNOPSYS_UNCONNECTED_340,
         SYNOPSYS_UNCONNECTED_341, SYNOPSYS_UNCONNECTED_342,
         SYNOPSYS_UNCONNECTED_343, SYNOPSYS_UNCONNECTED_344,
         SYNOPSYS_UNCONNECTED_345, SYNOPSYS_UNCONNECTED_346,
         SYNOPSYS_UNCONNECTED_347, SYNOPSYS_UNCONNECTED_348,
         SYNOPSYS_UNCONNECTED_349, SYNOPSYS_UNCONNECTED_350,
         SYNOPSYS_UNCONNECTED_351, SYNOPSYS_UNCONNECTED_352,
         SYNOPSYS_UNCONNECTED_353, SYNOPSYS_UNCONNECTED_354,
         SYNOPSYS_UNCONNECTED_355, SYNOPSYS_UNCONNECTED_356,
         SYNOPSYS_UNCONNECTED_357, SYNOPSYS_UNCONNECTED_358,
         SYNOPSYS_UNCONNECTED_359, SYNOPSYS_UNCONNECTED_360,
         SYNOPSYS_UNCONNECTED_361, SYNOPSYS_UNCONNECTED_362,
         SYNOPSYS_UNCONNECTED_363, SYNOPSYS_UNCONNECTED_364,
         SYNOPSYS_UNCONNECTED_365, SYNOPSYS_UNCONNECTED_366,
         SYNOPSYS_UNCONNECTED_367, SYNOPSYS_UNCONNECTED_368,
         SYNOPSYS_UNCONNECTED_369, SYNOPSYS_UNCONNECTED_370,
         SYNOPSYS_UNCONNECTED_371, SYNOPSYS_UNCONNECTED_372,
         SYNOPSYS_UNCONNECTED_373, SYNOPSYS_UNCONNECTED_374,
         SYNOPSYS_UNCONNECTED_375, SYNOPSYS_UNCONNECTED_376,
         SYNOPSYS_UNCONNECTED_377, SYNOPSYS_UNCONNECTED_378,
         SYNOPSYS_UNCONNECTED_379, SYNOPSYS_UNCONNECTED_380,
         SYNOPSYS_UNCONNECTED_381, SYNOPSYS_UNCONNECTED_382,
         SYNOPSYS_UNCONNECTED_383, SYNOPSYS_UNCONNECTED_384,
         SYNOPSYS_UNCONNECTED_385, SYNOPSYS_UNCONNECTED_386,
         SYNOPSYS_UNCONNECTED_387, SYNOPSYS_UNCONNECTED_388,
         SYNOPSYS_UNCONNECTED_389, SYNOPSYS_UNCONNECTED_390,
         SYNOPSYS_UNCONNECTED_391, SYNOPSYS_UNCONNECTED_392,
         SYNOPSYS_UNCONNECTED_393, SYNOPSYS_UNCONNECTED_394,
         SYNOPSYS_UNCONNECTED_395, SYNOPSYS_UNCONNECTED_396,
         SYNOPSYS_UNCONNECTED_397, SYNOPSYS_UNCONNECTED_398,
         SYNOPSYS_UNCONNECTED_399, SYNOPSYS_UNCONNECTED_400,
         SYNOPSYS_UNCONNECTED_401, SYNOPSYS_UNCONNECTED_402,
         SYNOPSYS_UNCONNECTED_403, SYNOPSYS_UNCONNECTED_404,
         SYNOPSYS_UNCONNECTED_405, SYNOPSYS_UNCONNECTED_406,
         SYNOPSYS_UNCONNECTED_407, SYNOPSYS_UNCONNECTED_408,
         SYNOPSYS_UNCONNECTED_409, SYNOPSYS_UNCONNECTED_410,
         SYNOPSYS_UNCONNECTED_411, SYNOPSYS_UNCONNECTED_412;
  wire   [26:2] boothout1;
  wire   [26:0] boothout2;
  wire   [26:0] boothout3;
  wire   [26:0] boothout4;
  wire   [26:0] boothout5;
  wire   [26:0] boothout6;
  wire   [26:0] boothout7;
  wire   [26:0] boothout8;
  wire   [26:0] boothout9;
  wire   [26:0] boothout10;
  wire   [26:0] boothout11;
  wire   [25:0] boothout12;
  wire   [22:0] boothout13;
  wire   [29:2] cout1;
  wire   [31:3] mulout1;
  wire   [35:8] cout2;
  wire   [37:6] mulout2;
  wire   [41:14] cout3;
  wire   [42:12] mulout3;
  wire   [46:20] cout4;
  wire   [47:18] mulout4;
  wire   [31:3] cout5;
  wire   [46:4] mulout5;
  wire   [37:9] cout6;
  wire   [42:6] mulout6;
  wire   [46:18] cout7;
  wire   [47:12] mulout7;
  wire   [38:4] cout8;
  wire   [46:5] mulout8;
  wire   [46:12] cout9;
  wire   [47:6] mulout9;
  wire   [46:5] cout10;
  wire   [47:6] mulout10;
  wire   [46:6] cout11;
  wire   [47:7] mulout11;
  wire   [47:0] a;
  wire   [47:8] b;

  booth27_0 booth1 ( .out1({boothout1, SYNOPSYS_UNCONNECTED_1, 
        SYNOPSYS_UNCONNECTED_2}), .in1({in1[1:0], 1'b0}), .in2({1'b0, 1'b0, 
        1'b1, in2[22:0]}) );
  booth27_90 booth2 ( .out1(boothout2), .in1(in1[3:1]), .in2({1'b0, 1'b0, 1'b1, 
        in2[22:0]}) );
  booth27_89 booth3 ( .out1(boothout3), .in1(in1[5:3]), .in2({1'b0, 1'b0, 1'b1, 
        in2[22:0]}) );
  booth27_88 booth4 ( .out1(boothout4), .in1(in1[7:5]), .in2({1'b0, 1'b0, 1'b1, 
        in2[22:0]}) );
  booth27_87 booth5 ( .out1(boothout5), .in1(in1[9:7]), .in2({1'b0, 1'b0, 1'b1, 
        in2[22:0]}) );
  booth27_86 booth6 ( .out1(boothout6), .in1(in1[11:9]), .in2({1'b0, 1'b0, 
        1'b1, in2[22:0]}) );
  booth27_85 booth7 ( .out1(boothout7), .in1(in1[13:11]), .in2({1'b0, 1'b0, 
        1'b1, in2[22:0]}) );
  booth27_84 booth8 ( .out1(boothout8), .in1(in1[15:13]), .in2({1'b0, 1'b0, 
        1'b1, in2[22:0]}) );
  booth27_83 booth9 ( .out1(boothout9), .in1(in1[17:15]), .in2({1'b0, 1'b0, 
        1'b1, in2[22:0]}) );
  booth27_82 booth10 ( .out1(boothout10), .in1(in1[19:17]), .in2({1'b0, 1'b0, 
        1'b1, in2[22:0]}) );
  booth27_81 booth11 ( .out1(boothout11), .in1(in1[21:19]), .in2({1'b0, 1'b0, 
        1'b1, in2[22:0]}) );
  booth27_80 booth12 ( .out1({SYNOPSYS_UNCONNECTED_3, boothout12}), .in1({1'b1, 
        in1[22:21]}), .in2({1'b0, 1'b0, 1'b1, in2[22:0]}) );
  booth27_79 booth13 ( .out1({SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, 
        SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, boothout13}), .in1({
        1'b0, 1'b0, 1'b1}), .in2({1'b0, 1'b0, 1'b1, in2[22:0]}) );
  csa51squ_0 csa51squ1 ( .cout({SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, 
        SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11, 
        SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13, 
        SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, 
        SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17, 
        SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19, 
        SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21, 
        SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_23, 
        SYNOPSYS_UNCONNECTED_24, SYNOPSYS_UNCONNECTED_25, 
        SYNOPSYS_UNCONNECTED_26, SYNOPSYS_UNCONNECTED_27, 
        SYNOPSYS_UNCONNECTED_28, cout1, SYNOPSYS_UNCONNECTED_29, 
        SYNOPSYS_UNCONNECTED_30}), .sumout({SYNOPSYS_UNCONNECTED_31, 
        SYNOPSYS_UNCONNECTED_32, SYNOPSYS_UNCONNECTED_33, 
        SYNOPSYS_UNCONNECTED_34, SYNOPSYS_UNCONNECTED_35, 
        SYNOPSYS_UNCONNECTED_36, SYNOPSYS_UNCONNECTED_37, 
        SYNOPSYS_UNCONNECTED_38, SYNOPSYS_UNCONNECTED_39, 
        SYNOPSYS_UNCONNECTED_40, SYNOPSYS_UNCONNECTED_41, 
        SYNOPSYS_UNCONNECTED_42, SYNOPSYS_UNCONNECTED_43, 
        SYNOPSYS_UNCONNECTED_44, SYNOPSYS_UNCONNECTED_45, 
        SYNOPSYS_UNCONNECTED_46, SYNOPSYS_UNCONNECTED_47, 
        SYNOPSYS_UNCONNECTED_48, SYNOPSYS_UNCONNECTED_49, mulout1[31], 
        SYNOPSYS_UNCONNECTED_50, mulout1[29:3], SYNOPSYS_UNCONNECTED_51, 
        SYNOPSYS_UNCONNECTED_52, SYNOPSYS_UNCONNECTED_53}), .in1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, boothout1, 
        1'b0, 1'b0}), .in2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, boothout2, 1'b0, 1'b0}), .in3({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, n3, 1'b0, boothout3[25:0], 1'b0, 1'b0, 1'b0, 1'b0})
         );
  csa51squ_83 csa51squ2 ( .cout({SYNOPSYS_UNCONNECTED_54, 
        SYNOPSYS_UNCONNECTED_55, SYNOPSYS_UNCONNECTED_56, 
        SYNOPSYS_UNCONNECTED_57, SYNOPSYS_UNCONNECTED_58, 
        SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_60, 
        SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_62, 
        SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_64, 
        SYNOPSYS_UNCONNECTED_65, SYNOPSYS_UNCONNECTED_66, 
        SYNOPSYS_UNCONNECTED_67, SYNOPSYS_UNCONNECTED_68, cout2, 
        SYNOPSYS_UNCONNECTED_69, SYNOPSYS_UNCONNECTED_70, 
        SYNOPSYS_UNCONNECTED_71, SYNOPSYS_UNCONNECTED_72, 
        SYNOPSYS_UNCONNECTED_73, SYNOPSYS_UNCONNECTED_74, 
        SYNOPSYS_UNCONNECTED_75, SYNOPSYS_UNCONNECTED_76}), .sumout({
        SYNOPSYS_UNCONNECTED_77, SYNOPSYS_UNCONNECTED_78, 
        SYNOPSYS_UNCONNECTED_79, SYNOPSYS_UNCONNECTED_80, 
        SYNOPSYS_UNCONNECTED_81, SYNOPSYS_UNCONNECTED_82, 
        SYNOPSYS_UNCONNECTED_83, SYNOPSYS_UNCONNECTED_84, 
        SYNOPSYS_UNCONNECTED_85, SYNOPSYS_UNCONNECTED_86, 
        SYNOPSYS_UNCONNECTED_87, SYNOPSYS_UNCONNECTED_88, 
        SYNOPSYS_UNCONNECTED_89, mulout2[37], SYNOPSYS_UNCONNECTED_90, 
        mulout2[35:6], SYNOPSYS_UNCONNECTED_91, SYNOPSYS_UNCONNECTED_92, 
        SYNOPSYS_UNCONNECTED_93, SYNOPSYS_UNCONNECTED_94, 
        SYNOPSYS_UNCONNECTED_95, SYNOPSYS_UNCONNECTED_96}), .in1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, boothout4, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, boothout5, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .in3({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n6, 1'b0, boothout6[25:0], 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_82 csa51squ3 ( .cout({SYNOPSYS_UNCONNECTED_97, 
        SYNOPSYS_UNCONNECTED_98, SYNOPSYS_UNCONNECTED_99, 
        SYNOPSYS_UNCONNECTED_100, SYNOPSYS_UNCONNECTED_101, 
        SYNOPSYS_UNCONNECTED_102, SYNOPSYS_UNCONNECTED_103, 
        SYNOPSYS_UNCONNECTED_104, SYNOPSYS_UNCONNECTED_105, cout3, 
        SYNOPSYS_UNCONNECTED_106, SYNOPSYS_UNCONNECTED_107, 
        SYNOPSYS_UNCONNECTED_108, SYNOPSYS_UNCONNECTED_109, 
        SYNOPSYS_UNCONNECTED_110, SYNOPSYS_UNCONNECTED_111, 
        SYNOPSYS_UNCONNECTED_112, SYNOPSYS_UNCONNECTED_113, 
        SYNOPSYS_UNCONNECTED_114, SYNOPSYS_UNCONNECTED_115, 
        SYNOPSYS_UNCONNECTED_116, SYNOPSYS_UNCONNECTED_117, 
        SYNOPSYS_UNCONNECTED_118, SYNOPSYS_UNCONNECTED_119}), .sumout({
        SYNOPSYS_UNCONNECTED_120, SYNOPSYS_UNCONNECTED_121, 
        SYNOPSYS_UNCONNECTED_122, SYNOPSYS_UNCONNECTED_123, 
        SYNOPSYS_UNCONNECTED_124, SYNOPSYS_UNCONNECTED_125, 
        SYNOPSYS_UNCONNECTED_126, SYNOPSYS_UNCONNECTED_127, mulout3, 
        SYNOPSYS_UNCONNECTED_128, SYNOPSYS_UNCONNECTED_129, 
        SYNOPSYS_UNCONNECTED_130, SYNOPSYS_UNCONNECTED_131, 
        SYNOPSYS_UNCONNECTED_132, SYNOPSYS_UNCONNECTED_133, 
        SYNOPSYS_UNCONNECTED_134, SYNOPSYS_UNCONNECTED_135, 
        SYNOPSYS_UNCONNECTED_136, SYNOPSYS_UNCONNECTED_137, 
        SYNOPSYS_UNCONNECTED_138, SYNOPSYS_UNCONNECTED_139}), .in1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, boothout7, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, boothout8, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .in3({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        boothout9, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_81 csa51squ4 ( .cout({SYNOPSYS_UNCONNECTED_140, 
        SYNOPSYS_UNCONNECTED_141, SYNOPSYS_UNCONNECTED_142, 
        SYNOPSYS_UNCONNECTED_143, cout4, SYNOPSYS_UNCONNECTED_144, 
        SYNOPSYS_UNCONNECTED_145, SYNOPSYS_UNCONNECTED_146, 
        SYNOPSYS_UNCONNECTED_147, SYNOPSYS_UNCONNECTED_148, 
        SYNOPSYS_UNCONNECTED_149, SYNOPSYS_UNCONNECTED_150, 
        SYNOPSYS_UNCONNECTED_151, SYNOPSYS_UNCONNECTED_152, 
        SYNOPSYS_UNCONNECTED_153, SYNOPSYS_UNCONNECTED_154, 
        SYNOPSYS_UNCONNECTED_155, SYNOPSYS_UNCONNECTED_156, 
        SYNOPSYS_UNCONNECTED_157, SYNOPSYS_UNCONNECTED_158, 
        SYNOPSYS_UNCONNECTED_159, SYNOPSYS_UNCONNECTED_160, 
        SYNOPSYS_UNCONNECTED_161, SYNOPSYS_UNCONNECTED_162, 
        SYNOPSYS_UNCONNECTED_163}), .sumout({SYNOPSYS_UNCONNECTED_164, 
        SYNOPSYS_UNCONNECTED_165, SYNOPSYS_UNCONNECTED_166, mulout4, 
        SYNOPSYS_UNCONNECTED_167, SYNOPSYS_UNCONNECTED_168, 
        SYNOPSYS_UNCONNECTED_169, SYNOPSYS_UNCONNECTED_170, 
        SYNOPSYS_UNCONNECTED_171, SYNOPSYS_UNCONNECTED_172, 
        SYNOPSYS_UNCONNECTED_173, SYNOPSYS_UNCONNECTED_174, 
        SYNOPSYS_UNCONNECTED_175, SYNOPSYS_UNCONNECTED_176, 
        SYNOPSYS_UNCONNECTED_177, SYNOPSYS_UNCONNECTED_178, 
        SYNOPSYS_UNCONNECTED_179, SYNOPSYS_UNCONNECTED_180, 
        SYNOPSYS_UNCONNECTED_181, SYNOPSYS_UNCONNECTED_182, 
        SYNOPSYS_UNCONNECTED_183, SYNOPSYS_UNCONNECTED_184}), .in1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, boothout10, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 1'b0, 1'b0, 1'b0, boothout11, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .in3({1'b0, 1'b0, 1'b0, boothout12, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_80 csa51squ5 ( .cout({SYNOPSYS_UNCONNECTED_185, 
        SYNOPSYS_UNCONNECTED_186, SYNOPSYS_UNCONNECTED_187, 
        SYNOPSYS_UNCONNECTED_188, SYNOPSYS_UNCONNECTED_189, 
        SYNOPSYS_UNCONNECTED_190, SYNOPSYS_UNCONNECTED_191, 
        SYNOPSYS_UNCONNECTED_192, SYNOPSYS_UNCONNECTED_193, 
        SYNOPSYS_UNCONNECTED_194, SYNOPSYS_UNCONNECTED_195, 
        SYNOPSYS_UNCONNECTED_196, SYNOPSYS_UNCONNECTED_197, 
        SYNOPSYS_UNCONNECTED_198, SYNOPSYS_UNCONNECTED_199, 
        SYNOPSYS_UNCONNECTED_200, SYNOPSYS_UNCONNECTED_201, 
        SYNOPSYS_UNCONNECTED_202, SYNOPSYS_UNCONNECTED_203, cout5, 
        SYNOPSYS_UNCONNECTED_204, SYNOPSYS_UNCONNECTED_205, 
        SYNOPSYS_UNCONNECTED_206}), .sumout({SYNOPSYS_UNCONNECTED_207, 
        SYNOPSYS_UNCONNECTED_208, SYNOPSYS_UNCONNECTED_209, 
        SYNOPSYS_UNCONNECTED_210, mulout5, SYNOPSYS_UNCONNECTED_211, 
        SYNOPSYS_UNCONNECTED_212, SYNOPSYS_UNCONNECTED_213, 
        SYNOPSYS_UNCONNECTED_214}), .in1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, cout1, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, mulout1[31], 1'b0, mulout1[29:3], 1'b0, 1'b0, 1'b0}), 
        .in3({1'b0, 1'b0, 1'b0, 1'b1, boothout13, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_79 csa51squ6 ( .cout({SYNOPSYS_UNCONNECTED_215, 
        SYNOPSYS_UNCONNECTED_216, SYNOPSYS_UNCONNECTED_217, 
        SYNOPSYS_UNCONNECTED_218, SYNOPSYS_UNCONNECTED_219, 
        SYNOPSYS_UNCONNECTED_220, SYNOPSYS_UNCONNECTED_221, 
        SYNOPSYS_UNCONNECTED_222, SYNOPSYS_UNCONNECTED_223, 
        SYNOPSYS_UNCONNECTED_224, SYNOPSYS_UNCONNECTED_225, 
        SYNOPSYS_UNCONNECTED_226, SYNOPSYS_UNCONNECTED_227, cout6, 
        SYNOPSYS_UNCONNECTED_228, SYNOPSYS_UNCONNECTED_229, 
        SYNOPSYS_UNCONNECTED_230, SYNOPSYS_UNCONNECTED_231, 
        SYNOPSYS_UNCONNECTED_232, SYNOPSYS_UNCONNECTED_233, 
        SYNOPSYS_UNCONNECTED_234, SYNOPSYS_UNCONNECTED_235, 
        SYNOPSYS_UNCONNECTED_236}), .sumout({SYNOPSYS_UNCONNECTED_237, 
        SYNOPSYS_UNCONNECTED_238, SYNOPSYS_UNCONNECTED_239, 
        SYNOPSYS_UNCONNECTED_240, SYNOPSYS_UNCONNECTED_241, 
        SYNOPSYS_UNCONNECTED_242, SYNOPSYS_UNCONNECTED_243, 
        SYNOPSYS_UNCONNECTED_244, mulout6, SYNOPSYS_UNCONNECTED_245, 
        SYNOPSYS_UNCONNECTED_246, SYNOPSYS_UNCONNECTED_247, 
        SYNOPSYS_UNCONNECTED_248, SYNOPSYS_UNCONNECTED_249, 
        SYNOPSYS_UNCONNECTED_250}), .in1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, cout2, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        mulout2[37], 1'b0, mulout2[35:6], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .in3({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, cout3, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  csa51squ_78 csa51squ7 ( .cout({SYNOPSYS_UNCONNECTED_251, 
        SYNOPSYS_UNCONNECTED_252, SYNOPSYS_UNCONNECTED_253, 
        SYNOPSYS_UNCONNECTED_254, cout7, SYNOPSYS_UNCONNECTED_255, 
        SYNOPSYS_UNCONNECTED_256, SYNOPSYS_UNCONNECTED_257, 
        SYNOPSYS_UNCONNECTED_258, SYNOPSYS_UNCONNECTED_259, 
        SYNOPSYS_UNCONNECTED_260, SYNOPSYS_UNCONNECTED_261, 
        SYNOPSYS_UNCONNECTED_262, SYNOPSYS_UNCONNECTED_263, 
        SYNOPSYS_UNCONNECTED_264, SYNOPSYS_UNCONNECTED_265, 
        SYNOPSYS_UNCONNECTED_266, SYNOPSYS_UNCONNECTED_267, 
        SYNOPSYS_UNCONNECTED_268, SYNOPSYS_UNCONNECTED_269, 
        SYNOPSYS_UNCONNECTED_270, SYNOPSYS_UNCONNECTED_271, 
        SYNOPSYS_UNCONNECTED_272}), .sumout({SYNOPSYS_UNCONNECTED_273, 
        SYNOPSYS_UNCONNECTED_274, SYNOPSYS_UNCONNECTED_275, mulout7, 
        SYNOPSYS_UNCONNECTED_276, SYNOPSYS_UNCONNECTED_277, 
        SYNOPSYS_UNCONNECTED_278, SYNOPSYS_UNCONNECTED_279, 
        SYNOPSYS_UNCONNECTED_280, SYNOPSYS_UNCONNECTED_281, 
        SYNOPSYS_UNCONNECTED_282, SYNOPSYS_UNCONNECTED_283, 
        SYNOPSYS_UNCONNECTED_284, SYNOPSYS_UNCONNECTED_285, 
        SYNOPSYS_UNCONNECTED_286, SYNOPSYS_UNCONNECTED_287}), .in1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mulout3, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 1'b0, 
        1'b0, cout4, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in3({1'b0, 1'b0, 1'b0, mulout4, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_77 csa51squ8 ( .cout({SYNOPSYS_UNCONNECTED_288, 
        SYNOPSYS_UNCONNECTED_289, SYNOPSYS_UNCONNECTED_290, 
        SYNOPSYS_UNCONNECTED_291, SYNOPSYS_UNCONNECTED_292, 
        SYNOPSYS_UNCONNECTED_293, SYNOPSYS_UNCONNECTED_294, 
        SYNOPSYS_UNCONNECTED_295, SYNOPSYS_UNCONNECTED_296, 
        SYNOPSYS_UNCONNECTED_297, SYNOPSYS_UNCONNECTED_298, 
        SYNOPSYS_UNCONNECTED_299, cout8, SYNOPSYS_UNCONNECTED_300, 
        SYNOPSYS_UNCONNECTED_301, SYNOPSYS_UNCONNECTED_302, 
        SYNOPSYS_UNCONNECTED_303}), .sumout({SYNOPSYS_UNCONNECTED_304, 
        SYNOPSYS_UNCONNECTED_305, SYNOPSYS_UNCONNECTED_306, 
        SYNOPSYS_UNCONNECTED_307, mulout8, SYNOPSYS_UNCONNECTED_308, 
        SYNOPSYS_UNCONNECTED_309, SYNOPSYS_UNCONNECTED_310, 
        SYNOPSYS_UNCONNECTED_311, SYNOPSYS_UNCONNECTED_312}), .in1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, cout5, 1'b0, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 
        1'b0, 1'b0, 1'b1, mulout5, 1'b0, 1'b0, 1'b0, 1'b0}), .in3({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, cout6, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_76 csa51squ9 ( .cout({SYNOPSYS_UNCONNECTED_313, 
        SYNOPSYS_UNCONNECTED_314, SYNOPSYS_UNCONNECTED_315, 
        SYNOPSYS_UNCONNECTED_316, cout9, SYNOPSYS_UNCONNECTED_317, 
        SYNOPSYS_UNCONNECTED_318, SYNOPSYS_UNCONNECTED_319, 
        SYNOPSYS_UNCONNECTED_320, SYNOPSYS_UNCONNECTED_321, 
        SYNOPSYS_UNCONNECTED_322, SYNOPSYS_UNCONNECTED_323, 
        SYNOPSYS_UNCONNECTED_324, SYNOPSYS_UNCONNECTED_325, 
        SYNOPSYS_UNCONNECTED_326, SYNOPSYS_UNCONNECTED_327, 
        SYNOPSYS_UNCONNECTED_328}), .sumout({SYNOPSYS_UNCONNECTED_329, 
        SYNOPSYS_UNCONNECTED_330, SYNOPSYS_UNCONNECTED_331, mulout9, 
        SYNOPSYS_UNCONNECTED_332, SYNOPSYS_UNCONNECTED_333, 
        SYNOPSYS_UNCONNECTED_334, SYNOPSYS_UNCONNECTED_335, 
        SYNOPSYS_UNCONNECTED_336, SYNOPSYS_UNCONNECTED_337}), .in1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mulout6, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .in2({1'b0, 1'b0, 1'b0, cout7, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .in3({1'b0, 1'b0, 1'b0, mulout7, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_75 csa51squ10 ( .cout({SYNOPSYS_UNCONNECTED_338, 
        SYNOPSYS_UNCONNECTED_339, SYNOPSYS_UNCONNECTED_340, 
        SYNOPSYS_UNCONNECTED_341, cout10, SYNOPSYS_UNCONNECTED_342, 
        SYNOPSYS_UNCONNECTED_343, SYNOPSYS_UNCONNECTED_344, 
        SYNOPSYS_UNCONNECTED_345, SYNOPSYS_UNCONNECTED_346}), .sumout({
        SYNOPSYS_UNCONNECTED_347, SYNOPSYS_UNCONNECTED_348, 
        SYNOPSYS_UNCONNECTED_349, mulout10, SYNOPSYS_UNCONNECTED_350, 
        SYNOPSYS_UNCONNECTED_351, SYNOPSYS_UNCONNECTED_352, 
        SYNOPSYS_UNCONNECTED_353, SYNOPSYS_UNCONNECTED_354, 
        SYNOPSYS_UNCONNECTED_355}), .in1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, cout8, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .in2({1'b0, 1'b0, 1'b0, 1'b1, mulout8, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .in3({1'b0, 1'b0, 1'b0, cout9, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_74 csa51squ11 ( .cout({SYNOPSYS_UNCONNECTED_356, 
        SYNOPSYS_UNCONNECTED_357, SYNOPSYS_UNCONNECTED_358, 
        SYNOPSYS_UNCONNECTED_359, cout11, SYNOPSYS_UNCONNECTED_360, 
        SYNOPSYS_UNCONNECTED_361, SYNOPSYS_UNCONNECTED_362, 
        SYNOPSYS_UNCONNECTED_363, SYNOPSYS_UNCONNECTED_364, 
        SYNOPSYS_UNCONNECTED_365}), .sumout({SYNOPSYS_UNCONNECTED_366, 
        SYNOPSYS_UNCONNECTED_367, SYNOPSYS_UNCONNECTED_368, mulout11, 
        SYNOPSYS_UNCONNECTED_369, SYNOPSYS_UNCONNECTED_370, 
        SYNOPSYS_UNCONNECTED_371, SYNOPSYS_UNCONNECTED_372, 
        SYNOPSYS_UNCONNECTED_373, SYNOPSYS_UNCONNECTED_374, 
        SYNOPSYS_UNCONNECTED_375}), .in1({1'b0, 1'b0, 1'b0, mulout9, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 1'b0, 1'b0, cout10, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in3({1'b0, 1'b0, 1'b0, mulout10, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_73 csa51squ12 ( .sumout({SYNOPSYS_UNCONNECTED_376, 
        SYNOPSYS_UNCONNECTED_377, SYNOPSYS_UNCONNECTED_378, N101, N100, N99, 
        N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, 
        N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, 
        N70, N69, N68, N67, N66, N65, N64, N63, N62, SYNOPSYS_UNCONNECTED_379, 
        SYNOPSYS_UNCONNECTED_380, SYNOPSYS_UNCONNECTED_381, 
        SYNOPSYS_UNCONNECTED_382, SYNOPSYS_UNCONNECTED_383, 
        SYNOPSYS_UNCONNECTED_384, SYNOPSYS_UNCONNECTED_385, 
        SYNOPSYS_UNCONNECTED_386}), .in1({1'b0, 1'b0, 1'b0, mulout11, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 1'b0, 1'b0, cout11, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in3({1'b1, 1'b0, 1'b1, 
        1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 
        1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .cout_46_(N50), .cout_44_(N48), .cout_42_(N46), .cout_40_(N44), .cout_38_(
        N42), .cout_36_(N40), .cout_34_(N38), .cout_32_(N36), .cout_30_(N34), 
        .cout_28_(N32), .cout_27_(N31), .cout_7__BAR(N11), .cout_8__BAR(N12), 
        .cout_9__BAR(N13), .cout_10__BAR(N14), .cout_11__BAR(N15), 
        .cout_12__BAR(N16), .cout_13__BAR(N17), .cout_14__BAR(N18), 
        .cout_15__BAR(N19), .cout_16__BAR(N20), .cout_17__BAR(N21), 
        .cout_18__BAR(N22), .cout_19__BAR(N23), .cout_20__BAR(N24), 
        .cout_21__BAR(N25), .cout_22__BAR(N26), .cout_23__BAR(N27), 
        .cout_24__BAR(N28), .cout_25__BAR(N29), .cout_26__BAR(N30), 
        .cout_29__BAR(N33), .cout_31__BAR(N35), .cout_33__BAR(N37), 
        .cout_35__BAR(N39), .cout_37__BAR(N41), .cout_39__BAR(N43), 
        .cout_41__BAR(N45), .cout_43__BAR(N47), .cout_45__BAR(N49) );
  cla51squ_0 cla51squ ( .out({SYNOPSYS_UNCONNECTED_387, 
        SYNOPSYS_UNCONNECTED_388, SYNOPSYS_UNCONNECTED_389, mulout[47:23], 
        SYNOPSYS_UNCONNECTED_390, SYNOPSYS_UNCONNECTED_391, 
        SYNOPSYS_UNCONNECTED_392, SYNOPSYS_UNCONNECTED_393, 
        SYNOPSYS_UNCONNECTED_394, SYNOPSYS_UNCONNECTED_395, 
        SYNOPSYS_UNCONNECTED_396, SYNOPSYS_UNCONNECTED_397, 
        SYNOPSYS_UNCONNECTED_398, SYNOPSYS_UNCONNECTED_399, 
        SYNOPSYS_UNCONNECTED_400, SYNOPSYS_UNCONNECTED_401, 
        SYNOPSYS_UNCONNECTED_402, SYNOPSYS_UNCONNECTED_403, 
        SYNOPSYS_UNCONNECTED_404, SYNOPSYS_UNCONNECTED_405, 
        SYNOPSYS_UNCONNECTED_406, SYNOPSYS_UNCONNECTED_407, 
        SYNOPSYS_UNCONNECTED_408, SYNOPSYS_UNCONNECTED_409, 
        SYNOPSYS_UNCONNECTED_410, SYNOPSYS_UNCONNECTED_411, 
        SYNOPSYS_UNCONNECTED_412}), .a({1'b0, 1'b0, 1'b0, a[47:8], 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({1'b0, 1'b0, 1'b0, b, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  DFFARX1 b_reg_47_ ( .D(N101), .CLK(clk), .RSTB(rst_n), .Q(b[47]) );
  DFFARX1 b_reg_46_ ( .D(N100), .CLK(clk), .RSTB(rst_n), .Q(b[46]) );
  DFFARX1 b_reg_45_ ( .D(N99), .CLK(clk), .RSTB(rst_n), .Q(b[45]) );
  DFFARX1 b_reg_44_ ( .D(N98), .CLK(clk), .RSTB(rst_n), .Q(b[44]) );
  DFFARX1 b_reg_43_ ( .D(N97), .CLK(clk), .RSTB(rst_n), .Q(b[43]) );
  DFFARX1 b_reg_42_ ( .D(N96), .CLK(clk), .RSTB(rst_n), .Q(b[42]) );
  DFFARX1 b_reg_41_ ( .D(N95), .CLK(clk), .RSTB(rst_n), .Q(b[41]) );
  DFFARX1 b_reg_40_ ( .D(N94), .CLK(clk), .RSTB(rst_n), .Q(b[40]) );
  DFFARX1 b_reg_39_ ( .D(N93), .CLK(clk), .RSTB(rst_n), .Q(b[39]) );
  DFFARX1 b_reg_38_ ( .D(N92), .CLK(clk), .RSTB(rst_n), .Q(b[38]) );
  DFFARX1 b_reg_37_ ( .D(N91), .CLK(clk), .RSTB(rst_n), .Q(b[37]) );
  DFFARX1 b_reg_36_ ( .D(N90), .CLK(clk), .RSTB(rst_n), .Q(b[36]) );
  DFFARX1 b_reg_35_ ( .D(N89), .CLK(clk), .RSTB(rst_n), .Q(b[35]) );
  DFFARX1 b_reg_34_ ( .D(N88), .CLK(clk), .RSTB(rst_n), .Q(b[34]) );
  DFFARX1 b_reg_33_ ( .D(N87), .CLK(clk), .RSTB(rst_n), .Q(b[33]) );
  DFFARX1 b_reg_32_ ( .D(N86), .CLK(clk), .RSTB(rst_n), .Q(b[32]) );
  DFFARX1 b_reg_31_ ( .D(N85), .CLK(clk), .RSTB(rst_n), .Q(b[31]) );
  DFFARX1 b_reg_30_ ( .D(N84), .CLK(clk), .RSTB(rst_n), .Q(b[30]) );
  DFFARX1 b_reg_29_ ( .D(N83), .CLK(clk), .RSTB(rst_n), .Q(b[29]) );
  DFFARX1 b_reg_28_ ( .D(N82), .CLK(clk), .RSTB(rst_n), .Q(b[28]) );
  DFFARX1 b_reg_27_ ( .D(N81), .CLK(clk), .RSTB(rst_n), .Q(b[27]) );
  DFFARX1 b_reg_26_ ( .D(N80), .CLK(clk), .RSTB(rst_n), .Q(b[26]) );
  DFFARX1 b_reg_25_ ( .D(N79), .CLK(clk), .RSTB(rst_n), .Q(b[25]) );
  DFFARX1 b_reg_24_ ( .D(N78), .CLK(clk), .RSTB(rst_n), .Q(b[24]) );
  DFFARX1 b_reg_23_ ( .D(N77), .CLK(clk), .RSTB(rst_n), .Q(b[23]) );
  DFFARX1 b_reg_22_ ( .D(N76), .CLK(clk), .RSTB(rst_n), .Q(b[22]) );
  DFFARX1 b_reg_21_ ( .D(N75), .CLK(clk), .RSTB(rst_n), .Q(b[21]) );
  DFFARX1 b_reg_20_ ( .D(N74), .CLK(clk), .RSTB(rst_n), .Q(b[20]) );
  DFFARX1 b_reg_19_ ( .D(N73), .CLK(clk), .RSTB(rst_n), .Q(b[19]) );
  DFFARX1 b_reg_18_ ( .D(N72), .CLK(clk), .RSTB(rst_n), .Q(b[18]) );
  DFFARX1 b_reg_17_ ( .D(N71), .CLK(clk), .RSTB(rst_n), .Q(b[17]) );
  DFFARX1 b_reg_16_ ( .D(N70), .CLK(clk), .RSTB(rst_n), .Q(b[16]) );
  DFFARX1 b_reg_15_ ( .D(N69), .CLK(clk), .RSTB(rst_n), .Q(b[15]) );
  DFFARX1 b_reg_14_ ( .D(N68), .CLK(clk), .RSTB(rst_n), .Q(b[14]) );
  DFFARX1 b_reg_13_ ( .D(N67), .CLK(clk), .RSTB(rst_n), .Q(b[13]) );
  DFFARX1 b_reg_12_ ( .D(N66), .CLK(clk), .RSTB(rst_n), .Q(b[12]) );
  DFFARX1 b_reg_11_ ( .D(N65), .CLK(clk), .RSTB(rst_n), .Q(b[11]) );
  DFFARX1 b_reg_10_ ( .D(N64), .CLK(clk), .RSTB(rst_n), .Q(b[10]) );
  DFFARX1 b_reg_9_ ( .D(N63), .CLK(clk), .RSTB(rst_n), .Q(b[9]) );
  DFFARX1 b_reg_8_ ( .D(N62), .CLK(clk), .RSTB(rst_n), .Q(b[8]) );
  DFFARX1 a_reg_47_ ( .D(N50), .CLK(clk), .RSTB(rst_n), .Q(a[47]) );
  DFFARX1 a_reg_46_ ( .D(n45), .CLK(clk), .RSTB(rst_n), .Q(a[46]) );
  DFFARX1 a_reg_45_ ( .D(N48), .CLK(clk), .RSTB(rst_n), .Q(a[45]) );
  DFFARX1 a_reg_44_ ( .D(n46), .CLK(clk), .RSTB(rst_n), .Q(a[44]) );
  DFFARX1 a_reg_43_ ( .D(N46), .CLK(clk), .RSTB(rst_n), .Q(a[43]) );
  DFFARX1 a_reg_42_ ( .D(n47), .CLK(clk), .RSTB(rst_n), .Q(a[42]) );
  DFFARX1 a_reg_41_ ( .D(N44), .CLK(clk), .RSTB(rst_n), .Q(a[41]) );
  DFFARX1 a_reg_40_ ( .D(n48), .CLK(clk), .RSTB(rst_n), .Q(a[40]) );
  DFFARX1 a_reg_39_ ( .D(N42), .CLK(clk), .RSTB(rst_n), .Q(a[39]) );
  DFFARX1 a_reg_38_ ( .D(n49), .CLK(clk), .RSTB(rst_n), .Q(a[38]) );
  DFFARX1 a_reg_37_ ( .D(N40), .CLK(clk), .RSTB(rst_n), .Q(a[37]) );
  DFFARX1 a_reg_36_ ( .D(n50), .CLK(clk), .RSTB(rst_n), .Q(a[36]) );
  DFFARX1 a_reg_35_ ( .D(N38), .CLK(clk), .RSTB(rst_n), .Q(a[35]) );
  DFFARX1 a_reg_34_ ( .D(n51), .CLK(clk), .RSTB(rst_n), .Q(a[34]) );
  DFFARX1 a_reg_33_ ( .D(N36), .CLK(clk), .RSTB(rst_n), .Q(a[33]) );
  DFFARX1 a_reg_32_ ( .D(n52), .CLK(clk), .RSTB(rst_n), .Q(a[32]) );
  DFFARX1 a_reg_31_ ( .D(N34), .CLK(clk), .RSTB(rst_n), .Q(a[31]) );
  DFFARX1 a_reg_30_ ( .D(n53), .CLK(clk), .RSTB(rst_n), .Q(a[30]) );
  DFFARX1 a_reg_29_ ( .D(N32), .CLK(clk), .RSTB(rst_n), .Q(a[29]) );
  DFFARX1 a_reg_28_ ( .D(N31), .CLK(clk), .RSTB(rst_n), .Q(a[28]) );
  DFFARX1 a_reg_27_ ( .D(n54), .CLK(clk), .RSTB(rst_n), .Q(a[27]) );
  DFFARX1 a_reg_26_ ( .D(n55), .CLK(clk), .RSTB(rst_n), .Q(a[26]) );
  DFFARX1 a_reg_25_ ( .D(n56), .CLK(clk), .RSTB(rst_n), .Q(a[25]) );
  DFFARX1 a_reg_24_ ( .D(n57), .CLK(clk), .RSTB(rst_n), .Q(a[24]) );
  DFFARX1 a_reg_23_ ( .D(n58), .CLK(clk), .RSTB(rst_n), .Q(a[23]) );
  DFFARX1 a_reg_22_ ( .D(n59), .CLK(clk), .RSTB(rst_n), .Q(a[22]) );
  DFFARX1 a_reg_21_ ( .D(n60), .CLK(clk), .RSTB(rst_n), .Q(a[21]) );
  DFFARX1 a_reg_20_ ( .D(n61), .CLK(clk), .RSTB(rst_n), .Q(a[20]) );
  DFFARX1 a_reg_19_ ( .D(n62), .CLK(clk), .RSTB(rst_n), .Q(a[19]) );
  DFFARX1 a_reg_18_ ( .D(n63), .CLK(clk), .RSTB(rst_n), .Q(a[18]) );
  DFFARX1 a_reg_17_ ( .D(n64), .CLK(clk), .RSTB(rst_n), .Q(a[17]) );
  DFFARX1 a_reg_16_ ( .D(n65), .CLK(clk), .RSTB(rst_n), .Q(a[16]) );
  DFFARX1 a_reg_15_ ( .D(n66), .CLK(clk), .RSTB(rst_n), .Q(a[15]) );
  DFFARX1 a_reg_14_ ( .D(n67), .CLK(clk), .RSTB(rst_n), .Q(a[14]) );
  DFFARX1 a_reg_13_ ( .D(n68), .CLK(clk), .RSTB(rst_n), .Q(a[13]) );
  DFFARX1 a_reg_12_ ( .D(n69), .CLK(clk), .RSTB(rst_n), .Q(a[12]) );
  DFFARX1 a_reg_11_ ( .D(n70), .CLK(clk), .RSTB(rst_n), .Q(a[11]) );
  DFFARX1 a_reg_10_ ( .D(n71), .CLK(clk), .RSTB(rst_n), .Q(a[10]) );
  DFFARX1 a_reg_9_ ( .D(n72), .CLK(clk), .RSTB(rst_n), .Q(a[9]) );
  DFFARX1 a_reg_8_ ( .D(n73), .CLK(clk), .RSTB(rst_n), .Q(a[8]) );
  INVX0 U5 ( .INP(boothout3[26]), .ZN(n3) );
  INVX0 U8 ( .INP(boothout6[26]), .ZN(n6) );
  INVX0 U54 ( .INP(N49), .ZN(n45) );
  INVX0 U55 ( .INP(N47), .ZN(n46) );
  INVX0 U56 ( .INP(N45), .ZN(n47) );
  INVX0 U57 ( .INP(N43), .ZN(n48) );
  INVX0 U58 ( .INP(N41), .ZN(n49) );
  INVX0 U59 ( .INP(N39), .ZN(n50) );
  INVX0 U60 ( .INP(N37), .ZN(n51) );
  INVX0 U61 ( .INP(N35), .ZN(n52) );
  INVX0 U62 ( .INP(N33), .ZN(n53) );
  INVX0 U63 ( .INP(N30), .ZN(n54) );
  INVX0 U64 ( .INP(N29), .ZN(n55) );
  INVX0 U65 ( .INP(N28), .ZN(n56) );
  INVX0 U66 ( .INP(N27), .ZN(n57) );
  INVX0 U67 ( .INP(N26), .ZN(n58) );
  INVX0 U68 ( .INP(N25), .ZN(n59) );
  INVX0 U69 ( .INP(N24), .ZN(n60) );
  INVX0 U70 ( .INP(N23), .ZN(n61) );
  INVX0 U71 ( .INP(N22), .ZN(n62) );
  INVX0 U72 ( .INP(N21), .ZN(n63) );
  INVX0 U73 ( .INP(N20), .ZN(n64) );
  INVX0 U74 ( .INP(N19), .ZN(n65) );
  INVX0 U75 ( .INP(N18), .ZN(n66) );
  INVX0 U76 ( .INP(N17), .ZN(n67) );
  INVX0 U77 ( .INP(N16), .ZN(n68) );
  INVX0 U78 ( .INP(N15), .ZN(n69) );
  INVX0 U79 ( .INP(N14), .ZN(n70) );
  INVX0 U80 ( .INP(N13), .ZN(n71) );
  INVX0 U81 ( .INP(N12), .ZN(n72) );
  INVX0 U82 ( .INP(N11), .ZN(n73) );
endmodule


module add_0 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(b), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(b), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_777 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  XOR3X1 U1 ( .IN1(b), .IN2(ci), .IN3(a), .Q(s) );
endmodule


module add_778 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_779 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_780 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_781 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_782 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_783 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module adder8_0 ( out, a, b, cin );
  output [7:0] out;
  input [7:0] a;
  input [7:0] b;
  input cin;

  wire   [6:0] c;

  add_0 add_01 ( .s(out[0]), .a(a[0]), .b(b[0]), .ci(1'b0), .co(c[0]) );
  add_783 add_02 ( .s(out[1]), .a(a[1]), .b(b[1]), .ci(c[0]), .co(c[1]) );
  add_782 add_03 ( .s(out[2]), .a(a[2]), .b(b[2]), .ci(c[1]), .co(c[2]) );
  add_781 add_04 ( .s(out[3]), .a(a[3]), .b(b[3]), .ci(c[2]), .co(c[3]) );
  add_780 add_05 ( .s(out[4]), .a(a[4]), .b(b[4]), .ci(c[3]), .co(c[4]) );
  add_779 add_06 ( .s(out[5]), .a(a[5]), .b(b[5]), .ci(c[4]), .co(c[5]) );
  add_778 add_07 ( .s(out[6]), .a(a[6]), .b(b[6]), .ci(c[5]), .co(c[6]) );
  add_777 add_08 ( .s(out[7]), .a(a[7]), .b(b[7]), .ci(c[6]) );
endmodule


module add_769 ( s, a, b, co, ci_BAR );
  input a, b, ci_BAR;
  output s, co;


  XOR2X1 U1 ( .IN1(a), .IN2(ci_BAR), .Q(s) );
endmodule


module add_770 ( s, a, b, ci, co_BAR );
  input a, b, ci;
  output s, co_BAR;


  NAND2X0 U1 ( .IN1(ci), .IN2(a), .QN(co_BAR) );
  OA21X1 U2 ( .IN1(ci), .IN2(a), .IN3(co_BAR), .Q(s) );
endmodule


module add_771 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_772 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_773 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_774 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_775 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  INVX0 U1 ( .INP(a), .ZN(s) );
  NBUFFX2 U2 ( .INP(a), .Z(co) );
endmodule


module add_776 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  NBUFFX2 U1 ( .INP(a), .Z(s) );
endmodule


module adder8_55 ( out, a, b, cin );
  output [7:0] out;
  input [7:0] a;
  input [7:0] b;
  input cin;

  wire   [6:1] c;

  add_776 add_01 ( .s(out[0]), .a(a[0]), .b(1'b1), .ci(1'b1) );
  add_775 add_02 ( .s(out[1]), .a(a[1]), .b(1'b0), .ci(1'b1), .co(c[1]) );
  add_774 add_03 ( .s(out[2]), .a(a[2]), .b(1'b0), .ci(c[1]), .co(c[2]) );
  add_773 add_04 ( .s(out[3]), .a(a[3]), .b(1'b0), .ci(c[2]), .co(c[3]) );
  add_772 add_05 ( .s(out[4]), .a(a[4]), .b(1'b0), .ci(c[3]), .co(c[4]) );
  add_771 add_06 ( .s(out[5]), .a(a[5]), .b(1'b0), .ci(c[4]), .co(c[5]) );
  add_770 add_07 ( .s(out[6]), .a(a[6]), .b(1'b0), .ci(c[5]), .co_BAR(c[6]) );
  add_769 add_08 ( .s(out[7]), .a(a[7]), .b(1'b1), .ci_BAR(c[6]) );
endmodule


module floating_point_multiple_0 ( clk, rst_n, input_factor_01, 
        input_factor_02, output_multiply );
  input [31:0] input_factor_01;
  input [31:0] input_factor_02;
  output [31:0] output_multiply;
  input clk, rst_n;
  wire   N5, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22,
         N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N48, N49, N50, N51,
         N52, N53, N54, N55, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22,
         SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24,
         SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26;
  wire   [47:23] base_multiply_result;
  wire   [47:23] mulout;
  wire   [7:0] exponent_factor_12;
  wire   [7:0] pre_mul_output_exponent;

  mul26_0 mul26_01 ( .clk(clk), .rst_n(rst_n), .in1({1'b0, 1'b0, 1'b1, 
        input_factor_01[22:0]}), .in2({1'b0, 1'b0, 1'b1, input_factor_02[22:0]}), .en(1'b1), .mulout({SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, 
        SYNOPSYS_UNCONNECTED_3, mulout, SYNOPSYS_UNCONNECTED_4, 
        SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, 
        SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, 
        SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11, 
        SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13, 
        SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, 
        SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17, 
        SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19, 
        SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21, 
        SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_23, 
        SYNOPSYS_UNCONNECTED_24, SYNOPSYS_UNCONNECTED_25, 
        SYNOPSYS_UNCONNECTED_26}) );
  adder8_0 adder8_01 ( .out(exponent_factor_12), .a(input_factor_01[30:23]), 
        .b(input_factor_02[30:23]), .cin(1'b0) );
  adder8_55 adder8_02 ( .out(pre_mul_output_exponent), .a(exponent_factor_12), 
        .b({1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0}), .cin(1'b1) );
  DFFARX1 mul_output_sign_reg ( .D(N5), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[31]) );
  DFFARX1 base_multiply_result_reg_47_ ( .D(mulout[47]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[47]) );
  DFFARX1 base_multiply_result_reg_46_ ( .D(mulout[46]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[46]) );
  DFFARX1 base_multiply_result_reg_45_ ( .D(mulout[45]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[45]) );
  DFFARX1 base_multiply_result_reg_44_ ( .D(mulout[44]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[44]) );
  DFFARX1 base_multiply_result_reg_43_ ( .D(mulout[43]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[43]) );
  DFFARX1 base_multiply_result_reg_42_ ( .D(mulout[42]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[42]) );
  DFFARX1 base_multiply_result_reg_41_ ( .D(mulout[41]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[41]) );
  DFFARX1 base_multiply_result_reg_40_ ( .D(mulout[40]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[40]) );
  DFFARX1 base_multiply_result_reg_39_ ( .D(mulout[39]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[39]) );
  DFFARX1 base_multiply_result_reg_38_ ( .D(mulout[38]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[38]) );
  DFFARX1 base_multiply_result_reg_37_ ( .D(mulout[37]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[37]) );
  DFFARX1 base_multiply_result_reg_36_ ( .D(mulout[36]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[36]) );
  DFFARX1 base_multiply_result_reg_35_ ( .D(mulout[35]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[35]) );
  DFFARX1 base_multiply_result_reg_34_ ( .D(mulout[34]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[34]) );
  DFFARX1 base_multiply_result_reg_33_ ( .D(mulout[33]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[33]) );
  DFFARX1 base_multiply_result_reg_32_ ( .D(mulout[32]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[32]) );
  DFFARX1 base_multiply_result_reg_31_ ( .D(mulout[31]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[31]) );
  DFFARX1 base_multiply_result_reg_30_ ( .D(mulout[30]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[30]) );
  DFFARX1 base_multiply_result_reg_29_ ( .D(mulout[29]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[29]) );
  DFFARX1 base_multiply_result_reg_28_ ( .D(mulout[28]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[28]) );
  DFFARX1 base_multiply_result_reg_27_ ( .D(mulout[27]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[27]) );
  DFFARX1 base_multiply_result_reg_26_ ( .D(mulout[26]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[26]) );
  DFFARX1 base_multiply_result_reg_25_ ( .D(mulout[25]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[25]) );
  DFFARX1 base_multiply_result_reg_24_ ( .D(mulout[24]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[24]) );
  DFFARX1 base_multiply_result_reg_23_ ( .D(mulout[23]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[23]) );
  DFFARX1 mul_output_significand_reg_22_ ( .D(N32), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[22]) );
  DFFARX1 mul_output_significand_reg_21_ ( .D(N31), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[21]) );
  DFFARX1 mul_output_significand_reg_20_ ( .D(N30), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[20]) );
  DFFARX1 mul_output_significand_reg_19_ ( .D(N29), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[19]) );
  DFFARX1 mul_output_significand_reg_18_ ( .D(N28), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[18]) );
  DFFARX1 mul_output_significand_reg_17_ ( .D(N27), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[17]) );
  DFFARX1 mul_output_significand_reg_16_ ( .D(N26), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[16]) );
  DFFARX1 mul_output_significand_reg_15_ ( .D(N25), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[15]) );
  DFFARX1 mul_output_significand_reg_14_ ( .D(N24), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[14]) );
  DFFARX1 mul_output_significand_reg_13_ ( .D(N23), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[13]) );
  DFFARX1 mul_output_significand_reg_12_ ( .D(N22), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[12]) );
  DFFARX1 mul_output_significand_reg_11_ ( .D(N21), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[11]) );
  DFFARX1 mul_output_significand_reg_10_ ( .D(N20), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[10]) );
  DFFARX1 mul_output_significand_reg_9_ ( .D(N19), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[9]) );
  DFFARX1 mul_output_significand_reg_8_ ( .D(N18), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[8]) );
  DFFARX1 mul_output_significand_reg_7_ ( .D(N17), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[7]) );
  DFFARX1 mul_output_significand_reg_6_ ( .D(N16), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[6]) );
  DFFARX1 mul_output_significand_reg_5_ ( .D(N15), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[5]) );
  DFFARX1 mul_output_significand_reg_4_ ( .D(N14), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[4]) );
  DFFARX1 mul_output_significand_reg_3_ ( .D(N13), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[3]) );
  DFFARX1 mul_output_significand_reg_2_ ( .D(N12), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[2]) );
  DFFARX1 mul_output_significand_reg_1_ ( .D(N11), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[1]) );
  DFFARX1 mul_output_significand_reg_0_ ( .D(N10), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[0]) );
  DFFARX1 mul_output_exponent_reg_7_ ( .D(N55), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[30]) );
  DFFARX1 mul_output_exponent_reg_6_ ( .D(N54), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[29]) );
  DFFARX1 mul_output_exponent_reg_5_ ( .D(N53), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[28]) );
  DFFARX1 mul_output_exponent_reg_4_ ( .D(N52), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[27]) );
  DFFARX1 mul_output_exponent_reg_3_ ( .D(N51), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[26]) );
  DFFARX1 mul_output_exponent_reg_2_ ( .D(N50), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[25]) );
  DFFARX1 mul_output_exponent_reg_1_ ( .D(N49), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[24]) );
  DFFARX1 mul_output_exponent_reg_0_ ( .D(N48), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[23]) );
  AND2X1 U3 ( .IN1(base_multiply_result[47]), .IN2(n35), .Q(n32) );
  INVX0 U4 ( .INP(n1), .ZN(n2) );
  OR2X1 U5 ( .IN1(base_multiply_result[47]), .IN2(n23), .Q(n1) );
  NOR4X0 U6 ( .IN1(input_factor_01[0]), .IN2(input_factor_01[10]), .IN3(
        input_factor_01[11]), .IN4(input_factor_01[12]), .QN(n6) );
  NOR4X0 U7 ( .IN1(input_factor_01[13]), .IN2(input_factor_01[14]), .IN3(
        input_factor_01[15]), .IN4(input_factor_01[16]), .QN(n5) );
  NOR4X0 U8 ( .IN1(input_factor_01[17]), .IN2(input_factor_01[18]), .IN3(
        input_factor_01[19]), .IN4(input_factor_01[1]), .QN(n4) );
  NOR4X0 U9 ( .IN1(input_factor_01[20]), .IN2(input_factor_01[21]), .IN3(
        input_factor_01[22]), .IN4(input_factor_01[23]), .QN(n3) );
  NAND4X0 U10 ( .IN1(n6), .IN2(n5), .IN3(n4), .IN4(n3), .QN(n22) );
  NOR4X0 U11 ( .IN1(input_factor_01[24]), .IN2(input_factor_01[25]), .IN3(
        input_factor_01[26]), .IN4(input_factor_01[27]), .QN(n10) );
  NOR4X0 U12 ( .IN1(input_factor_01[28]), .IN2(input_factor_01[29]), .IN3(
        input_factor_01[2]), .IN4(input_factor_01[30]), .QN(n9) );
  NOR4X0 U13 ( .IN1(input_factor_01[31]), .IN2(input_factor_01[3]), .IN3(
        input_factor_01[4]), .IN4(input_factor_01[5]), .QN(n8) );
  NOR4X0 U14 ( .IN1(input_factor_01[6]), .IN2(input_factor_01[7]), .IN3(
        input_factor_01[8]), .IN4(input_factor_01[9]), .QN(n7) );
  NAND4X0 U15 ( .IN1(n10), .IN2(n9), .IN3(n8), .IN4(n7), .QN(n21) );
  NOR4X0 U16 ( .IN1(input_factor_02[0]), .IN2(input_factor_02[10]), .IN3(
        input_factor_02[11]), .IN4(input_factor_02[12]), .QN(n14) );
  NOR4X0 U17 ( .IN1(input_factor_02[13]), .IN2(input_factor_02[14]), .IN3(
        input_factor_02[15]), .IN4(input_factor_02[16]), .QN(n13) );
  NOR4X0 U18 ( .IN1(input_factor_02[17]), .IN2(input_factor_02[18]), .IN3(
        input_factor_02[19]), .IN4(input_factor_02[1]), .QN(n12) );
  NOR4X0 U19 ( .IN1(input_factor_02[20]), .IN2(input_factor_02[21]), .IN3(
        input_factor_02[22]), .IN4(input_factor_02[23]), .QN(n11) );
  NAND4X0 U20 ( .IN1(n14), .IN2(n13), .IN3(n12), .IN4(n11), .QN(n20) );
  NOR4X0 U21 ( .IN1(input_factor_02[24]), .IN2(input_factor_02[25]), .IN3(
        input_factor_02[26]), .IN4(input_factor_02[27]), .QN(n18) );
  NOR4X0 U22 ( .IN1(input_factor_02[28]), .IN2(input_factor_02[29]), .IN3(
        input_factor_02[2]), .IN4(input_factor_02[30]), .QN(n17) );
  NOR4X0 U23 ( .IN1(input_factor_02[31]), .IN2(input_factor_02[3]), .IN3(
        input_factor_02[4]), .IN4(input_factor_02[5]), .QN(n16) );
  NOR4X0 U24 ( .IN1(input_factor_02[6]), .IN2(input_factor_02[7]), .IN3(
        input_factor_02[8]), .IN4(input_factor_02[9]), .QN(n15) );
  NAND4X0 U25 ( .IN1(n18), .IN2(n17), .IN3(n16), .IN4(n15), .QN(n19) );
  OA22X1 U26 ( .IN1(n22), .IN2(n21), .IN3(n20), .IN4(n19), .Q(n35) );
  INVX0 U27 ( .INP(n35), .ZN(n23) );
  AO22X1 U28 ( .IN1(n2), .IN2(base_multiply_result[23]), .IN3(n32), .IN4(
        base_multiply_result[24]), .Q(N10) );
  AO22X1 U29 ( .IN1(n2), .IN2(base_multiply_result[24]), .IN3(n32), .IN4(
        base_multiply_result[25]), .Q(N11) );
  AO22X1 U30 ( .IN1(n2), .IN2(base_multiply_result[25]), .IN3(n32), .IN4(
        base_multiply_result[26]), .Q(N12) );
  AO22X1 U31 ( .IN1(n2), .IN2(base_multiply_result[26]), .IN3(n32), .IN4(
        base_multiply_result[27]), .Q(N13) );
  AO22X1 U32 ( .IN1(n2), .IN2(base_multiply_result[27]), .IN3(n32), .IN4(
        base_multiply_result[28]), .Q(N14) );
  AO22X1 U33 ( .IN1(n2), .IN2(base_multiply_result[28]), .IN3(n32), .IN4(
        base_multiply_result[29]), .Q(N15) );
  AO22X1 U34 ( .IN1(n2), .IN2(base_multiply_result[29]), .IN3(n32), .IN4(
        base_multiply_result[30]), .Q(N16) );
  AO22X1 U35 ( .IN1(n2), .IN2(base_multiply_result[30]), .IN3(n32), .IN4(
        base_multiply_result[31]), .Q(N17) );
  AO22X1 U36 ( .IN1(n2), .IN2(base_multiply_result[31]), .IN3(n32), .IN4(
        base_multiply_result[32]), .Q(N18) );
  AO22X1 U37 ( .IN1(n2), .IN2(base_multiply_result[32]), .IN3(n32), .IN4(
        base_multiply_result[33]), .Q(N19) );
  AO22X1 U38 ( .IN1(n2), .IN2(base_multiply_result[33]), .IN3(n32), .IN4(
        base_multiply_result[34]), .Q(N20) );
  AO22X1 U39 ( .IN1(n2), .IN2(base_multiply_result[34]), .IN3(n32), .IN4(
        base_multiply_result[35]), .Q(N21) );
  AO22X1 U40 ( .IN1(n2), .IN2(base_multiply_result[35]), .IN3(n32), .IN4(
        base_multiply_result[36]), .Q(N22) );
  AO22X1 U41 ( .IN1(n2), .IN2(base_multiply_result[36]), .IN3(n32), .IN4(
        base_multiply_result[37]), .Q(N23) );
  AO22X1 U42 ( .IN1(n2), .IN2(base_multiply_result[37]), .IN3(n32), .IN4(
        base_multiply_result[38]), .Q(N24) );
  AO22X1 U43 ( .IN1(n2), .IN2(base_multiply_result[38]), .IN3(n32), .IN4(
        base_multiply_result[39]), .Q(N25) );
  AO22X1 U44 ( .IN1(n2), .IN2(base_multiply_result[39]), .IN3(n32), .IN4(
        base_multiply_result[40]), .Q(N26) );
  AO22X1 U45 ( .IN1(n2), .IN2(base_multiply_result[40]), .IN3(n32), .IN4(
        base_multiply_result[41]), .Q(N27) );
  AO22X1 U46 ( .IN1(n2), .IN2(base_multiply_result[41]), .IN3(n32), .IN4(
        base_multiply_result[42]), .Q(N28) );
  AO22X1 U47 ( .IN1(n2), .IN2(base_multiply_result[42]), .IN3(n32), .IN4(
        base_multiply_result[43]), .Q(N29) );
  AO22X1 U48 ( .IN1(n2), .IN2(base_multiply_result[43]), .IN3(n32), .IN4(
        base_multiply_result[44]), .Q(N30) );
  AO22X1 U49 ( .IN1(n2), .IN2(base_multiply_result[44]), .IN3(n32), .IN4(
        base_multiply_result[45]), .Q(N31) );
  AO22X1 U50 ( .IN1(n2), .IN2(base_multiply_result[45]), .IN3(n32), .IN4(
        base_multiply_result[46]), .Q(N32) );
  MUX21X1 U51 ( .IN1(n2), .IN2(n32), .S(pre_mul_output_exponent[0]), .Q(N48)
         );
  AO21X1 U52 ( .IN1(pre_mul_output_exponent[0]), .IN2(n2), .IN3(n32), .Q(n24)
         );
  NOR3X0 U53 ( .IN1(pre_mul_output_exponent[1]), .IN2(
        pre_mul_output_exponent[0]), .IN3(n1), .QN(n27) );
  AO21X1 U54 ( .IN1(pre_mul_output_exponent[1]), .IN2(n24), .IN3(n27), .Q(N49)
         );
  INVX0 U55 ( .INP(input_factor_01[31]), .ZN(n26) );
  INVX0 U56 ( .INP(input_factor_02[31]), .ZN(n25) );
  OA221X1 U57 ( .IN1(input_factor_01[31]), .IN2(input_factor_02[31]), .IN3(n26), .IN4(n25), .IN5(n35), .Q(N5) );
  AO221X1 U58 ( .IN1(n2), .IN2(pre_mul_output_exponent[1]), .IN3(n2), .IN4(
        pre_mul_output_exponent[0]), .IN5(n32), .Q(n28) );
  MUX21X1 U59 ( .IN1(n27), .IN2(n28), .S(pre_mul_output_exponent[2]), .Q(N50)
         );
  AND2X1 U60 ( .IN1(n2), .IN2(pre_mul_output_exponent[2]), .Q(n29) );
  OR4X1 U61 ( .IN1(pre_mul_output_exponent[1]), .IN2(
        pre_mul_output_exponent[0]), .IN3(pre_mul_output_exponent[3]), .IN4(
        pre_mul_output_exponent[2]), .Q(n34) );
  NOR2X0 U62 ( .IN1(n1), .IN2(n34), .QN(n31) );
  AO221X1 U63 ( .IN1(pre_mul_output_exponent[3]), .IN2(n29), .IN3(
        pre_mul_output_exponent[3]), .IN4(n28), .IN5(n31), .Q(N51) );
  OA21X1 U64 ( .IN1(base_multiply_result[47]), .IN2(n34), .IN3(n35), .Q(n30)
         );
  MUX21X1 U65 ( .IN1(n31), .IN2(n30), .S(pre_mul_output_exponent[4]), .Q(N52)
         );
  AO221X1 U66 ( .IN1(n2), .IN2(pre_mul_output_exponent[4]), .IN3(n2), .IN4(n34), .IN5(n32), .Q(n33) );
  NOR4X0 U67 ( .IN1(pre_mul_output_exponent[5]), .IN2(
        pre_mul_output_exponent[4]), .IN3(n34), .IN4(n1), .QN(n37) );
  AO21X1 U68 ( .IN1(pre_mul_output_exponent[5]), .IN2(n33), .IN3(n37), .Q(N53)
         );
  OR3X1 U69 ( .IN1(pre_mul_output_exponent[5]), .IN2(
        pre_mul_output_exponent[4]), .IN3(n34), .Q(n36) );
  OA21X1 U70 ( .IN1(base_multiply_result[47]), .IN2(n36), .IN3(n35), .Q(n39)
         );
  INVX0 U71 ( .INP(n37), .ZN(n38) );
  NOR2X0 U72 ( .IN1(pre_mul_output_exponent[6]), .IN2(n38), .QN(n41) );
  AO21X1 U73 ( .IN1(pre_mul_output_exponent[6]), .IN2(n39), .IN3(n41), .Q(N54)
         );
  AO21X1 U74 ( .IN1(n2), .IN2(pre_mul_output_exponent[6]), .IN3(n39), .Q(n40)
         );
  MUX21X1 U75 ( .IN1(n41), .IN2(n40), .S(pre_mul_output_exponent[7]), .Q(N55)
         );
endmodule


module add_729 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_730 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_731 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_732 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_733 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_734 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_735 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_736 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_737 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_738 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_739 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_740 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_741 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_742 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_743 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_744 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_745 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_746 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_747 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_748 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_749 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_750 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_751 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_752 ( s, a, ci, co, b_BAR );
  input a, ci, b_BAR;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(b_BAR), .IN2(n1), .QN(co) );
  INVX0 U2 ( .INP(a), .ZN(n1) );
  MUX21X1 U3 ( .IN1(a), .IN2(n1), .S(b_BAR), .Q(s) );
endmodule


module adder24_0 ( clk, rst_n, a, b, cin, out );
  input [23:0] a;
  input [23:0] b;
  output [24:0] out;
  input clk, rst_n, cin;
  wire   c_tmp, n_1_net_, n_2_net_, n_3_net_, n_4_net_, n_5_net_, n_6_net_,
         n_7_net_, n_8_net_, n_9_net_, n_10_net_, n_11_net_, n_12_net_,
         n_13_net_, n_14_net_, n_15_net_, n_16_net_, n_17_net_, n_18_net_,
         n_19_net_, n_20_net_, n_21_net_, n_22_net_, n_23_net_;
  wire   [24:0] s;
  wire   [23:0] c;

  add_752 add_01 ( .s(s[0]), .a(a[0]), .ci(1'b1), .co(c[0]), .b_BAR(b[0]) );
  add_751 add_02 ( .s(s[1]), .a(a[1]), .b(n_1_net_), .ci(c[0]), .co(c[1]) );
  add_750 add_03 ( .s(s[2]), .a(a[2]), .b(n_2_net_), .ci(c[1]), .co(c[2]) );
  add_749 add_04 ( .s(s[3]), .a(a[3]), .b(n_3_net_), .ci(c[2]), .co(c[3]) );
  add_748 add_05 ( .s(s[4]), .a(a[4]), .b(n_4_net_), .ci(c[3]), .co(c[4]) );
  add_747 add_06 ( .s(s[5]), .a(a[5]), .b(n_5_net_), .ci(c[4]), .co(c[5]) );
  add_746 add_07 ( .s(s[6]), .a(a[6]), .b(n_6_net_), .ci(c[5]), .co(c[6]) );
  add_745 add_08 ( .s(s[7]), .a(a[7]), .b(n_7_net_), .ci(c[6]), .co(c[7]) );
  add_744 add_09 ( .s(s[8]), .a(a[8]), .b(n_8_net_), .ci(c[7]), .co(c[8]) );
  add_743 add_10 ( .s(s[9]), .a(a[9]), .b(n_9_net_), .ci(c[8]), .co(c[9]) );
  add_742 add_11 ( .s(s[10]), .a(a[10]), .b(n_10_net_), .ci(c[9]), .co(c[10])
         );
  add_741 add_12 ( .s(s[11]), .a(a[11]), .b(n_11_net_), .ci(c_tmp), .co(c[11])
         );
  add_740 add_13 ( .s(s[12]), .a(a[12]), .b(n_12_net_), .ci(c[11]), .co(c[12])
         );
  add_739 add_14 ( .s(s[13]), .a(a[13]), .b(n_13_net_), .ci(c[12]), .co(c[13])
         );
  add_738 add_15 ( .s(s[14]), .a(a[14]), .b(n_14_net_), .ci(c[13]), .co(c[14])
         );
  add_737 add_16 ( .s(s[15]), .a(a[15]), .b(n_15_net_), .ci(c[14]), .co(c[15])
         );
  add_736 add_17 ( .s(s[16]), .a(a[16]), .b(n_16_net_), .ci(c[15]), .co(c[16])
         );
  add_735 add_18 ( .s(s[17]), .a(a[17]), .b(n_17_net_), .ci(c[16]), .co(c[17])
         );
  add_734 add_19 ( .s(s[18]), .a(a[18]), .b(n_18_net_), .ci(c[17]), .co(c[18])
         );
  add_733 add_20 ( .s(s[19]), .a(a[19]), .b(n_19_net_), .ci(c[18]), .co(c[19])
         );
  add_732 add_21 ( .s(s[20]), .a(a[20]), .b(n_20_net_), .ci(c[19]), .co(c[20])
         );
  add_731 add_22 ( .s(s[21]), .a(a[21]), .b(n_21_net_), .ci(c[20]), .co(c[21])
         );
  add_730 add_23 ( .s(s[22]), .a(a[22]), .b(n_22_net_), .ci(c[21]), .co(c[22])
         );
  add_729 add_24 ( .s(s[23]), .a(a[23]), .b(n_23_net_), .ci(c[22]), .co(c[23])
         );
  DFFARX1 out_reg_10_ ( .D(s[10]), .CLK(clk), .RSTB(rst_n), .Q(out[10]) );
  DFFARX1 out_reg_9_ ( .D(s[9]), .CLK(clk), .RSTB(rst_n), .Q(out[9]) );
  DFFARX1 out_reg_8_ ( .D(s[8]), .CLK(clk), .RSTB(rst_n), .Q(out[8]) );
  DFFARX1 out_reg_7_ ( .D(s[7]), .CLK(clk), .RSTB(rst_n), .Q(out[7]) );
  DFFARX1 out_reg_6_ ( .D(s[6]), .CLK(clk), .RSTB(rst_n), .Q(out[6]) );
  DFFARX1 out_reg_5_ ( .D(s[5]), .CLK(clk), .RSTB(rst_n), .Q(out[5]) );
  DFFARX1 out_reg_4_ ( .D(s[4]), .CLK(clk), .RSTB(rst_n), .Q(out[4]) );
  DFFARX1 out_reg_3_ ( .D(s[3]), .CLK(clk), .RSTB(rst_n), .Q(out[3]) );
  DFFARX1 out_reg_2_ ( .D(s[2]), .CLK(clk), .RSTB(rst_n), .Q(out[2]) );
  DFFARX1 out_reg_1_ ( .D(s[1]), .CLK(clk), .RSTB(rst_n), .Q(out[1]) );
  DFFARX1 out_reg_0_ ( .D(s[0]), .CLK(clk), .RSTB(rst_n), .Q(out[0]) );
  DFFARX1 c_tmp_reg ( .D(c[10]), .CLK(clk), .RSTB(rst_n), .Q(c_tmp) );
  DFFARX1 out_reg_24_ ( .D(s[24]), .CLK(clk), .RSTB(rst_n), .Q(out[24]) );
  DFFARX1 out_reg_23_ ( .D(s[23]), .CLK(clk), .RSTB(rst_n), .Q(out[23]) );
  DFFARX1 out_reg_22_ ( .D(s[22]), .CLK(clk), .RSTB(rst_n), .Q(out[22]) );
  DFFARX1 out_reg_21_ ( .D(s[21]), .CLK(clk), .RSTB(rst_n), .Q(out[21]) );
  DFFARX1 out_reg_20_ ( .D(s[20]), .CLK(clk), .RSTB(rst_n), .Q(out[20]) );
  DFFARX1 out_reg_19_ ( .D(s[19]), .CLK(clk), .RSTB(rst_n), .Q(out[19]) );
  DFFARX1 out_reg_18_ ( .D(s[18]), .CLK(clk), .RSTB(rst_n), .Q(out[18]) );
  DFFARX1 out_reg_17_ ( .D(s[17]), .CLK(clk), .RSTB(rst_n), .Q(out[17]) );
  DFFARX1 out_reg_16_ ( .D(s[16]), .CLK(clk), .RSTB(rst_n), .Q(out[16]) );
  DFFARX1 out_reg_15_ ( .D(s[15]), .CLK(clk), .RSTB(rst_n), .Q(out[15]) );
  DFFARX1 out_reg_14_ ( .D(s[14]), .CLK(clk), .RSTB(rst_n), .Q(out[14]) );
  DFFARX1 out_reg_13_ ( .D(s[13]), .CLK(clk), .RSTB(rst_n), .Q(out[13]) );
  DFFARX1 out_reg_12_ ( .D(s[12]), .CLK(clk), .RSTB(rst_n), .Q(out[12]) );
  DFFARX1 out_reg_11_ ( .D(s[11]), .CLK(clk), .RSTB(rst_n), .Q(out[11]) );
  INVX0 U3 ( .INP(b[1]), .ZN(n_1_net_) );
  INVX0 U4 ( .INP(b[2]), .ZN(n_2_net_) );
  INVX0 U5 ( .INP(b[3]), .ZN(n_3_net_) );
  INVX0 U6 ( .INP(b[4]), .ZN(n_4_net_) );
  INVX0 U7 ( .INP(b[5]), .ZN(n_5_net_) );
  INVX0 U8 ( .INP(b[6]), .ZN(n_6_net_) );
  INVX0 U9 ( .INP(b[7]), .ZN(n_7_net_) );
  INVX0 U10 ( .INP(b[8]), .ZN(n_8_net_) );
  INVX0 U11 ( .INP(b[9]), .ZN(n_9_net_) );
  INVX0 U12 ( .INP(b[10]), .ZN(n_10_net_) );
  INVX0 U13 ( .INP(c[23]), .ZN(s[24]) );
  INVX0 U14 ( .INP(b[11]), .ZN(n_11_net_) );
  INVX0 U15 ( .INP(b[12]), .ZN(n_12_net_) );
  INVX0 U16 ( .INP(b[13]), .ZN(n_13_net_) );
  INVX0 U17 ( .INP(b[14]), .ZN(n_14_net_) );
  INVX0 U18 ( .INP(b[15]), .ZN(n_15_net_) );
  INVX0 U19 ( .INP(b[16]), .ZN(n_16_net_) );
  INVX0 U20 ( .INP(b[17]), .ZN(n_17_net_) );
  INVX0 U21 ( .INP(b[18]), .ZN(n_18_net_) );
  INVX0 U22 ( .INP(b[19]), .ZN(n_19_net_) );
  INVX0 U23 ( .INP(b[20]), .ZN(n_20_net_) );
  INVX0 U24 ( .INP(b[21]), .ZN(n_21_net_) );
  INVX0 U25 ( .INP(b[22]), .ZN(n_22_net_) );
  INVX0 U26 ( .INP(b[23]), .ZN(n_23_net_) );
endmodule


module add_705 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_706 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_707 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_708 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_709 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_710 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_711 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_712 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_713 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_714 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_715 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_716 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_717 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_718 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_719 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_720 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_721 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_722 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_723 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_724 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_725 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_726 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_727 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_728 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(b), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(b), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module adder24_13 ( clk, rst_n, a, b, cin, out );
  input [23:0] a;
  input [23:0] b;
  output [24:0] out;
  input clk, rst_n, cin;
  wire   c_tmp;
  wire   [24:0] s;
  wire   [22:0] c;

  add_728 add_01 ( .s(s[0]), .a(a[0]), .b(b[0]), .ci(1'b0), .co(c[0]) );
  add_727 add_02 ( .s(s[1]), .a(a[1]), .b(b[1]), .ci(c[0]), .co(c[1]) );
  add_726 add_03 ( .s(s[2]), .a(a[2]), .b(b[2]), .ci(c[1]), .co(c[2]) );
  add_725 add_04 ( .s(s[3]), .a(a[3]), .b(b[3]), .ci(c[2]), .co(c[3]) );
  add_724 add_05 ( .s(s[4]), .a(a[4]), .b(b[4]), .ci(c[3]), .co(c[4]) );
  add_723 add_06 ( .s(s[5]), .a(a[5]), .b(b[5]), .ci(c[4]), .co(c[5]) );
  add_722 add_07 ( .s(s[6]), .a(a[6]), .b(b[6]), .ci(c[5]), .co(c[6]) );
  add_721 add_08 ( .s(s[7]), .a(a[7]), .b(b[7]), .ci(c[6]), .co(c[7]) );
  add_720 add_09 ( .s(s[8]), .a(a[8]), .b(b[8]), .ci(c[7]), .co(c[8]) );
  add_719 add_10 ( .s(s[9]), .a(a[9]), .b(b[9]), .ci(c[8]), .co(c[9]) );
  add_718 add_11 ( .s(s[10]), .a(a[10]), .b(b[10]), .ci(c[9]), .co(c[10]) );
  add_717 add_12 ( .s(s[11]), .a(a[11]), .b(b[11]), .ci(c_tmp), .co(c[11]) );
  add_716 add_13 ( .s(s[12]), .a(a[12]), .b(b[12]), .ci(c[11]), .co(c[12]) );
  add_715 add_14 ( .s(s[13]), .a(a[13]), .b(b[13]), .ci(c[12]), .co(c[13]) );
  add_714 add_15 ( .s(s[14]), .a(a[14]), .b(b[14]), .ci(c[13]), .co(c[14]) );
  add_713 add_16 ( .s(s[15]), .a(a[15]), .b(b[15]), .ci(c[14]), .co(c[15]) );
  add_712 add_17 ( .s(s[16]), .a(a[16]), .b(b[16]), .ci(c[15]), .co(c[16]) );
  add_711 add_18 ( .s(s[17]), .a(a[17]), .b(b[17]), .ci(c[16]), .co(c[17]) );
  add_710 add_19 ( .s(s[18]), .a(a[18]), .b(b[18]), .ci(c[17]), .co(c[18]) );
  add_709 add_20 ( .s(s[19]), .a(a[19]), .b(b[19]), .ci(c[18]), .co(c[19]) );
  add_708 add_21 ( .s(s[20]), .a(a[20]), .b(b[20]), .ci(c[19]), .co(c[20]) );
  add_707 add_22 ( .s(s[21]), .a(a[21]), .b(b[21]), .ci(c[20]), .co(c[21]) );
  add_706 add_23 ( .s(s[22]), .a(a[22]), .b(b[22]), .ci(c[21]), .co(c[22]) );
  add_705 add_24 ( .s(s[23]), .a(a[23]), .b(b[23]), .ci(c[22]), .co(s[24]) );
  DFFARX1 out_reg_10_ ( .D(s[10]), .CLK(clk), .RSTB(rst_n), .Q(out[10]) );
  DFFARX1 out_reg_9_ ( .D(s[9]), .CLK(clk), .RSTB(rst_n), .Q(out[9]) );
  DFFARX1 out_reg_8_ ( .D(s[8]), .CLK(clk), .RSTB(rst_n), .Q(out[8]) );
  DFFARX1 out_reg_7_ ( .D(s[7]), .CLK(clk), .RSTB(rst_n), .Q(out[7]) );
  DFFARX1 out_reg_6_ ( .D(s[6]), .CLK(clk), .RSTB(rst_n), .Q(out[6]) );
  DFFARX1 out_reg_5_ ( .D(s[5]), .CLK(clk), .RSTB(rst_n), .Q(out[5]) );
  DFFARX1 out_reg_4_ ( .D(s[4]), .CLK(clk), .RSTB(rst_n), .Q(out[4]) );
  DFFARX1 out_reg_3_ ( .D(s[3]), .CLK(clk), .RSTB(rst_n), .Q(out[3]) );
  DFFARX1 out_reg_2_ ( .D(s[2]), .CLK(clk), .RSTB(rst_n), .Q(out[2]) );
  DFFARX1 out_reg_1_ ( .D(s[1]), .CLK(clk), .RSTB(rst_n), .Q(out[1]) );
  DFFARX1 out_reg_0_ ( .D(s[0]), .CLK(clk), .RSTB(rst_n), .Q(out[0]) );
  DFFARX1 c_tmp_reg ( .D(c[10]), .CLK(clk), .RSTB(rst_n), .Q(c_tmp) );
  DFFARX1 out_reg_24_ ( .D(s[24]), .CLK(clk), .RSTB(rst_n), .Q(out[24]) );
  DFFARX1 out_reg_23_ ( .D(s[23]), .CLK(clk), .RSTB(rst_n), .Q(out[23]) );
  DFFARX1 out_reg_22_ ( .D(s[22]), .CLK(clk), .RSTB(rst_n), .Q(out[22]) );
  DFFARX1 out_reg_21_ ( .D(s[21]), .CLK(clk), .RSTB(rst_n), .Q(out[21]) );
  DFFARX1 out_reg_20_ ( .D(s[20]), .CLK(clk), .RSTB(rst_n), .Q(out[20]) );
  DFFARX1 out_reg_19_ ( .D(s[19]), .CLK(clk), .RSTB(rst_n), .Q(out[19]) );
  DFFARX1 out_reg_18_ ( .D(s[18]), .CLK(clk), .RSTB(rst_n), .Q(out[18]) );
  DFFARX1 out_reg_17_ ( .D(s[17]), .CLK(clk), .RSTB(rst_n), .Q(out[17]) );
  DFFARX1 out_reg_16_ ( .D(s[16]), .CLK(clk), .RSTB(rst_n), .Q(out[16]) );
  DFFARX1 out_reg_15_ ( .D(s[15]), .CLK(clk), .RSTB(rst_n), .Q(out[15]) );
  DFFARX1 out_reg_14_ ( .D(s[14]), .CLK(clk), .RSTB(rst_n), .Q(out[14]) );
  DFFARX1 out_reg_13_ ( .D(s[13]), .CLK(clk), .RSTB(rst_n), .Q(out[13]) );
  DFFARX1 out_reg_12_ ( .D(s[12]), .CLK(clk), .RSTB(rst_n), .Q(out[12]) );
  DFFARX1 out_reg_11_ ( .D(s[11]), .CLK(clk), .RSTB(rst_n), .Q(out[11]) );
endmodule


module add_673 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  XNOR2X1 U1 ( .IN1(ci), .IN2(a), .Q(s) );
endmodule


module add_674 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_675 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_676 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_677 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_678 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_679 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_680 ( s, a, ci, co, b_BAR );
  input a, ci, b_BAR;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(b_BAR), .IN2(n1), .QN(co) );
  INVX0 U2 ( .INP(a), .ZN(n1) );
  MUX21X1 U3 ( .IN1(a), .IN2(n1), .S(b_BAR), .Q(s) );
endmodule


module adder8_49 ( out, a, b, cin );
  output [7:0] out;
  input [7:0] a;
  input [7:0] b;
  input cin;
  wire   n_1_net_, n_2_net_, n_4_net_;
  wire   [6:0] c;

  add_680 add_01 ( .s(out[0]), .a(a[0]), .ci(1'b1), .co(c[0]), .b_BAR(b[0]) );
  add_679 add_02 ( .s(out[1]), .a(a[1]), .b(n_1_net_), .ci(c[0]), .co(c[1]) );
  add_678 add_03 ( .s(out[2]), .a(a[2]), .b(n_2_net_), .ci(c[1]), .co(c[2]) );
  add_677 add_04 ( .s(out[3]), .a(a[3]), .b(1'b1), .ci(c[2]), .co(c[3]) );
  add_676 add_05 ( .s(out[4]), .a(a[4]), .b(n_4_net_), .ci(c[3]), .co(c[4]) );
  add_675 add_06 ( .s(out[5]), .a(a[5]), .b(1'b1), .ci(c[4]), .co(c[5]) );
  add_674 add_07 ( .s(out[6]), .a(a[6]), .b(1'b1), .ci(c[5]), .co(c[6]) );
  add_673 add_08 ( .s(out[7]), .a(a[7]), .b(1'b1), .ci(c[6]) );
  INVX0 U1 ( .INP(b[1]), .ZN(n_1_net_) );
  INVX0 U2 ( .INP(b[2]), .ZN(n_2_net_) );
  INVX0 U3 ( .INP(b[4]), .ZN(n_4_net_) );
endmodule


module add_681 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  XNOR2X1 U1 ( .IN1(ci), .IN2(a), .Q(s) );
endmodule


module add_682 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_683 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_684 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_685 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_686 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_687 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_688 ( s, a, ci, co, b_BAR );
  input a, ci, b_BAR;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(b_BAR), .IN2(n1), .QN(co) );
  INVX0 U2 ( .INP(a), .ZN(n1) );
  MUX21X1 U3 ( .IN1(a), .IN2(n1), .S(b_BAR), .Q(s) );
endmodule


module adder8_50 ( out, a, b, cin );
  output [7:0] out;
  input [7:0] a;
  input [7:0] b;
  input cin;
  wire   n_1_net_, n_2_net_, n_3_net_;
  wire   [6:0] c;

  add_688 add_01 ( .s(out[0]), .a(a[0]), .ci(1'b1), .co(c[0]), .b_BAR(b[0]) );
  add_687 add_02 ( .s(out[1]), .a(a[1]), .b(n_1_net_), .ci(c[0]), .co(c[1]) );
  add_686 add_03 ( .s(out[2]), .a(a[2]), .b(n_2_net_), .ci(c[1]), .co(c[2]) );
  add_685 add_04 ( .s(out[3]), .a(a[3]), .b(n_3_net_), .ci(c[2]), .co(c[3]) );
  add_684 add_05 ( .s(out[4]), .a(a[4]), .b(1'b1), .ci(c[3]), .co(c[4]) );
  add_683 add_06 ( .s(out[5]), .a(a[5]), .b(1'b1), .ci(c[4]), .co(c[5]) );
  add_682 add_07 ( .s(out[6]), .a(a[6]), .b(1'b1), .ci(c[5]), .co(c[6]) );
  add_681 add_08 ( .s(out[7]), .a(a[7]), .b(1'b1), .ci(c[6]) );
  INVX0 U1 ( .INP(b[1]), .ZN(n_1_net_) );
  INVX0 U2 ( .INP(b[2]), .ZN(n_2_net_) );
  INVX0 U3 ( .INP(b[3]), .ZN(n_3_net_) );
endmodule


module add_689 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  XNOR2X1 U1 ( .IN1(ci), .IN2(a), .Q(s) );
endmodule


module add_690 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_691 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_692 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_693 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_694 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_695 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_696 ( s, a, ci, co, b_BAR );
  input a, ci, b_BAR;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(b_BAR), .IN2(n1), .QN(co) );
  INVX0 U2 ( .INP(a), .ZN(n1) );
  MUX21X1 U3 ( .IN1(a), .IN2(n1), .S(b_BAR), .Q(s) );
endmodule


module adder8_51 ( out, a, b, cin );
  output [7:0] out;
  input [7:0] a;
  input [7:0] b;
  input cin;
  wire   n_1_net_, n_2_net_, n_3_net_;
  wire   [6:0] c;

  add_696 add_01 ( .s(out[0]), .a(a[0]), .ci(1'b1), .co(c[0]), .b_BAR(b[0]) );
  add_695 add_02 ( .s(out[1]), .a(a[1]), .b(n_1_net_), .ci(c[0]), .co(c[1]) );
  add_694 add_03 ( .s(out[2]), .a(a[2]), .b(n_2_net_), .ci(c[1]), .co(c[2]) );
  add_693 add_04 ( .s(out[3]), .a(a[3]), .b(n_3_net_), .ci(c[2]), .co(c[3]) );
  add_692 add_05 ( .s(out[4]), .a(a[4]), .b(1'b1), .ci(c[3]), .co(c[4]) );
  add_691 add_06 ( .s(out[5]), .a(a[5]), .b(1'b1), .ci(c[4]), .co(c[5]) );
  add_690 add_07 ( .s(out[6]), .a(a[6]), .b(1'b1), .ci(c[5]), .co(c[6]) );
  add_689 add_08 ( .s(out[7]), .a(a[7]), .b(1'b1), .ci(c[6]) );
  INVX0 U1 ( .INP(b[1]), .ZN(n_1_net_) );
  INVX0 U2 ( .INP(b[2]), .ZN(n_2_net_) );
  INVX0 U3 ( .INP(b[3]), .ZN(n_3_net_) );
endmodule


module add_697 ( s, a, b, co, ci_BAR );
  input a, b, ci_BAR;
  output s, co;


  XNOR2X1 U1 ( .IN1(a), .IN2(ci_BAR), .Q(s) );
endmodule


module add_698 ( s, a, b, ci, co_BAR );
  input a, b, ci;
  output s, co_BAR;


  NAND2X0 U1 ( .IN1(ci), .IN2(a), .QN(co_BAR) );
  OA21X1 U2 ( .IN1(ci), .IN2(a), .IN3(co_BAR), .Q(s) );
endmodule


module add_699 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_700 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_701 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_702 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_703 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_704 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(b), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(b), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module adder8_52 ( out, a, b, cin );
  output [7:0] out;
  input [7:0] a;
  input [7:0] b;
  input cin;

  wire   [6:0] c;

  add_704 add_01 ( .s(out[0]), .a(a[0]), .b(b[0]), .ci(1'b0), .co(c[0]) );
  add_703 add_02 ( .s(out[1]), .a(a[1]), .b(1'b0), .ci(c[0]), .co(c[1]) );
  add_702 add_03 ( .s(out[2]), .a(a[2]), .b(1'b0), .ci(c[1]), .co(c[2]) );
  add_701 add_04 ( .s(out[3]), .a(a[3]), .b(1'b0), .ci(c[2]), .co(c[3]) );
  add_700 add_05 ( .s(out[4]), .a(a[4]), .b(1'b0), .ci(c[3]), .co(c[4]) );
  add_699 add_06 ( .s(out[5]), .a(a[5]), .b(1'b0), .ci(c[4]), .co(c[5]) );
  add_698 add_07 ( .s(out[6]), .a(a[6]), .b(1'b0), .ci(c[5]), .co_BAR(c[6]) );
  add_697 add_08 ( .s(out[7]), .a(a[7]), .b(1'b0), .ci_BAR(c[6]) );
endmodule


module add_753 ( s, a, ci, co, b_BAR );
  input a, ci, b_BAR;
  output s, co;


  XNOR3X1 U1 ( .IN1(b_BAR), .IN2(ci), .IN3(a), .Q(s) );
endmodule


module add_754 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_755 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_756 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_757 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_758 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_759 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_760 ( s, a, ci, co, b_BAR );
  input a, ci, b_BAR;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(b_BAR), .IN2(n1), .QN(co) );
  INVX0 U2 ( .INP(a), .ZN(n1) );
  MUX21X1 U3 ( .IN1(a), .IN2(n1), .S(b_BAR), .Q(s) );
endmodule


module adder8_53 ( out, a, b, cin );
  output [7:0] out;
  input [7:0] a;
  input [7:0] b;
  input cin;
  wire   n_1_net_, n_2_net_, n_3_net_, n_4_net_, n_5_net_, n_6_net_;
  wire   [6:0] c;

  add_760 add_01 ( .s(out[0]), .a(a[0]), .ci(1'b1), .co(c[0]), .b_BAR(b[0]) );
  add_759 add_02 ( .s(out[1]), .a(a[1]), .b(n_1_net_), .ci(c[0]), .co(c[1]) );
  add_758 add_03 ( .s(out[2]), .a(a[2]), .b(n_2_net_), .ci(c[1]), .co(c[2]) );
  add_757 add_04 ( .s(out[3]), .a(a[3]), .b(n_3_net_), .ci(c[2]), .co(c[3]) );
  add_756 add_05 ( .s(out[4]), .a(a[4]), .b(n_4_net_), .ci(c[3]), .co(c[4]) );
  add_755 add_06 ( .s(out[5]), .a(a[5]), .b(n_5_net_), .ci(c[4]), .co(c[5]) );
  add_754 add_07 ( .s(out[6]), .a(a[6]), .b(n_6_net_), .ci(c[5]), .co(c[6]) );
  add_753 add_08 ( .s(out[7]), .a(a[7]), .ci(c[6]), .b_BAR(b[7]) );
  INVX0 U1 ( .INP(b[1]), .ZN(n_1_net_) );
  INVX0 U2 ( .INP(b[2]), .ZN(n_2_net_) );
  INVX0 U3 ( .INP(b[3]), .ZN(n_3_net_) );
  INVX0 U4 ( .INP(b[4]), .ZN(n_4_net_) );
  INVX0 U5 ( .INP(b[5]), .ZN(n_5_net_) );
  INVX0 U6 ( .INP(b[6]), .ZN(n_6_net_) );
endmodule


module add_761 ( s, a, ci, co, b_BAR );
  input a, ci, b_BAR;
  output s, co;


  XNOR3X1 U1 ( .IN1(b_BAR), .IN2(ci), .IN3(a), .Q(s) );
endmodule


module add_762 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_763 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_764 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_765 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_766 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_767 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_768 ( s, a, ci, co, b_BAR );
  input a, ci, b_BAR;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(b_BAR), .IN2(n1), .QN(co) );
  INVX0 U2 ( .INP(a), .ZN(n1) );
  MUX21X1 U3 ( .IN1(a), .IN2(n1), .S(b_BAR), .Q(s) );
endmodule


module adder8_54 ( out, a, b, cin );
  output [7:0] out;
  input [7:0] a;
  input [7:0] b;
  input cin;
  wire   n_1_net_, n_2_net_, n_3_net_, n_4_net_, n_5_net_, n_6_net_;
  wire   [6:0] c;

  add_768 add_01 ( .s(out[0]), .a(a[0]), .ci(1'b1), .co(c[0]), .b_BAR(b[0]) );
  add_767 add_02 ( .s(out[1]), .a(a[1]), .b(n_1_net_), .ci(c[0]), .co(c[1]) );
  add_766 add_03 ( .s(out[2]), .a(a[2]), .b(n_2_net_), .ci(c[1]), .co(c[2]) );
  add_765 add_04 ( .s(out[3]), .a(a[3]), .b(n_3_net_), .ci(c[2]), .co(c[3]) );
  add_764 add_05 ( .s(out[4]), .a(a[4]), .b(n_4_net_), .ci(c[3]), .co(c[4]) );
  add_763 add_06 ( .s(out[5]), .a(a[5]), .b(n_5_net_), .ci(c[4]), .co(c[5]) );
  add_762 add_07 ( .s(out[6]), .a(a[6]), .b(n_6_net_), .ci(c[5]), .co(c[6]) );
  add_761 add_08 ( .s(out[7]), .a(a[7]), .ci(c[6]), .b_BAR(b[7]) );
  INVX0 U1 ( .INP(b[1]), .ZN(n_1_net_) );
  INVX0 U2 ( .INP(b[2]), .ZN(n_2_net_) );
  INVX0 U3 ( .INP(b[3]), .ZN(n_3_net_) );
  INVX0 U4 ( .INP(b[4]), .ZN(n_4_net_) );
  INVX0 U5 ( .INP(b[5]), .ZN(n_5_net_) );
  INVX0 U6 ( .INP(b[6]), .ZN(n_6_net_) );
endmodule


module floating_point_adder_0 ( clk, rst_n, input_factor_01, input_factor_02, 
        output_adder );
  input [31:0] input_factor_01;
  input [31:0] input_factor_02;
  output [31:0] output_adder;
  input clk, rst_n;
  wire   N34, N35, N36, N37, N38, N39, N40, N41, N152, N153, N154, N155, N156,
         N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, N167,
         N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178,
         N179, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189,
         N190, N191, N192, N193, N194, N195, N196, N197, N198,
         add_sub_result_24_, N211, shift_temp_01_0_, N226, N227, N228, N229,
         N230, N231, N232, N233, N234, N235, N236, N237, N238, N239, N240,
         N241, N242, N243, N244, N245, N246, N247, N248, N256, N257, N258,
         N260, N261, N262, N263, N264, N265, N266, N267, N268, N269, N270,
         N271, N272, N273, N274, N275, N276, N277, N278, N279, N280, N281,
         N306, N307, N308, N346, N347, N348, N349, N350, N351, N352, N353,
         N354, N355, N380, N381, N382, N383, N384, N385, N386, N387, N388,
         N389, N390, N391, N392, N393, N394, N395, N396, N397, N398, N399,
         N400, N401, N402, N403, N404, N405, N406, N407, N408, N409, N410, n78,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n138, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850;
  wire   [7:0] exp_diff_value;
  wire   [7:0] exponent_factor_21;
  wire   [7:0] exponent_factor_12;
  wire   [23:0] shift_smaller_factor;
  wire   [22:0] larger_factor;
  wire   [7:0] larger_exponent;
  wire   [24:0] add_result;
  wire   [24:0] sub_result;
  wire   [22:0] pre_sig_res_01;
  wire   [3:0] shift_temp_02;
  wire   [22:1] pre_sig_res_02;
  wire   [2:0] shift_temp_03;
  wire   [22:9] pre_sig_res_03;
  wire   [4:0] shift_temp_04;
  wire   [22:16] pre_sig_res_04;
  wire   [7:0] add_output_exponent_w1;
  wire   [7:0] add_output_exponent_w2;
  wire   [7:0] add_output_exponent_w3;
  wire   [7:0] add_output_exponent_w4;

  adder8_54 adder8_01 ( .out(exponent_factor_21), .a(input_factor_02[30:23]), 
        .b(input_factor_01[30:23]), .cin(1'b1) );
  adder8_53 adder8_02 ( .out(exponent_factor_12), .a(input_factor_01[30:23]), 
        .b(input_factor_02[30:23]), .cin(1'b1) );
  adder24_0 adder24_01 ( .clk(clk), .rst_n(rst_n), .a({shift_temp_04[4], 
        larger_factor}), .b(shift_smaller_factor), .cin(1'b1), .out(sub_result) );
  adder24_13 adder24_02 ( .clk(clk), .rst_n(rst_n), .a({shift_temp_04[4], 
        larger_factor}), .b(shift_smaller_factor), .cin(1'b0), .out(add_result) );
  adder8_52 adder8_03 ( .out(add_output_exponent_w1), .a(larger_exponent), .b(
        {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, shift_temp_01_0_}), .cin(
        1'b0) );
  adder8_51 adder8_04 ( .out(add_output_exponent_w2), .a(larger_exponent), .b(
        {1'b0, 1'b0, 1'b0, 1'b0, shift_temp_02}), .cin(1'b1) );
  adder8_50 adder8_05 ( .out(add_output_exponent_w3), .a(larger_exponent), .b(
        {1'b0, 1'b0, 1'b0, 1'b0, shift_temp_04[4], shift_temp_03}), .cin(1'b1)
         );
  adder8_49 adder8_06 ( .out(add_output_exponent_w4), .a(larger_exponent), .b(
        {1'b0, 1'b0, 1'b0, shift_temp_04[4], 1'b0, shift_temp_04[2:0]}), .cin(
        1'b1) );
  DFFARX1 exp_diff_value_reg_7_ ( .D(N41), .CLK(clk), .RSTB(rst_n), .Q(
        exp_diff_value[7]) );
  DFFARX1 exp_diff_value_reg_6_ ( .D(N40), .CLK(clk), .RSTB(rst_n), .Q(
        exp_diff_value[6]) );
  DFFARX1 exp_diff_value_reg_5_ ( .D(N39), .CLK(clk), .RSTB(rst_n), .Q(
        exp_diff_value[5]) );
  DFFARX1 exp_diff_value_reg_4_ ( .D(N38), .CLK(clk), .RSTB(rst_n), .Q(
        exp_diff_value[4]) );
  DFFARX1 exp_diff_value_reg_3_ ( .D(N37), .CLK(clk), .RSTB(rst_n), .Q(
        exp_diff_value[3]), .QN(n4) );
  DFFARX1 exp_diff_value_reg_2_ ( .D(N36), .CLK(clk), .RSTB(rst_n), .Q(
        exp_diff_value[2]), .QN(n2) );
  DFFARX1 exp_diff_value_reg_1_ ( .D(N35), .CLK(clk), .RSTB(rst_n), .Q(
        exp_diff_value[1]), .QN(n3) );
  DFFARX1 exp_diff_value_reg_0_ ( .D(N34), .CLK(clk), .RSTB(rst_n), .Q(
        exp_diff_value[0]), .QN(n1) );
  DFFARX1 larger_factor_reg_22_ ( .D(N198), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[22]) );
  DFFARX1 larger_factor_reg_21_ ( .D(N197), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[21]) );
  DFFARX1 larger_factor_reg_20_ ( .D(N196), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[20]) );
  DFFARX1 larger_factor_reg_19_ ( .D(N195), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[19]) );
  DFFARX1 larger_factor_reg_18_ ( .D(N194), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[18]) );
  DFFARX1 larger_factor_reg_17_ ( .D(N193), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[17]) );
  DFFARX1 larger_factor_reg_16_ ( .D(N192), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[16]) );
  DFFARX1 larger_factor_reg_15_ ( .D(N191), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[15]) );
  DFFARX1 larger_factor_reg_14_ ( .D(N190), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[14]) );
  DFFARX1 larger_factor_reg_13_ ( .D(N189), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[13]) );
  DFFARX1 larger_factor_reg_12_ ( .D(N188), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[12]) );
  DFFARX1 larger_factor_reg_11_ ( .D(N187), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[11]) );
  DFFARX1 larger_factor_reg_10_ ( .D(N186), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[10]) );
  DFFARX1 larger_factor_reg_9_ ( .D(N185), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[9]) );
  DFFARX1 larger_factor_reg_8_ ( .D(N184), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[8]) );
  DFFARX1 larger_factor_reg_7_ ( .D(N183), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[7]) );
  DFFARX1 larger_factor_reg_6_ ( .D(N182), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[6]) );
  DFFARX1 larger_factor_reg_5_ ( .D(N181), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[5]) );
  DFFARX1 larger_factor_reg_4_ ( .D(N180), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[4]) );
  DFFARX1 larger_factor_reg_3_ ( .D(N179), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[3]) );
  DFFARX1 larger_factor_reg_2_ ( .D(N178), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[2]) );
  DFFARX1 larger_factor_reg_1_ ( .D(N177), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[1]) );
  DFFARX1 larger_factor_reg_0_ ( .D(N176), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[0]) );
  DFFARX1 shift_smaller_factor_reg_23_ ( .D(N175), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[23]) );
  DFFARX1 shift_smaller_factor_reg_22_ ( .D(N174), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[22]) );
  DFFARX1 shift_smaller_factor_reg_21_ ( .D(N173), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[21]) );
  DFFARX1 shift_smaller_factor_reg_20_ ( .D(N172), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[20]) );
  DFFARX1 shift_smaller_factor_reg_19_ ( .D(N171), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[19]) );
  DFFARX1 shift_smaller_factor_reg_18_ ( .D(N170), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[18]) );
  DFFARX1 shift_smaller_factor_reg_17_ ( .D(N169), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[17]) );
  DFFARX1 shift_smaller_factor_reg_16_ ( .D(N168), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[16]) );
  DFFARX1 shift_smaller_factor_reg_15_ ( .D(N167), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[15]) );
  DFFARX1 shift_smaller_factor_reg_14_ ( .D(N166), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[14]) );
  DFFARX1 shift_smaller_factor_reg_13_ ( .D(N165), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[13]) );
  DFFARX1 shift_smaller_factor_reg_12_ ( .D(N164), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[12]) );
  DFFARX1 shift_smaller_factor_reg_11_ ( .D(N163), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[11]) );
  DFFARX1 shift_smaller_factor_reg_10_ ( .D(N162), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[10]) );
  DFFARX1 shift_smaller_factor_reg_9_ ( .D(N161), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[9]) );
  DFFARX1 shift_smaller_factor_reg_8_ ( .D(N160), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[8]) );
  DFFARX1 shift_smaller_factor_reg_7_ ( .D(N159), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[7]) );
  DFFARX1 shift_smaller_factor_reg_6_ ( .D(N158), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[6]) );
  DFFARX1 shift_smaller_factor_reg_5_ ( .D(N157), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[5]) );
  DFFARX1 shift_smaller_factor_reg_4_ ( .D(N156), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[4]) );
  DFFARX1 shift_smaller_factor_reg_3_ ( .D(N155), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[3]) );
  DFFARX1 shift_smaller_factor_reg_2_ ( .D(N154), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[2]) );
  DFFARX1 shift_smaller_factor_reg_1_ ( .D(N153), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[1]) );
  DFFARX1 shift_smaller_factor_reg_0_ ( .D(N152), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[0]) );
  DFFX1 larger_exponent_reg_7_ ( .D(n115), .CLK(clk), .Q(larger_exponent[7])
         );
  DFFX1 larger_exponent_reg_6_ ( .D(n114), .CLK(clk), .Q(larger_exponent[6])
         );
  DFFX1 larger_exponent_reg_5_ ( .D(n113), .CLK(clk), .Q(larger_exponent[5])
         );
  DFFX1 larger_exponent_reg_4_ ( .D(n112), .CLK(clk), .Q(larger_exponent[4])
         );
  DFFX1 larger_exponent_reg_3_ ( .D(n111), .CLK(clk), .Q(larger_exponent[3])
         );
  DFFX1 larger_exponent_reg_2_ ( .D(n110), .CLK(clk), .Q(larger_exponent[2])
         );
  DFFX1 larger_exponent_reg_1_ ( .D(n109), .CLK(clk), .Q(larger_exponent[1])
         );
  DFFX1 larger_exponent_reg_0_ ( .D(n108), .CLK(clk), .Q(larger_exponent[0])
         );
  DFFARX1 shift_temp_04_reg_4_ ( .D(1'b1), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_04[4]) );
  DFFARX1 shift_temp_01_reg_0_ ( .D(add_sub_result_24_), .CLK(clk), .RSTB(
        rst_n), .Q(shift_temp_01_0_) );
  DFFARX1 pre_sig_res_02_reg_1_ ( .D(N260), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[1]) );
  DFFARX1 pre_sig_res_02_reg_2_ ( .D(N261), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[2]) );
  DFFARX1 pre_sig_res_02_reg_3_ ( .D(N262), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[3]) );
  DFFARX1 pre_sig_res_02_reg_4_ ( .D(N263), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[4]) );
  DFFARX1 pre_sig_res_02_reg_5_ ( .D(N264), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[5]) );
  DFFARX1 pre_sig_res_02_reg_6_ ( .D(N265), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[6]) );
  DFFARX1 pre_sig_res_02_reg_7_ ( .D(N266), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[7]) );
  DFFARX1 shift_temp_02_reg_2_ ( .D(N258), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_02[2]) );
  DFFASX1 shift_temp_02_reg_3_ ( .D(n138), .CLK(clk), .SETB(rst_n), .QN(
        shift_temp_02[3]) );
  DFFARX1 pre_sig_res_02_reg_8_ ( .D(N267), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[8]) );
  DFFARX1 pre_sig_res_02_reg_9_ ( .D(N268), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[9]) );
  DFFARX1 pre_sig_res_02_reg_10_ ( .D(N269), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[10]) );
  DFFARX1 pre_sig_res_02_reg_11_ ( .D(N270), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[11]) );
  DFFARX1 pre_sig_res_02_reg_12_ ( .D(N271), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[12]) );
  DFFARX1 pre_sig_res_02_reg_13_ ( .D(N272), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[13]) );
  DFFARX1 pre_sig_res_02_reg_14_ ( .D(N273), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[14]) );
  DFFARX1 pre_sig_res_02_reg_15_ ( .D(N274), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[15]) );
  DFFARX1 pre_sig_res_02_reg_16_ ( .D(N275), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[16]) );
  DFFARX1 pre_sig_res_02_reg_17_ ( .D(N276), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[17]) );
  DFFARX1 pre_sig_res_02_reg_18_ ( .D(N277), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[18]) );
  DFFARX1 pre_sig_res_02_reg_19_ ( .D(N278), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[19]) );
  DFFARX1 pre_sig_res_02_reg_20_ ( .D(N279), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[20]) );
  DFFARX1 pre_sig_res_02_reg_21_ ( .D(N280), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[21]) );
  DFFARX1 pre_sig_res_02_reg_22_ ( .D(N281), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[22]) );
  DFFARX1 shift_temp_02_reg_1_ ( .D(N257), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_02[1]) );
  DFFARX1 shift_temp_02_reg_0_ ( .D(N256), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_02[0]) );
  DFFX1 pre_sig_res_03_reg_9_ ( .D(n107), .CLK(clk), .Q(pre_sig_res_03[9]) );
  DFFX1 pre_sig_res_03_reg_10_ ( .D(n106), .CLK(clk), .Q(pre_sig_res_03[10])
         );
  DFFX1 pre_sig_res_03_reg_12_ ( .D(n105), .CLK(clk), .Q(pre_sig_res_03[12])
         );
  DFFX1 pre_sig_res_03_reg_11_ ( .D(n104), .CLK(clk), .Q(pre_sig_res_03[11])
         );
  DFFX1 pre_sig_res_03_reg_13_ ( .D(n103), .CLK(clk), .Q(pre_sig_res_03[13])
         );
  DFFX1 pre_sig_res_03_reg_14_ ( .D(n102), .CLK(clk), .Q(pre_sig_res_03[14])
         );
  DFFARX1 shift_temp_03_reg_2_ ( .D(N308), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_03[2]) );
  DFFARX1 shift_temp_03_reg_0_ ( .D(N306), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_03[0]) );
  DFFARX1 shift_temp_03_reg_1_ ( .D(N307), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_03[1]) );
  DFFX1 pre_sig_res_03_reg_15_ ( .D(n101), .CLK(clk), .Q(pre_sig_res_03[15])
         );
  DFFX1 pre_sig_res_03_reg_16_ ( .D(n100), .CLK(clk), .Q(pre_sig_res_03[16])
         );
  DFFX1 pre_sig_res_03_reg_17_ ( .D(n99), .CLK(clk), .Q(pre_sig_res_03[17]) );
  DFFX1 pre_sig_res_03_reg_18_ ( .D(n98), .CLK(clk), .Q(pre_sig_res_03[18]) );
  DFFX1 pre_sig_res_03_reg_19_ ( .D(n97), .CLK(clk), .Q(pre_sig_res_03[19]) );
  DFFX1 pre_sig_res_03_reg_20_ ( .D(n96), .CLK(clk), .Q(pre_sig_res_03[20]) );
  DFFX1 pre_sig_res_03_reg_21_ ( .D(n95), .CLK(clk), .Q(pre_sig_res_03[21]) );
  DFFX1 pre_sig_res_03_reg_22_ ( .D(n94), .CLK(clk), .Q(pre_sig_res_03[22]) );
  DFFARX1 pre_sig_res_04_reg_16_ ( .D(N349), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_04[16]) );
  DFFARX1 pre_sig_res_04_reg_17_ ( .D(N350), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_04[17]) );
  DFFARX1 pre_sig_res_04_reg_18_ ( .D(N351), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_04[18]) );
  DFFARX1 pre_sig_res_04_reg_19_ ( .D(N352), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_04[19]) );
  DFFARX1 pre_sig_res_04_reg_20_ ( .D(N353), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_04[20]) );
  DFFARX1 pre_sig_res_04_reg_21_ ( .D(N354), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_04[21]) );
  DFFARX1 pre_sig_res_04_reg_22_ ( .D(N355), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_04[22]) );
  DFFARX1 add_output_sign_reg ( .D(N211), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[31]) );
  DFFARX1 pre_sig_res_01_reg_0_ ( .D(N226), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[0]) );
  DFFARX1 pre_sig_res_01_reg_1_ ( .D(N227), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[1]) );
  DFFARX1 pre_sig_res_01_reg_2_ ( .D(N228), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[2]) );
  DFFARX1 pre_sig_res_01_reg_3_ ( .D(N229), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[3]) );
  DFFARX1 pre_sig_res_01_reg_4_ ( .D(N230), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[4]) );
  DFFARX1 pre_sig_res_01_reg_5_ ( .D(N231), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[5]) );
  DFFARX1 pre_sig_res_01_reg_6_ ( .D(N232), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[6]) );
  DFFARX1 pre_sig_res_01_reg_7_ ( .D(N233), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[7]) );
  DFFARX1 pre_sig_res_01_reg_8_ ( .D(N234), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[8]) );
  DFFARX1 pre_sig_res_01_reg_9_ ( .D(N235), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[9]) );
  DFFARX1 pre_sig_res_01_reg_10_ ( .D(N236), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[10]) );
  DFFARX1 pre_sig_res_01_reg_11_ ( .D(N237), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[11]) );
  DFFARX1 pre_sig_res_01_reg_12_ ( .D(N238), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[12]) );
  DFFARX1 pre_sig_res_01_reg_13_ ( .D(N239), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[13]) );
  DFFARX1 pre_sig_res_01_reg_14_ ( .D(N240), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[14]) );
  DFFARX1 pre_sig_res_01_reg_15_ ( .D(N241), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[15]) );
  DFFARX1 pre_sig_res_01_reg_16_ ( .D(N242), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[16]) );
  DFFARX1 pre_sig_res_01_reg_17_ ( .D(N243), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[17]) );
  DFFARX1 pre_sig_res_01_reg_18_ ( .D(N244), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[18]) );
  DFFARX1 pre_sig_res_01_reg_19_ ( .D(N245), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[19]) );
  DFFARX1 pre_sig_res_01_reg_20_ ( .D(N246), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[20]) );
  DFFARX1 pre_sig_res_01_reg_21_ ( .D(N247), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[21]) );
  DFFARX1 pre_sig_res_01_reg_22_ ( .D(N248), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[22]) );
  DFFARX1 shift_temp_04_reg_2_ ( .D(N348), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_04[2]) );
  DFFARX1 shift_temp_04_reg_1_ ( .D(N347), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_04[1]) );
  DFFARX1 shift_temp_04_reg_0_ ( .D(N346), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_04[0]) );
  DFFARX1 add_output_exponent_reg_7_ ( .D(N387), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[30]) );
  DFFARX1 add_output_exponent_reg_6_ ( .D(N386), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[29]) );
  DFFARX1 add_output_exponent_reg_5_ ( .D(N385), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[28]) );
  DFFARX1 add_output_exponent_reg_4_ ( .D(N384), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[27]) );
  DFFARX1 add_output_exponent_reg_3_ ( .D(N383), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[26]) );
  DFFARX1 add_output_exponent_reg_2_ ( .D(N382), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[25]) );
  DFFARX1 add_output_exponent_reg_1_ ( .D(N381), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[24]) );
  DFFARX1 add_output_exponent_reg_0_ ( .D(N380), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[23]) );
  DFFARX1 add_output_significands_reg_22_ ( .D(N410), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[22]) );
  DFFARX1 add_output_significands_reg_21_ ( .D(N409), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[21]) );
  DFFARX1 add_output_significands_reg_20_ ( .D(N408), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[20]) );
  DFFARX1 add_output_significands_reg_19_ ( .D(N407), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[19]) );
  DFFARX1 add_output_significands_reg_18_ ( .D(N406), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[18]) );
  DFFARX1 add_output_significands_reg_17_ ( .D(N405), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[17]) );
  DFFARX1 add_output_significands_reg_16_ ( .D(N404), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[16]) );
  DFFARX1 add_output_significands_reg_15_ ( .D(N403), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[15]) );
  DFFARX1 add_output_significands_reg_14_ ( .D(N402), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[14]) );
  DFFARX1 add_output_significands_reg_13_ ( .D(N401), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[13]) );
  DFFARX1 add_output_significands_reg_12_ ( .D(N400), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[12]) );
  DFFARX1 add_output_significands_reg_11_ ( .D(N399), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[11]) );
  DFFARX1 add_output_significands_reg_10_ ( .D(N398), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[10]) );
  DFFARX1 add_output_significands_reg_9_ ( .D(N397), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[9]) );
  DFFARX1 add_output_significands_reg_8_ ( .D(N396), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[8]) );
  DFFARX1 add_output_significands_reg_7_ ( .D(N395), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[7]) );
  DFFARX1 add_output_significands_reg_6_ ( .D(N394), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[6]) );
  DFFARX1 add_output_significands_reg_5_ ( .D(N393), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[5]) );
  DFFARX1 add_output_significands_reg_4_ ( .D(N392), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[4]) );
  DFFARX1 add_output_significands_reg_3_ ( .D(N391), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[3]) );
  DFFARX1 add_output_significands_reg_2_ ( .D(N390), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[2]) );
  DFFARX1 add_output_significands_reg_1_ ( .D(N389), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[1]) );
  DFFARX1 add_output_significands_reg_0_ ( .D(N388), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[0]) );
  INVX1 U5 ( .INP(rst_n), .ZN(n78) );
  NAND2X0 U3 ( .IN1(n507), .IN2(n420), .QN(n589) );
  NAND2X0 U4 ( .IN1(n287), .IN2(n848), .QN(n266) );
  NAND2X0 U6 ( .IN1(input_factor_02[16]), .IN2(n391), .QN(n52) );
  NAND2X0 U7 ( .IN1(input_factor_02[25]), .IN2(n566), .QN(n55) );
  NAND2X0 U8 ( .IN1(n571), .IN2(input_factor_02[24]), .QN(n56) );
  NAND2X0 U9 ( .IN1(input_factor_02[26]), .IN2(n569), .QN(n62) );
  NAND2X0 U10 ( .IN1(n570), .IN2(input_factor_02[28]), .QN(n63) );
  NAND2X0 U11 ( .IN1(input_factor_02[27]), .IN2(n568), .QN(n65) );
  NAND2X0 U12 ( .IN1(input_factor_02[29]), .IN2(n567), .QN(n70) );
  NAND2X0 U13 ( .IN1(n832), .IN2(n547), .QN(n404) );
  NAND2X0 U14 ( .IN1(n802), .IN2(n539), .QN(n403) );
  NAND2X0 U15 ( .IN1(n795), .IN2(n540), .QN(n402) );
  NAND2X0 U16 ( .IN1(n771), .IN2(n745), .QN(n586) );
  NAND2X0 U17 ( .IN1(n424), .IN2(n517), .QN(n400) );
  NAND2X0 U18 ( .IN1(n515), .IN2(n427), .QN(n399) );
  NAND2X0 U19 ( .IN1(n398), .IN2(n595), .QN(n426) );
  NAND2X0 U20 ( .IN1(n118), .IN2(n117), .QN(n233) );
  NAND2X0 U21 ( .IN1(n150), .IN2(n149), .QN(n250) );
  NAND2X0 U22 ( .IN1(n179), .IN2(n178), .QN(n268) );
  NAND2X0 U23 ( .IN1(n215), .IN2(n214), .QN(n288) );
  NAND2X0 U24 ( .IN1(n116), .IN2(n93), .QN(n224) );
  NAND2X0 U25 ( .IN1(n375), .IN2(n233), .QN(n234) );
  NAND2X0 U26 ( .IN1(n148), .IN2(n147), .QN(n244) );
  NAND2X0 U27 ( .IN1(n375), .IN2(n250), .QN(n251) );
  NAND2X0 U28 ( .IN1(n177), .IN2(n176), .QN(n261) );
  NAND2X0 U29 ( .IN1(n375), .IN2(n268), .QN(n269) );
  NAND2X0 U30 ( .IN1(n726), .IN2(n287), .QN(n270) );
  NAND2X0 U31 ( .IN1(exp_diff_value[0]), .IN2(n3), .QN(n213) );
  NAND2X0 U32 ( .IN1(exp_diff_value[1]), .IN2(exp_diff_value[0]), .QN(n212) );
  NAND2X0 U33 ( .IN1(exp_diff_value[1]), .IN2(n1), .QN(n211) );
  NAND2X0 U34 ( .IN1(n210), .IN2(n209), .QN(n280) );
  NAND2X0 U35 ( .IN1(n375), .IN2(n288), .QN(n289) );
  NAND2X0 U36 ( .IN1(n52), .IN2(n53), .QN(n14) );
  NAND2X0 U37 ( .IN1(n4), .IN2(n2), .QN(n294) );
  NAND2X0 U38 ( .IN1(n394), .IN2(n74), .QN(n397) );
  NAND2X0 U39 ( .IN1(n734), .IN2(pre_sig_res_01[9]), .QN(n652) );
  NAND2X0 U40 ( .IN1(n734), .IN2(pre_sig_res_01[10]), .QN(n658) );
  NAND2X0 U41 ( .IN1(n734), .IN2(pre_sig_res_01[11]), .QN(n664) );
  NAND2X0 U42 ( .IN1(n734), .IN2(pre_sig_res_01[12]), .QN(n670) );
  NAND2X0 U43 ( .IN1(n734), .IN2(pre_sig_res_01[13]), .QN(n676) );
  NAND2X0 U44 ( .IN1(n734), .IN2(pre_sig_res_01[14]), .QN(n682) );
  NAND2X0 U45 ( .IN1(n734), .IN2(pre_sig_res_01[15]), .QN(n688) );
  NAND2X0 U46 ( .IN1(n734), .IN2(pre_sig_res_01[16]), .QN(n692) );
  NAND2X0 U47 ( .IN1(n734), .IN2(pre_sig_res_01[17]), .QN(n698) );
  NAND2X0 U48 ( .IN1(n734), .IN2(pre_sig_res_01[18]), .QN(n704) );
  NAND2X0 U49 ( .IN1(n734), .IN2(pre_sig_res_01[19]), .QN(n710) );
  NAND2X0 U50 ( .IN1(n734), .IN2(pre_sig_res_01[20]), .QN(n716) );
  NAND2X0 U51 ( .IN1(n734), .IN2(pre_sig_res_01[21]), .QN(n722) );
  NAND2X0 U52 ( .IN1(n734), .IN2(pre_sig_res_01[22]), .QN(n735) );
  NAND2X0 U53 ( .IN1(n734), .IN2(add_output_exponent_w1[0]), .QN(n596) );
  NAND2X0 U54 ( .IN1(n734), .IN2(add_output_exponent_w1[1]), .QN(n600) );
  NAND2X0 U55 ( .IN1(n734), .IN2(add_output_exponent_w1[2]), .QN(n604) );
  NAND2X0 U56 ( .IN1(n734), .IN2(add_output_exponent_w1[3]), .QN(n608) );
  NAND2X0 U57 ( .IN1(n734), .IN2(add_output_exponent_w1[4]), .QN(n612) );
  NAND2X0 U58 ( .IN1(n734), .IN2(add_output_exponent_w1[5]), .QN(n616) );
  NAND2X0 U59 ( .IN1(n734), .IN2(add_output_exponent_w1[6]), .QN(n620) );
  NAND2X0 U60 ( .IN1(n734), .IN2(add_output_exponent_w1[7]), .QN(n624) );
  NAND2X0 U61 ( .IN1(n541), .IN2(n842), .QN(n559) );
  NAND2X0 U62 ( .IN1(n538), .IN2(n547), .QN(n544) );
  NAND2X0 U63 ( .IN1(n397), .IN2(n396), .QN(n416) );
  NAND2X0 U64 ( .IN1(n539), .IN2(n815), .QN(n557) );
  NAND2X0 U65 ( .IN1(n540), .IN2(n782), .QN(n558) );
  NAND2X0 U66 ( .IN1(n787), .IN2(n771), .QN(n746) );
  NAND2X0 U67 ( .IN1(n745), .IN2(n758), .QN(n820) );
  NAND2X0 U68 ( .IN1(n537), .IN2(n525), .QN(n749) );
  NAND2X0 U69 ( .IN1(n537), .IN2(n529), .QN(n742) );
  NAND2X0 U70 ( .IN1(n420), .IN2(n419), .QN(n519) );
  NAND2X0 U71 ( .IN1(n437), .IN2(n844), .QN(n434) );
  NAND2X0 U72 ( .IN1(n424), .IN2(n421), .QN(n508) );
  NAND2X0 U73 ( .IN1(n427), .IN2(n422), .QN(n512) );
  NAND2X0 U74 ( .IN1(n423), .IN2(n595), .QN(n510) );
  NAND2X0 U75 ( .IN1(n90), .IN2(n89), .QN(n119) );
  NAND2X0 U76 ( .IN1(n144), .IN2(n143), .QN(n151) );
  NAND2X0 U77 ( .IN1(n173), .IN2(n172), .QN(n180) );
  NAND2X0 U78 ( .IN1(n287), .IN2(n4), .QN(n190) );
  NAND2X0 U79 ( .IN1(n848), .IN2(n393), .QN(n290) );
  NAND2X0 U80 ( .IN1(n726), .IN2(n393), .QN(n232) );
  NAND2X0 U81 ( .IN1(n206), .IN2(n205), .QN(n216) );
  NAND2X0 U82 ( .IN1(n92), .IN2(n91), .QN(n226) );
  NAND2X0 U83 ( .IN1(n234), .IN2(n235), .QN(n12) );
  NAND2X0 U84 ( .IN1(n146), .IN2(n145), .QN(n245) );
  NAND2X0 U85 ( .IN1(n251), .IN2(n252), .QN(n10) );
  NAND2X0 U86 ( .IN1(n175), .IN2(n174), .QN(n262) );
  NAND2X0 U87 ( .IN1(n269), .IN2(n271), .QN(n8) );
  NAND2X0 U88 ( .IN1(n373), .IN2(n227), .QN(n285) );
  NAND2X0 U89 ( .IN1(n208), .IN2(n207), .QN(n281) );
  NAND2X0 U90 ( .IN1(n289), .IN2(n292), .QN(n6) );
  NAND2X0 U91 ( .IN1(exp_diff_value[3]), .IN2(n373), .QN(n349) );
  NAND2X0 U92 ( .IN1(n328), .IN2(n2), .QN(n342) );
  NAND2X0 U93 ( .IN1(n350), .IN2(n349), .QN(n351) );
  NAND2X0 U94 ( .IN1(n373), .IN2(n4), .QN(n367) );
  NAND2X0 U95 ( .IN1(n375), .IN2(n4), .QN(n369) );
  NAND2X0 U96 ( .IN1(n384), .IN2(n76), .QN(n396) );
  NAND2X0 U97 ( .IN1(n392), .IN2(n375), .QN(n387) );
  NAND2X0 U98 ( .IN1(n373), .IN2(n392), .QN(n385) );
  NAND2X0 U99 ( .IN1(n629), .IN2(n628), .QN(N389) );
  NAND2X0 U100 ( .IN1(n631), .IN2(n630), .QN(N390) );
  NAND2X0 U101 ( .IN1(n633), .IN2(n632), .QN(N391) );
  NAND2X0 U102 ( .IN1(n635), .IN2(n634), .QN(N392) );
  NAND2X0 U103 ( .IN1(n637), .IN2(n636), .QN(N393) );
  NAND2X0 U104 ( .IN1(n639), .IN2(n638), .QN(N394) );
  NAND2X0 U105 ( .IN1(n643), .IN2(n642), .QN(N395) );
  NAND2X0 U106 ( .IN1(n647), .IN2(n646), .QN(N396) );
  NAND2X0 U107 ( .IN1(n732), .IN2(pre_sig_res_03[9]), .QN(n650) );
  NAND2X0 U108 ( .IN1(n731), .IN2(pre_sig_res_02[9]), .QN(n651) );
  NAND2X0 U109 ( .IN1(n732), .IN2(pre_sig_res_03[10]), .QN(n656) );
  NAND2X0 U110 ( .IN1(n731), .IN2(pre_sig_res_02[10]), .QN(n657) );
  NAND2X0 U111 ( .IN1(n732), .IN2(pre_sig_res_03[11]), .QN(n662) );
  NAND2X0 U112 ( .IN1(n731), .IN2(pre_sig_res_02[11]), .QN(n663) );
  NAND2X0 U113 ( .IN1(n732), .IN2(pre_sig_res_03[12]), .QN(n668) );
  NAND2X0 U114 ( .IN1(n731), .IN2(pre_sig_res_02[12]), .QN(n669) );
  NAND2X0 U115 ( .IN1(n732), .IN2(pre_sig_res_03[13]), .QN(n674) );
  NAND2X0 U116 ( .IN1(n731), .IN2(pre_sig_res_02[13]), .QN(n675) );
  NAND2X0 U117 ( .IN1(n732), .IN2(pre_sig_res_03[14]), .QN(n680) );
  NAND2X0 U118 ( .IN1(n731), .IN2(pre_sig_res_02[14]), .QN(n681) );
  NAND2X0 U119 ( .IN1(n732), .IN2(pre_sig_res_03[15]), .QN(n686) );
  NAND2X0 U120 ( .IN1(n731), .IN2(pre_sig_res_02[15]), .QN(n687) );
  NAND2X0 U121 ( .IN1(n733), .IN2(pre_sig_res_04[16]), .QN(n693) );
  NAND2X0 U122 ( .IN1(n733), .IN2(pre_sig_res_04[17]), .QN(n699) );
  NAND2X0 U123 ( .IN1(n733), .IN2(pre_sig_res_04[18]), .QN(n705) );
  NAND2X0 U124 ( .IN1(n733), .IN2(pre_sig_res_04[19]), .QN(n711) );
  NAND2X0 U125 ( .IN1(n733), .IN2(pre_sig_res_04[20]), .QN(n717) );
  NAND2X0 U126 ( .IN1(n733), .IN2(pre_sig_res_04[21]), .QN(n723) );
  NAND2X0 U127 ( .IN1(n733), .IN2(pre_sig_res_04[22]), .QN(n736) );
  NAND2X0 U128 ( .IN1(n733), .IN2(add_output_exponent_w4[0]), .QN(n597) );
  NAND2X0 U129 ( .IN1(n733), .IN2(add_output_exponent_w4[1]), .QN(n601) );
  NAND2X0 U130 ( .IN1(n733), .IN2(add_output_exponent_w4[2]), .QN(n605) );
  NAND2X0 U131 ( .IN1(n733), .IN2(add_output_exponent_w4[3]), .QN(n609) );
  NAND2X0 U132 ( .IN1(n733), .IN2(add_output_exponent_w4[4]), .QN(n613) );
  NAND2X0 U133 ( .IN1(n733), .IN2(add_output_exponent_w4[5]), .QN(n617) );
  NAND2X0 U134 ( .IN1(n733), .IN2(add_output_exponent_w4[6]), .QN(n621) );
  NAND2X0 U135 ( .IN1(n733), .IN2(add_output_exponent_w4[7]), .QN(n625) );
  NAND2X0 U136 ( .IN1(n544), .IN2(n543), .QN(N348) );
  NAND2X0 U137 ( .IN1(n561), .IN2(n822), .QN(n562) );
  NAND2X0 U138 ( .IN1(n561), .IN2(n842), .QN(n552) );
  NAND2X0 U139 ( .IN1(n561), .IN2(n844), .QN(n548) );
  NAND2X0 U140 ( .IN1(n546), .IN2(n545), .QN(N352) );
  NAND2X0 U141 ( .IN1(pre_sig_res_03[22]), .IN2(n846), .QN(n751) );
  NAND2X0 U142 ( .IN1(n835), .IN2(n750), .QN(n752) );
  NAND2X0 U143 ( .IN1(pre_sig_res_03[21]), .IN2(n846), .QN(n759) );
  NAND2X0 U144 ( .IN1(n835), .IN2(n758), .QN(n760) );
  NAND2X0 U145 ( .IN1(pre_sig_res_03[20]), .IN2(n846), .QN(n767) );
  NAND2X0 U146 ( .IN1(n835), .IN2(n766), .QN(n768) );
  NAND2X0 U147 ( .IN1(pre_sig_res_03[19]), .IN2(n846), .QN(n775) );
  NAND2X0 U148 ( .IN1(n835), .IN2(n774), .QN(n776) );
  NAND2X0 U149 ( .IN1(pre_sig_res_03[18]), .IN2(n846), .QN(n783) );
  NAND2X0 U150 ( .IN1(n835), .IN2(n782), .QN(n784) );
  NAND2X0 U151 ( .IN1(pre_sig_res_03[17]), .IN2(n846), .QN(n791) );
  NAND2X0 U152 ( .IN1(n835), .IN2(n790), .QN(n792) );
  NAND2X0 U153 ( .IN1(pre_sig_res_03[16]), .IN2(n846), .QN(n798) );
  NAND2X0 U154 ( .IN1(n835), .IN2(n815), .QN(n799) );
  NAND2X0 U155 ( .IN1(pre_sig_res_03[15]), .IN2(n846), .QN(n807) );
  NAND2X0 U156 ( .IN1(n835), .IN2(n823), .QN(n808) );
  NAND2X0 U157 ( .IN1(n742), .IN2(n749), .QN(n530) );
  NAND2X0 U158 ( .IN1(pre_sig_res_03[14]), .IN2(n78), .QN(n817) );
  NAND2X0 U159 ( .IN1(n845), .IN2(n815), .QN(n816) );
  NAND2X0 U160 ( .IN1(n835), .IN2(n814), .QN(n818) );
  NAND2X0 U161 ( .IN1(pre_sig_res_03[13]), .IN2(n846), .QN(n825) );
  NAND2X0 U162 ( .IN1(n845), .IN2(n823), .QN(n824) );
  NAND2X0 U163 ( .IN1(n835), .IN2(n822), .QN(n826) );
  NAND2X0 U164 ( .IN1(n830), .IN2(n829), .QN(n104) );
  NAND2X0 U165 ( .IN1(pre_sig_res_03[12]), .IN2(n846), .QN(n838) );
  NAND2X0 U166 ( .IN1(n835), .IN2(n842), .QN(n840) );
  NAND2X0 U167 ( .IN1(n437), .IN2(n842), .QN(n438) );
  NAND2X0 U168 ( .IN1(n442), .IN2(n823), .QN(n433) );
  NAND2X0 U169 ( .IN1(n443), .IN2(n822), .QN(n430) );
  NAND2X0 U170 ( .IN1(n429), .IN2(n428), .QN(N263) );
  NAND2X0 U171 ( .IN1(n740), .IN2(n739), .QN(n741) );
  NAND2X0 U172 ( .IN1(n51), .IN2(input_factor_02[0]), .QN(n124) );
  NAND2X0 U173 ( .IN1(n296), .IN2(input_factor_01[1]), .QN(n156) );
  NAND2X0 U174 ( .IN1(n296), .IN2(input_factor_01[2]), .QN(n185) );
  NAND2X0 U175 ( .IN1(n296), .IN2(input_factor_01[3]), .QN(n221) );
  NAND2X0 U176 ( .IN1(input_factor_01[4]), .IN2(n296), .QN(n238) );
  NAND2X0 U177 ( .IN1(input_factor_01[5]), .IN2(n296), .QN(n255) );
  NAND2X0 U178 ( .IN1(input_factor_01[6]), .IN2(n296), .QN(n274) );
  NAND2X0 U179 ( .IN1(input_factor_01[7]), .IN2(n296), .QN(n297) );
  NAND2X0 U180 ( .IN1(n358), .IN2(n357), .QN(N168) );
  NAND2X0 U181 ( .IN1(n362), .IN2(n361), .QN(N169) );
  NAND2X0 U182 ( .IN1(n366), .IN2(n365), .QN(N170) );
  NAND2X0 U183 ( .IN1(n372), .IN2(n371), .QN(N171) );
  NAND2X0 U184 ( .IN1(n378), .IN2(n377), .QN(N172) );
  NAND2X0 U185 ( .IN1(n383), .IN2(n382), .QN(N173) );
  NAND2X0 U186 ( .IN1(n390), .IN2(n389), .QN(N174) );
  NAND2X0 U187 ( .IN1(n395), .IN2(n394), .QN(N175) );
  INVX0 U188 ( .INP(n416), .ZN(n415) );
  NAND2X0 U189 ( .IN1(input_factor_01[23]), .IN2(n584), .QN(n54) );
  NOR2X0 U190 ( .IN1(n848), .IN2(n78), .QN(n849) );
  NOR2X0 U191 ( .IN1(n847), .IN2(n846), .QN(n850) );
  INVX0 U192 ( .INP(n588), .ZN(n138) );
  INVX0 U193 ( .INP(n442), .ZN(n514) );
  NOR2X0 U194 ( .IN1(n749), .IN2(n846), .QN(n835) );
  INVX0 U195 ( .INP(n843), .ZN(n833) );
  INVX0 U196 ( .INP(n822), .ZN(n834) );
  INVX0 U197 ( .INP(n823), .ZN(n812) );
  INVX0 U198 ( .INP(n790), .ZN(n803) );
  NOR2X0 U199 ( .IN1(n592), .IN2(n594), .QN(n732) );
  INVX0 U200 ( .INP(n766), .ZN(n779) );
  INVX0 U201 ( .INP(n589), .ZN(n537) );
  INVX0 U202 ( .INP(n774), .ZN(n787) );
  INVX0 U203 ( .INP(n729), .ZN(n641) );
  NOR2X0 U204 ( .IN1(n595), .IN2(n594), .QN(n734) );
  NOR2X0 U205 ( .IN1(n591), .IN2(n594), .QN(n731) );
  INVX0 U206 ( .INP(n640), .ZN(n728) );
  INVX0 U207 ( .INP(n479), .ZN(n590) );
  NAND2X0 U208 ( .IN1(exp_diff_value[2]), .IN2(n4), .QN(n225) );
  INVX0 U209 ( .INP(n397), .ZN(n726) );
  NOR2X0 U210 ( .IN1(n384), .IN2(n74), .QN(n848) );
  NOR2X0 U211 ( .IN1(exp_diff_value[1]), .IN2(exp_diff_value[0]), .QN(n391) );
  INVX0 U212 ( .INP(n213), .ZN(n199) );
  INVX0 U213 ( .INP(n211), .ZN(n198) );
  INVX0 U214 ( .INP(n296), .ZN(n379) );
  NOR2X0 U215 ( .IN1(n414), .IN2(n413), .QN(n640) );
  INVX0 U216 ( .INP(n421), .ZN(n517) );
  NOR2X0 U217 ( .IN1(add_sub_result_24_), .IN2(n418), .QN(n595) );
  MUX21X1 U218 ( .IN1(add_result[24]), .IN2(sub_result[24]), .S(n16), .Q(
        add_sub_result_24_) );
  INVX0 U219 ( .INP(n419), .ZN(n507) );
  INVX0 U220 ( .INP(n17), .ZN(n16) );
  INVX0 U221 ( .INP(n526), .ZN(n17) );
  INVX0 U222 ( .INP(n758), .ZN(n771) );
  INVX0 U223 ( .INP(n782), .ZN(n795) );
  INVX0 U224 ( .INP(n815), .ZN(n802) );
  INVX0 U225 ( .INP(n814), .ZN(n832) );
  INVX0 U226 ( .INP(n842), .ZN(n828) );
  INVX0 U227 ( .INP(n844), .ZN(n836) );
  MUX21X1 U228 ( .IN1(input_factor_01[31]), .IN2(n574), .S(input_factor_02[31]), .Q(n526) );
  INVX0 U229 ( .INP(input_factor_01[31]), .ZN(n574) );
  INVX0 U230 ( .INP(input_factor_02[22]), .ZN(n730) );
  INVX0 U231 ( .INP(n394), .ZN(n384) );
  INVX0 U232 ( .INP(input_factor_02[30]), .ZN(n740) );
  NAND4X0 U233 ( .IN1(n28), .IN2(n27), .IN3(n26), .IN4(n54), .QN(n394) );
  INVX0 U234 ( .INP(n470), .ZN(n744) );
  INVX0 U235 ( .INP(n465), .ZN(n755) );
  INVX0 U236 ( .INP(n845), .ZN(n831) );
  INVX0 U237 ( .INP(n750), .ZN(n763) );
  OR2X1 U238 ( .IN1(n586), .IN2(n779), .Q(n811) );
  NAND4X0 U239 ( .IN1(n582), .IN2(n581), .IN3(n580), .IN4(n579), .QN(n729) );
  NAND3X0 U240 ( .IN1(n517), .IN2(n424), .IN3(n488), .QN(n506) );
  NOR2X0 U241 ( .IN1(n7), .IN2(n8), .QN(n273) );
  NOR2X0 U242 ( .IN1(n388), .IN2(n270), .QN(n7) );
  NOR2X0 U243 ( .IN1(n5), .IN2(n6), .QN(n295) );
  NOR2X0 U244 ( .IN1(n290), .IN2(n291), .QN(n5) );
  NOR2X0 U245 ( .IN1(n9), .IN2(n10), .QN(n254) );
  NOR2X0 U246 ( .IN1(n270), .IN2(n381), .QN(n9) );
  NOR2X0 U247 ( .IN1(n11), .IN2(n12), .QN(n237) );
  NOR2X0 U248 ( .IN1(n376), .IN2(n270), .QN(n11) );
  INVX0 U249 ( .INP(n391), .ZN(n15) );
  NOR2X0 U250 ( .IN1(n13), .IN2(n14), .QN(n222) );
  NOR2X0 U251 ( .IN1(n709), .IN2(n212), .QN(n13) );
  INVX0 U252 ( .INP(n212), .ZN(n200) );
  MUX21X1 U253 ( .IN1(add_result[1]), .IN2(sub_result[1]), .S(n526), .Q(n842)
         );
  INVX0 U255 ( .INP(input_factor_01[30]), .ZN(n739) );
  INVX0 U256 ( .INP(input_factor_02[23]), .ZN(n584) );
  OA222X1 U257 ( .IN1(input_factor_02[30]), .IN2(n739), .IN3(n740), .IN4(
        input_factor_01[30]), .IN5(input_factor_01[23]), .IN6(n584), .Q(n28)
         );
  INVX0 U258 ( .INP(input_factor_01[24]), .ZN(n571) );
  INVX0 U259 ( .INP(n56), .ZN(n19) );
  NOR2X0 U260 ( .IN1(input_factor_02[24]), .IN2(n571), .QN(n58) );
  INVX0 U261 ( .INP(input_factor_01[28]), .ZN(n570) );
  NOR2X0 U262 ( .IN1(input_factor_02[28]), .IN2(n570), .QN(n69) );
  INVX0 U263 ( .INP(n63), .ZN(n18) );
  NOR4X0 U264 ( .IN1(n19), .IN2(n58), .IN3(n69), .IN4(n18), .QN(n27) );
  INVX0 U265 ( .INP(input_factor_01[26]), .ZN(n569) );
  NOR2X0 U266 ( .IN1(n569), .IN2(input_factor_02[26]), .QN(n59) );
  INVX0 U267 ( .INP(n59), .ZN(n21) );
  INVX0 U268 ( .INP(input_factor_01[27]), .ZN(n568) );
  NOR2X0 U269 ( .IN1(n568), .IN2(input_factor_02[27]), .QN(n66) );
  INVX0 U270 ( .INP(n66), .ZN(n20) );
  NAND4X0 U271 ( .IN1(n62), .IN2(n21), .IN3(n65), .IN4(n20), .QN(n25) );
  INVX0 U272 ( .INP(input_factor_01[29]), .ZN(n567) );
  NOR2X0 U273 ( .IN1(n567), .IN2(input_factor_02[29]), .QN(n67) );
  INVX0 U274 ( .INP(n67), .ZN(n23) );
  INVX0 U275 ( .INP(input_factor_01[25]), .ZN(n566) );
  NOR2X0 U276 ( .IN1(n566), .IN2(input_factor_02[25]), .QN(n61) );
  INVX0 U277 ( .INP(n61), .ZN(n22) );
  NAND4X0 U278 ( .IN1(n70), .IN2(n23), .IN3(n55), .IN4(n22), .QN(n24) );
  NOR2X0 U279 ( .IN1(n25), .IN2(n24), .QN(n26) );
  INVX0 U280 ( .INP(input_factor_02[21]), .ZN(n721) );
  INVX0 U281 ( .INP(input_factor_02[20]), .ZN(n715) );
  INVX0 U282 ( .INP(input_factor_02[19]), .ZN(n709) );
  INVX0 U283 ( .INP(input_factor_02[18]), .ZN(n703) );
  INVX0 U284 ( .INP(input_factor_02[17]), .ZN(n697) );
  INVX0 U285 ( .INP(input_factor_02[16]), .ZN(n691) );
  INVX0 U286 ( .INP(input_factor_02[15]), .ZN(n685) );
  INVX0 U287 ( .INP(input_factor_02[14]), .ZN(n679) );
  INVX0 U288 ( .INP(input_factor_02[13]), .ZN(n673) );
  INVX0 U289 ( .INP(input_factor_02[12]), .ZN(n667) );
  INVX0 U290 ( .INP(input_factor_02[11]), .ZN(n661) );
  INVX0 U291 ( .INP(input_factor_02[10]), .ZN(n655) );
  INVX0 U292 ( .INP(input_factor_02[9]), .ZN(n649) );
  INVX0 U293 ( .INP(input_factor_02[8]), .ZN(n645) );
  INVX0 U294 ( .INP(input_factor_02[7]), .ZN(n293) );
  INVX0 U295 ( .INP(input_factor_02[6]), .ZN(n272) );
  INVX0 U296 ( .INP(input_factor_02[5]), .ZN(n253) );
  INVX0 U297 ( .INP(input_factor_02[4]), .ZN(n236) );
  INVX0 U298 ( .INP(input_factor_02[3]), .ZN(n204) );
  INVX0 U299 ( .INP(input_factor_02[2]), .ZN(n171) );
  INVX0 U300 ( .INP(input_factor_01[0]), .ZN(n77) );
  NOR2X0 U301 ( .IN1(input_factor_02[0]), .IN2(n77), .QN(n29) );
  INVX0 U302 ( .INP(input_factor_02[1]), .ZN(n142) );
  AO222X1 U303 ( .IN1(input_factor_01[1]), .IN2(n29), .IN3(input_factor_01[1]), 
        .IN4(n142), .IN5(n29), .IN6(n142), .Q(n30) );
  AO222X1 U304 ( .IN1(input_factor_01[2]), .IN2(n171), .IN3(input_factor_01[2]), .IN4(n30), .IN5(n171), .IN6(n30), .Q(n31) );
  AO222X1 U305 ( .IN1(input_factor_01[3]), .IN2(n204), .IN3(input_factor_01[3]), .IN4(n31), .IN5(n204), .IN6(n31), .Q(n32) );
  AO222X1 U306 ( .IN1(input_factor_01[4]), .IN2(n236), .IN3(input_factor_01[4]), .IN4(n32), .IN5(n236), .IN6(n32), .Q(n33) );
  AO222X1 U307 ( .IN1(input_factor_01[5]), .IN2(n253), .IN3(input_factor_01[5]), .IN4(n33), .IN5(n253), .IN6(n33), .Q(n34) );
  AO222X1 U308 ( .IN1(input_factor_01[6]), .IN2(n272), .IN3(input_factor_01[6]), .IN4(n34), .IN5(n272), .IN6(n34), .Q(n35) );
  AO222X1 U309 ( .IN1(input_factor_01[7]), .IN2(n293), .IN3(input_factor_01[7]), .IN4(n35), .IN5(n293), .IN6(n35), .Q(n36) );
  AO222X1 U310 ( .IN1(input_factor_01[8]), .IN2(n645), .IN3(input_factor_01[8]), .IN4(n36), .IN5(n645), .IN6(n36), .Q(n37) );
  AO222X1 U311 ( .IN1(input_factor_01[9]), .IN2(n649), .IN3(input_factor_01[9]), .IN4(n37), .IN5(n649), .IN6(n37), .Q(n38) );
  AO222X1 U312 ( .IN1(input_factor_01[10]), .IN2(n655), .IN3(
        input_factor_01[10]), .IN4(n38), .IN5(n655), .IN6(n38), .Q(n39) );
  AO222X1 U313 ( .IN1(input_factor_01[11]), .IN2(n661), .IN3(
        input_factor_01[11]), .IN4(n39), .IN5(n661), .IN6(n39), .Q(n40) );
  AO222X1 U314 ( .IN1(input_factor_01[12]), .IN2(n667), .IN3(
        input_factor_01[12]), .IN4(n40), .IN5(n667), .IN6(n40), .Q(n41) );
  AO222X1 U315 ( .IN1(input_factor_01[13]), .IN2(n673), .IN3(
        input_factor_01[13]), .IN4(n41), .IN5(n673), .IN6(n41), .Q(n42) );
  AO222X1 U316 ( .IN1(input_factor_01[14]), .IN2(n679), .IN3(
        input_factor_01[14]), .IN4(n42), .IN5(n679), .IN6(n42), .Q(n43) );
  AO222X1 U317 ( .IN1(input_factor_01[15]), .IN2(n685), .IN3(
        input_factor_01[15]), .IN4(n43), .IN5(n685), .IN6(n43), .Q(n44) );
  AO222X1 U318 ( .IN1(input_factor_01[16]), .IN2(n691), .IN3(
        input_factor_01[16]), .IN4(n44), .IN5(n691), .IN6(n44), .Q(n45) );
  AO222X1 U319 ( .IN1(input_factor_01[17]), .IN2(n697), .IN3(
        input_factor_01[17]), .IN4(n45), .IN5(n697), .IN6(n45), .Q(n46) );
  AO222X1 U320 ( .IN1(input_factor_01[18]), .IN2(n703), .IN3(
        input_factor_01[18]), .IN4(n46), .IN5(n703), .IN6(n46), .Q(n47) );
  AO222X1 U321 ( .IN1(input_factor_01[19]), .IN2(n709), .IN3(
        input_factor_01[19]), .IN4(n47), .IN5(n709), .IN6(n47), .Q(n48) );
  AO222X1 U322 ( .IN1(input_factor_01[20]), .IN2(n715), .IN3(
        input_factor_01[20]), .IN4(n48), .IN5(n715), .IN6(n48), .Q(n49) );
  AO222X1 U323 ( .IN1(input_factor_01[21]), .IN2(n721), .IN3(
        input_factor_01[21]), .IN4(n49), .IN5(n721), .IN6(n49), .Q(n50) );
  AO222X1 U324 ( .IN1(input_factor_01[22]), .IN2(n730), .IN3(
        input_factor_01[22]), .IN4(n50), .IN5(n730), .IN6(n50), .Q(n76) );
  INVX0 U325 ( .INP(n396), .ZN(n51) );
  OA22X1 U326 ( .IN1(n697), .IN2(n213), .IN3(n703), .IN4(n211), .Q(n53) );
  AO222X1 U327 ( .IN1(n715), .IN2(n391), .IN3(n721), .IN4(n199), .IN5(n730), 
        .IN6(n198), .Q(n376) );
  MUX21X1 U328 ( .IN1(n222), .IN2(n376), .S(exp_diff_value[2]), .Q(n356) );
  INVX0 U329 ( .INP(n54), .ZN(n57) );
  OA221X1 U330 ( .IN1(n58), .IN2(n57), .IN3(n58), .IN4(n56), .IN5(n55), .Q(n60) );
  AO221X1 U331 ( .IN1(n62), .IN2(n61), .IN3(n62), .IN4(n60), .IN5(n59), .Q(n64) );
  OA221X1 U332 ( .IN1(n66), .IN2(n65), .IN3(n66), .IN4(n64), .IN5(n63), .Q(n68) );
  AO221X1 U333 ( .IN1(n70), .IN2(n69), .IN3(n70), .IN4(n68), .IN5(n67), .Q(n71) );
  AO222X1 U334 ( .IN1(input_factor_01[30]), .IN2(n740), .IN3(
        input_factor_01[30]), .IN4(n71), .IN5(n740), .IN6(n71), .Q(n74) );
  AO22X1 U335 ( .IN1(input_factor_01[18]), .IN2(n198), .IN3(
        input_factor_01[16]), .IN4(n391), .Q(n73) );
  AO22X1 U336 ( .IN1(input_factor_01[19]), .IN2(n200), .IN3(
        input_factor_01[17]), .IN4(n199), .Q(n72) );
  NOR2X0 U337 ( .IN1(n73), .IN2(n72), .QN(n228) );
  INVX0 U338 ( .INP(input_factor_01[22]), .ZN(n727) );
  INVX0 U339 ( .INP(input_factor_01[21]), .ZN(n720) );
  INVX0 U340 ( .INP(input_factor_01[20]), .ZN(n714) );
  AO222X1 U341 ( .IN1(n198), .IN2(n727), .IN3(n199), .IN4(n720), .IN5(n391), 
        .IN6(n714), .Q(n374) );
  MUX21X1 U342 ( .IN1(n228), .IN2(n374), .S(exp_diff_value[2]), .Q(n355) );
  INVX0 U343 ( .INP(n848), .ZN(n847) );
  OA22X1 U344 ( .IN1(n356), .IN2(n397), .IN3(n355), .IN4(n847), .Q(n79) );
  NOR3X0 U345 ( .IN1(exp_diff_value[5]), .IN2(exp_diff_value[6]), .IN3(
        exp_diff_value[7]), .QN(n75) );
  AND2X1 U346 ( .IN1(exp_diff_value[4]), .IN2(n75), .Q(n287) );
  NOR2X0 U347 ( .IN1(n394), .IN2(n76), .QN(n296) );
  OA22X1 U348 ( .IN1(n79), .IN2(n190), .IN3(n77), .IN4(n379), .Q(n123) );
  AO22X1 U349 ( .IN1(input_factor_01[10]), .IN2(n198), .IN3(input_factor_01[8]), .IN4(n391), .Q(n81) );
  AO22X1 U350 ( .IN1(input_factor_01[11]), .IN2(n200), .IN3(input_factor_01[9]), .IN4(n199), .Q(n80) );
  NOR2X0 U351 ( .IN1(n81), .IN2(n80), .QN(n230) );
  AO22X1 U352 ( .IN1(input_factor_01[14]), .IN2(n198), .IN3(
        input_factor_01[12]), .IN4(n391), .Q(n83) );
  AO22X1 U353 ( .IN1(input_factor_01[15]), .IN2(n200), .IN3(
        input_factor_01[13]), .IN4(n199), .Q(n82) );
  NOR2X0 U354 ( .IN1(n83), .IN2(n82), .QN(n229) );
  MUX21X1 U355 ( .IN1(n230), .IN2(n229), .S(exp_diff_value[2]), .Q(n303) );
  AO22X1 U356 ( .IN1(input_factor_01[2]), .IN2(n198), .IN3(input_factor_01[0]), 
        .IN4(n391), .Q(n85) );
  AO22X1 U357 ( .IN1(input_factor_01[3]), .IN2(n200), .IN3(input_factor_01[1]), 
        .IN4(n199), .Q(n84) );
  NOR2X0 U358 ( .IN1(n85), .IN2(n84), .QN(n88) );
  AO22X1 U359 ( .IN1(input_factor_01[6]), .IN2(n198), .IN3(input_factor_01[4]), 
        .IN4(n391), .Q(n87) );
  AO22X1 U360 ( .IN1(input_factor_01[7]), .IN2(n200), .IN3(input_factor_01[5]), 
        .IN4(n199), .Q(n86) );
  NOR2X0 U361 ( .IN1(n87), .IN2(n86), .QN(n231) );
  OA222X1 U362 ( .IN1(n4), .IN2(n303), .IN3(n294), .IN4(n88), .IN5(n225), 
        .IN6(n231), .Q(n121) );
  NOR4X0 U363 ( .IN1(exp_diff_value[4]), .IN2(exp_diff_value[5]), .IN3(
        exp_diff_value[6]), .IN4(exp_diff_value[7]), .QN(n393) );
  AOI22X1 U364 ( .IN1(input_factor_02[0]), .IN2(n391), .IN3(input_factor_02[2]), .IN4(n198), .QN(n90) );
  OA22X1 U365 ( .IN1(n142), .IN2(n213), .IN3(n204), .IN4(n212), .Q(n89) );
  INVX0 U366 ( .INP(n294), .ZN(n392) );
  OA22X1 U367 ( .IN1(n645), .IN2(n15), .IN3(n655), .IN4(n211), .Q(n92) );
  OA22X1 U368 ( .IN1(n649), .IN2(n213), .IN3(n661), .IN4(n212), .Q(n91) );
  OA22X1 U369 ( .IN1(n667), .IN2(n15), .IN3(n679), .IN4(n211), .Q(n116) );
  OA22X1 U370 ( .IN1(n673), .IN2(n213), .IN3(n685), .IN4(n212), .Q(n93) );
  MUX21X1 U371 ( .IN1(n226), .IN2(n224), .S(exp_diff_value[2]), .Q(n301) );
  OA22X1 U372 ( .IN1(n236), .IN2(n15), .IN3(n272), .IN4(n211), .Q(n118) );
  OA22X1 U373 ( .IN1(n253), .IN2(n213), .IN3(n293), .IN4(n212), .Q(n117) );
  INVX0 U374 ( .INP(n225), .ZN(n227) );
  AOI222X1 U375 ( .IN1(n119), .IN2(n392), .IN3(exp_diff_value[3]), .IN4(n301), 
        .IN5(n233), .IN6(n227), .QN(n120) );
  OA22X1 U376 ( .IN1(n121), .IN2(n290), .IN3(n120), .IN4(n232), .Q(n122) );
  NAND3X0 U377 ( .IN1(n124), .IN2(n123), .IN3(n122), .QN(N152) );
  AO22X1 U378 ( .IN1(input_factor_02[17]), .IN2(n391), .IN3(
        input_factor_02[19]), .IN4(n198), .Q(n126) );
  AO22X1 U379 ( .IN1(input_factor_02[18]), .IN2(n199), .IN3(
        input_factor_02[20]), .IN4(n200), .Q(n125) );
  NOR2X0 U380 ( .IN1(n126), .IN2(n125), .QN(n242) );
  AO22X1 U381 ( .IN1(input_factor_02[21]), .IN2(n1), .IN3(input_factor_02[22]), 
        .IN4(n199), .Q(n127) );
  NOR2X0 U382 ( .IN1(n198), .IN2(n127), .QN(n381) );
  MUX21X1 U383 ( .IN1(n242), .IN2(n381), .S(exp_diff_value[2]), .Q(n360) );
  AO22X1 U384 ( .IN1(input_factor_01[19]), .IN2(n198), .IN3(
        input_factor_01[17]), .IN4(n391), .Q(n129) );
  AO22X1 U385 ( .IN1(input_factor_01[20]), .IN2(n200), .IN3(
        input_factor_01[18]), .IN4(n199), .Q(n128) );
  NOR2X0 U386 ( .IN1(n129), .IN2(n128), .QN(n246) );
  AO22X1 U387 ( .IN1(input_factor_01[22]), .IN2(n199), .IN3(
        input_factor_01[21]), .IN4(n1), .Q(n130) );
  NOR2X0 U388 ( .IN1(n198), .IN2(n130), .QN(n380) );
  MUX21X1 U389 ( .IN1(n246), .IN2(n380), .S(exp_diff_value[2]), .Q(n359) );
  OA22X1 U390 ( .IN1(n397), .IN2(n360), .IN3(n847), .IN4(n359), .Q(n131) );
  OA22X1 U391 ( .IN1(n131), .IN2(n190), .IN3(n142), .IN4(n396), .Q(n155) );
  AO22X1 U392 ( .IN1(input_factor_01[11]), .IN2(n198), .IN3(input_factor_01[9]), .IN4(n391), .Q(n133) );
  AO22X1 U393 ( .IN1(input_factor_01[12]), .IN2(n200), .IN3(
        input_factor_01[10]), .IN4(n199), .Q(n132) );
  NOR2X0 U394 ( .IN1(n133), .IN2(n132), .QN(n248) );
  AO22X1 U395 ( .IN1(input_factor_01[15]), .IN2(n198), .IN3(
        input_factor_01[13]), .IN4(n391), .Q(n135) );
  AO22X1 U396 ( .IN1(input_factor_01[16]), .IN2(n200), .IN3(
        input_factor_01[14]), .IN4(n199), .Q(n134) );
  NOR2X0 U397 ( .IN1(n135), .IN2(n134), .QN(n247) );
  MUX21X1 U398 ( .IN1(n248), .IN2(n247), .S(exp_diff_value[2]), .Q(n309) );
  AO22X1 U399 ( .IN1(input_factor_01[3]), .IN2(n198), .IN3(input_factor_01[1]), 
        .IN4(n391), .Q(n137) );
  AO22X1 U400 ( .IN1(input_factor_01[4]), .IN2(n200), .IN3(input_factor_01[2]), 
        .IN4(n199), .Q(n136) );
  NOR2X0 U401 ( .IN1(n137), .IN2(n136), .QN(n141) );
  AO22X1 U402 ( .IN1(input_factor_01[7]), .IN2(n198), .IN3(input_factor_01[5]), 
        .IN4(n391), .Q(n140) );
  AO22X1 U403 ( .IN1(input_factor_01[8]), .IN2(n200), .IN3(input_factor_01[6]), 
        .IN4(n199), .Q(n139) );
  NOR2X0 U404 ( .IN1(n140), .IN2(n139), .QN(n249) );
  OA222X1 U405 ( .IN1(n4), .IN2(n309), .IN3(n294), .IN4(n141), .IN5(n225), 
        .IN6(n249), .Q(n153) );
  OA22X1 U406 ( .IN1(n142), .IN2(n15), .IN3(n204), .IN4(n211), .Q(n144) );
  OA22X1 U407 ( .IN1(n171), .IN2(n213), .IN3(n236), .IN4(n212), .Q(n143) );
  OA22X1 U408 ( .IN1(n649), .IN2(n15), .IN3(n661), .IN4(n211), .Q(n146) );
  OA22X1 U409 ( .IN1(n655), .IN2(n213), .IN3(n667), .IN4(n212), .Q(n145) );
  OA22X1 U410 ( .IN1(n673), .IN2(n15), .IN3(n685), .IN4(n211), .Q(n148) );
  OA22X1 U411 ( .IN1(n691), .IN2(n212), .IN3(n679), .IN4(n213), .Q(n147) );
  MUX21X1 U412 ( .IN1(n245), .IN2(n244), .S(exp_diff_value[2]), .Q(n307) );
  OA22X1 U413 ( .IN1(n253), .IN2(n15), .IN3(n293), .IN4(n211), .Q(n150) );
  OA22X1 U414 ( .IN1(n272), .IN2(n213), .IN3(n645), .IN4(n212), .Q(n149) );
  AOI222X1 U415 ( .IN1(n151), .IN2(n392), .IN3(exp_diff_value[3]), .IN4(n307), 
        .IN5(n250), .IN6(n227), .QN(n152) );
  OA22X1 U416 ( .IN1(n153), .IN2(n290), .IN3(n152), .IN4(n232), .Q(n154) );
  NAND3X0 U417 ( .IN1(n156), .IN2(n155), .IN3(n154), .QN(N153) );
  AO22X1 U418 ( .IN1(input_factor_02[18]), .IN2(n391), .IN3(
        input_factor_02[20]), .IN4(n198), .Q(n158) );
  AO22X1 U419 ( .IN1(input_factor_02[19]), .IN2(n199), .IN3(
        input_factor_02[21]), .IN4(n200), .Q(n157) );
  NOR2X0 U420 ( .IN1(n158), .IN2(n157), .QN(n259) );
  AO21X1 U421 ( .IN1(n730), .IN2(n1), .IN3(exp_diff_value[1]), .Q(n388) );
  MUX21X1 U422 ( .IN1(n259), .IN2(n388), .S(exp_diff_value[2]), .Q(n364) );
  AO22X1 U423 ( .IN1(input_factor_01[20]), .IN2(n198), .IN3(
        input_factor_01[18]), .IN4(n391), .Q(n160) );
  AO22X1 U424 ( .IN1(input_factor_01[21]), .IN2(n200), .IN3(
        input_factor_01[19]), .IN4(n199), .Q(n159) );
  NOR2X0 U425 ( .IN1(n160), .IN2(n159), .QN(n263) );
  AO21X1 U426 ( .IN1(n727), .IN2(n1), .IN3(exp_diff_value[1]), .Q(n386) );
  MUX21X1 U427 ( .IN1(n263), .IN2(n386), .S(exp_diff_value[2]), .Q(n363) );
  OA22X1 U428 ( .IN1(n364), .IN2(n397), .IN3(n363), .IN4(n847), .Q(n161) );
  OA22X1 U429 ( .IN1(n161), .IN2(n190), .IN3(n171), .IN4(n396), .Q(n184) );
  AO22X1 U430 ( .IN1(input_factor_01[12]), .IN2(n198), .IN3(
        input_factor_01[10]), .IN4(n391), .Q(n163) );
  AO22X1 U431 ( .IN1(input_factor_01[13]), .IN2(n200), .IN3(
        input_factor_01[11]), .IN4(n199), .Q(n162) );
  NOR2X0 U432 ( .IN1(n163), .IN2(n162), .QN(n265) );
  AO22X1 U433 ( .IN1(input_factor_01[16]), .IN2(n198), .IN3(
        input_factor_01[14]), .IN4(n391), .Q(n165) );
  AO22X1 U434 ( .IN1(input_factor_01[17]), .IN2(n200), .IN3(
        input_factor_01[15]), .IN4(n199), .Q(n164) );
  NOR2X0 U435 ( .IN1(n165), .IN2(n164), .QN(n264) );
  MUX21X1 U436 ( .IN1(n265), .IN2(n264), .S(exp_diff_value[2]), .Q(n315) );
  AO22X1 U437 ( .IN1(input_factor_01[4]), .IN2(n198), .IN3(input_factor_01[2]), 
        .IN4(n391), .Q(n167) );
  AO22X1 U438 ( .IN1(input_factor_01[5]), .IN2(n200), .IN3(input_factor_01[3]), 
        .IN4(n199), .Q(n166) );
  NOR2X0 U439 ( .IN1(n167), .IN2(n166), .QN(n170) );
  AO22X1 U440 ( .IN1(input_factor_01[8]), .IN2(n198), .IN3(input_factor_01[6]), 
        .IN4(n391), .Q(n169) );
  AO22X1 U441 ( .IN1(input_factor_01[9]), .IN2(n200), .IN3(input_factor_01[7]), 
        .IN4(n199), .Q(n168) );
  NOR2X0 U442 ( .IN1(n169), .IN2(n168), .QN(n267) );
  OA222X1 U443 ( .IN1(n4), .IN2(n315), .IN3(n294), .IN4(n170), .IN5(n225), 
        .IN6(n267), .Q(n182) );
  OA22X1 U444 ( .IN1(n171), .IN2(n15), .IN3(n236), .IN4(n211), .Q(n173) );
  OA22X1 U445 ( .IN1(n204), .IN2(n213), .IN3(n253), .IN4(n212), .Q(n172) );
  OA22X1 U446 ( .IN1(n655), .IN2(n15), .IN3(n667), .IN4(n211), .Q(n175) );
  OA22X1 U447 ( .IN1(n661), .IN2(n213), .IN3(n673), .IN4(n212), .Q(n174) );
  OA22X1 U448 ( .IN1(n691), .IN2(n211), .IN3(n679), .IN4(n15), .Q(n177) );
  OA22X1 U449 ( .IN1(n697), .IN2(n212), .IN3(n685), .IN4(n213), .Q(n176) );
  MUX21X1 U450 ( .IN1(n262), .IN2(n261), .S(exp_diff_value[2]), .Q(n313) );
  OA22X1 U451 ( .IN1(n272), .IN2(n15), .IN3(n645), .IN4(n211), .Q(n179) );
  OA22X1 U452 ( .IN1(n293), .IN2(n213), .IN3(n649), .IN4(n212), .Q(n178) );
  AOI222X1 U453 ( .IN1(n180), .IN2(n392), .IN3(exp_diff_value[3]), .IN4(n313), 
        .IN5(n268), .IN6(n227), .QN(n181) );
  OA22X1 U454 ( .IN1(n182), .IN2(n290), .IN3(n181), .IN4(n232), .Q(n183) );
  NAND3X0 U455 ( .IN1(n185), .IN2(n184), .IN3(n183), .QN(N154) );
  AO22X1 U456 ( .IN1(input_factor_02[19]), .IN2(n391), .IN3(
        input_factor_02[21]), .IN4(n198), .Q(n187) );
  AO22X1 U457 ( .IN1(input_factor_02[20]), .IN2(n199), .IN3(
        input_factor_02[22]), .IN4(n200), .Q(n186) );
  NOR2X0 U458 ( .IN1(n187), .IN2(n186), .QN(n278) );
  MUX21X1 U459 ( .IN1(n278), .IN2(n15), .S(exp_diff_value[2]), .Q(n370) );
  AO22X1 U460 ( .IN1(input_factor_01[21]), .IN2(n198), .IN3(
        input_factor_01[19]), .IN4(n391), .Q(n189) );
  AO22X1 U461 ( .IN1(input_factor_01[22]), .IN2(n200), .IN3(
        input_factor_01[20]), .IN4(n199), .Q(n188) );
  NOR2X0 U462 ( .IN1(n189), .IN2(n188), .QN(n283) );
  MUX21X1 U463 ( .IN1(n283), .IN2(n15), .S(exp_diff_value[2]), .Q(n368) );
  OA22X1 U464 ( .IN1(n370), .IN2(n397), .IN3(n368), .IN4(n847), .Q(n191) );
  OA22X1 U465 ( .IN1(n191), .IN2(n190), .IN3(n204), .IN4(n396), .Q(n220) );
  AO22X1 U466 ( .IN1(input_factor_01[13]), .IN2(n198), .IN3(
        input_factor_01[11]), .IN4(n391), .Q(n193) );
  AO22X1 U467 ( .IN1(input_factor_01[14]), .IN2(n200), .IN3(
        input_factor_01[12]), .IN4(n199), .Q(n192) );
  NOR2X0 U468 ( .IN1(n193), .IN2(n192), .QN(n286) );
  AO22X1 U469 ( .IN1(input_factor_01[17]), .IN2(n198), .IN3(
        input_factor_01[15]), .IN4(n391), .Q(n195) );
  AO22X1 U470 ( .IN1(input_factor_01[18]), .IN2(n200), .IN3(
        input_factor_01[16]), .IN4(n199), .Q(n194) );
  NOR2X0 U471 ( .IN1(n195), .IN2(n194), .QN(n284) );
  MUX21X1 U472 ( .IN1(n286), .IN2(n284), .S(exp_diff_value[2]), .Q(n321) );
  AO22X1 U473 ( .IN1(input_factor_01[5]), .IN2(n198), .IN3(input_factor_01[3]), 
        .IN4(n391), .Q(n197) );
  AO22X1 U474 ( .IN1(input_factor_01[6]), .IN2(n200), .IN3(input_factor_01[4]), 
        .IN4(n199), .Q(n196) );
  NOR2X0 U475 ( .IN1(n197), .IN2(n196), .QN(n203) );
  AO22X1 U476 ( .IN1(input_factor_01[9]), .IN2(n198), .IN3(input_factor_01[7]), 
        .IN4(n391), .Q(n202) );
  AO22X1 U477 ( .IN1(input_factor_01[10]), .IN2(n200), .IN3(input_factor_01[8]), .IN4(n199), .Q(n201) );
  NOR2X0 U478 ( .IN1(n202), .IN2(n201), .QN(n291) );
  OA222X1 U479 ( .IN1(n4), .IN2(n321), .IN3(n294), .IN4(n203), .IN5(n225), 
        .IN6(n291), .Q(n218) );
  OA22X1 U480 ( .IN1(n204), .IN2(n15), .IN3(n253), .IN4(n211), .Q(n206) );
  OA22X1 U481 ( .IN1(n236), .IN2(n213), .IN3(n272), .IN4(n212), .Q(n205) );
  OA22X1 U482 ( .IN1(n661), .IN2(n15), .IN3(n673), .IN4(n211), .Q(n208) );
  OA22X1 U483 ( .IN1(n667), .IN2(n213), .IN3(n679), .IN4(n212), .Q(n207) );
  OA22X1 U484 ( .IN1(n697), .IN2(n211), .IN3(n685), .IN4(n15), .Q(n210) );
  OA22X1 U485 ( .IN1(n691), .IN2(n213), .IN3(n703), .IN4(n212), .Q(n209) );
  MUX21X1 U486 ( .IN1(n281), .IN2(n280), .S(exp_diff_value[2]), .Q(n319) );
  OA22X1 U487 ( .IN1(n293), .IN2(n15), .IN3(n649), .IN4(n211), .Q(n215) );
  OA22X1 U488 ( .IN1(n645), .IN2(n213), .IN3(n655), .IN4(n212), .Q(n214) );
  AOI222X1 U489 ( .IN1(n216), .IN2(n392), .IN3(exp_diff_value[3]), .IN4(n319), 
        .IN5(n288), .IN6(n227), .QN(n217) );
  OA22X1 U490 ( .IN1(n218), .IN2(n290), .IN3(n217), .IN4(n232), .Q(n219) );
  NAND3X0 U491 ( .IN1(n221), .IN2(n220), .IN3(n219), .QN(N155) );
  INVX0 U492 ( .INP(n222), .ZN(n223) );
  MUX21X1 U493 ( .IN1(n224), .IN2(n223), .S(exp_diff_value[2]), .Q(n325) );
  NOR2X0 U494 ( .IN1(n4), .IN2(n232), .QN(n328) );
  NOR2X0 U495 ( .IN1(n225), .IN2(n232), .QN(n282) );
  AOI22X1 U496 ( .IN1(n325), .IN2(n328), .IN3(n282), .IN4(n226), .QN(n241) );
  INVX0 U497 ( .INP(n290), .ZN(n373) );
  MUX21X1 U498 ( .IN1(n229), .IN2(n228), .S(exp_diff_value[2]), .Q(n327) );
  OA22X1 U499 ( .IN1(n230), .IN2(n285), .IN3(n327), .IN4(n349), .Q(n240) );
  OA22X1 U500 ( .IN1(n231), .IN2(n290), .IN3(n374), .IN4(n266), .Q(n235) );
  INVX0 U501 ( .INP(n232), .ZN(n375) );
  OA22X1 U502 ( .IN1(n237), .IN2(n294), .IN3(n236), .IN4(n396), .Q(n239) );
  NAND4X0 U503 ( .IN1(n241), .IN2(n240), .IN3(n239), .IN4(n238), .QN(N156) );
  INVX0 U504 ( .INP(n242), .ZN(n243) );
  MUX21X1 U505 ( .IN1(n244), .IN2(n243), .S(exp_diff_value[2]), .Q(n332) );
  AOI22X1 U506 ( .IN1(n332), .IN2(n328), .IN3(n282), .IN4(n245), .QN(n258) );
  MUX21X1 U507 ( .IN1(n247), .IN2(n246), .S(exp_diff_value[2]), .Q(n334) );
  OA22X1 U508 ( .IN1(n248), .IN2(n285), .IN3(n334), .IN4(n349), .Q(n257) );
  OA22X1 U509 ( .IN1(n380), .IN2(n266), .IN3(n249), .IN4(n290), .Q(n252) );
  OA22X1 U510 ( .IN1(n254), .IN2(n294), .IN3(n253), .IN4(n396), .Q(n256) );
  NAND4X0 U511 ( .IN1(n258), .IN2(n257), .IN3(n256), .IN4(n255), .QN(N157) );
  INVX0 U512 ( .INP(n259), .ZN(n260) );
  MUX21X1 U513 ( .IN1(n261), .IN2(n260), .S(exp_diff_value[2]), .Q(n338) );
  AOI22X1 U514 ( .IN1(n338), .IN2(n328), .IN3(n282), .IN4(n262), .QN(n277) );
  MUX21X1 U515 ( .IN1(n264), .IN2(n263), .S(exp_diff_value[2]), .Q(n340) );
  OA22X1 U516 ( .IN1(n265), .IN2(n285), .IN3(n340), .IN4(n349), .Q(n276) );
  OA22X1 U517 ( .IN1(n267), .IN2(n290), .IN3(n386), .IN4(n266), .Q(n271) );
  OA22X1 U518 ( .IN1(n273), .IN2(n294), .IN3(n272), .IN4(n396), .Q(n275) );
  NAND4X0 U519 ( .IN1(n277), .IN2(n276), .IN3(n275), .IN4(n274), .QN(N158) );
  INVX0 U520 ( .INP(n278), .ZN(n279) );
  MUX21X1 U521 ( .IN1(n280), .IN2(n279), .S(exp_diff_value[2]), .Q(n346) );
  AOI22X1 U522 ( .IN1(n346), .IN2(n328), .IN3(n282), .IN4(n281), .QN(n300) );
  MUX21X1 U523 ( .IN1(n284), .IN2(n283), .S(exp_diff_value[2]), .Q(n348) );
  OA22X1 U524 ( .IN1(n286), .IN2(n285), .IN3(n348), .IN4(n349), .Q(n299) );
  NAND3X0 U525 ( .IN1(n287), .IN2(n391), .IN3(n394), .QN(n292) );
  OA22X1 U526 ( .IN1(n295), .IN2(n294), .IN3(n293), .IN4(n396), .Q(n298) );
  NAND4X0 U527 ( .IN1(n300), .IN2(n299), .IN3(n298), .IN4(n297), .QN(N159) );
  INVX0 U528 ( .INP(n328), .ZN(n350) );
  OA22X1 U529 ( .IN1(n355), .IN2(n349), .IN3(n356), .IN4(n350), .Q(n306) );
  INVX0 U530 ( .INP(n301), .ZN(n302) );
  OA22X1 U531 ( .IN1(n303), .IN2(n367), .IN3(n302), .IN4(n369), .Q(n305) );
  INVX0 U532 ( .INP(input_factor_01[8]), .ZN(n644) );
  OA22X1 U533 ( .IN1(n645), .IN2(n396), .IN3(n644), .IN4(n379), .Q(n304) );
  NAND3X0 U534 ( .IN1(n306), .IN2(n305), .IN3(n304), .QN(N160) );
  OA22X1 U535 ( .IN1(n360), .IN2(n350), .IN3(n359), .IN4(n349), .Q(n312) );
  INVX0 U536 ( .INP(n307), .ZN(n308) );
  OA22X1 U537 ( .IN1(n309), .IN2(n367), .IN3(n308), .IN4(n369), .Q(n311) );
  INVX0 U538 ( .INP(input_factor_01[9]), .ZN(n648) );
  OA22X1 U539 ( .IN1(n649), .IN2(n396), .IN3(n648), .IN4(n379), .Q(n310) );
  NAND3X0 U540 ( .IN1(n312), .IN2(n311), .IN3(n310), .QN(N161) );
  OA22X1 U541 ( .IN1(n363), .IN2(n349), .IN3(n364), .IN4(n350), .Q(n318) );
  INVX0 U542 ( .INP(n313), .ZN(n314) );
  OA22X1 U543 ( .IN1(n315), .IN2(n367), .IN3(n314), .IN4(n369), .Q(n317) );
  INVX0 U544 ( .INP(input_factor_01[10]), .ZN(n654) );
  OA22X1 U545 ( .IN1(n655), .IN2(n396), .IN3(n654), .IN4(n379), .Q(n316) );
  NAND3X0 U546 ( .IN1(n318), .IN2(n317), .IN3(n316), .QN(N162) );
  OA22X1 U547 ( .IN1(n368), .IN2(n349), .IN3(n370), .IN4(n350), .Q(n324) );
  INVX0 U548 ( .INP(n319), .ZN(n320) );
  OA22X1 U549 ( .IN1(n321), .IN2(n367), .IN3(n320), .IN4(n369), .Q(n323) );
  INVX0 U550 ( .INP(input_factor_01[11]), .ZN(n660) );
  OA22X1 U551 ( .IN1(n661), .IN2(n396), .IN3(n660), .IN4(n379), .Q(n322) );
  NAND3X0 U552 ( .IN1(n324), .IN2(n323), .IN3(n322), .QN(N163) );
  INVX0 U553 ( .INP(n325), .ZN(n326) );
  OA22X1 U554 ( .IN1(n327), .IN2(n367), .IN3(n326), .IN4(n369), .Q(n331) );
  OR2X1 U555 ( .IN1(n349), .IN2(exp_diff_value[2]), .Q(n341) );
  OA22X1 U556 ( .IN1(n376), .IN2(n342), .IN3(n374), .IN4(n341), .Q(n330) );
  INVX0 U557 ( .INP(input_factor_01[12]), .ZN(n666) );
  OA22X1 U558 ( .IN1(n667), .IN2(n396), .IN3(n666), .IN4(n379), .Q(n329) );
  NAND3X0 U559 ( .IN1(n331), .IN2(n330), .IN3(n329), .QN(N164) );
  INVX0 U560 ( .INP(n332), .ZN(n333) );
  OA22X1 U561 ( .IN1(n334), .IN2(n367), .IN3(n333), .IN4(n369), .Q(n337) );
  OA22X1 U562 ( .IN1(n380), .IN2(n341), .IN3(n381), .IN4(n342), .Q(n336) );
  INVX0 U563 ( .INP(input_factor_01[13]), .ZN(n672) );
  OA22X1 U564 ( .IN1(n673), .IN2(n396), .IN3(n672), .IN4(n379), .Q(n335) );
  NAND3X0 U565 ( .IN1(n337), .IN2(n336), .IN3(n335), .QN(N165) );
  INVX0 U566 ( .INP(n338), .ZN(n339) );
  OA22X1 U567 ( .IN1(n340), .IN2(n367), .IN3(n339), .IN4(n369), .Q(n345) );
  OA22X1 U568 ( .IN1(n388), .IN2(n342), .IN3(n386), .IN4(n341), .Q(n344) );
  INVX0 U569 ( .INP(input_factor_01[14]), .ZN(n678) );
  OA22X1 U570 ( .IN1(n679), .IN2(n396), .IN3(n678), .IN4(n379), .Q(n343) );
  NAND3X0 U571 ( .IN1(n345), .IN2(n344), .IN3(n343), .QN(N166) );
  INVX0 U572 ( .INP(n346), .ZN(n347) );
  OA22X1 U573 ( .IN1(n348), .IN2(n367), .IN3(n347), .IN4(n369), .Q(n354) );
  INVX0 U574 ( .INP(input_factor_01[15]), .ZN(n684) );
  OA22X1 U575 ( .IN1(n685), .IN2(n396), .IN3(n684), .IN4(n379), .Q(n353) );
  NAND3X0 U576 ( .IN1(n351), .IN2(n2), .IN3(n391), .QN(n352) );
  NAND3X0 U577 ( .IN1(n354), .IN2(n353), .IN3(n352), .QN(N167) );
  INVX0 U578 ( .INP(input_factor_01[16]), .ZN(n690) );
  OA22X1 U579 ( .IN1(n355), .IN2(n367), .IN3(n690), .IN4(n379), .Q(n358) );
  OA22X1 U580 ( .IN1(n356), .IN2(n369), .IN3(n691), .IN4(n396), .Q(n357) );
  INVX0 U581 ( .INP(input_factor_01[17]), .ZN(n696) );
  OA22X1 U582 ( .IN1(n696), .IN2(n379), .IN3(n359), .IN4(n367), .Q(n362) );
  OA22X1 U583 ( .IN1(n697), .IN2(n396), .IN3(n360), .IN4(n369), .Q(n361) );
  INVX0 U584 ( .INP(input_factor_01[18]), .ZN(n702) );
  OA22X1 U585 ( .IN1(n363), .IN2(n367), .IN3(n702), .IN4(n379), .Q(n366) );
  OA22X1 U586 ( .IN1(n364), .IN2(n369), .IN3(n703), .IN4(n396), .Q(n365) );
  INVX0 U587 ( .INP(input_factor_01[19]), .ZN(n708) );
  OA22X1 U588 ( .IN1(n368), .IN2(n367), .IN3(n708), .IN4(n379), .Q(n372) );
  OA22X1 U589 ( .IN1(n370), .IN2(n369), .IN3(n709), .IN4(n396), .Q(n371) );
  OA22X1 U590 ( .IN1(n714), .IN2(n379), .IN3(n374), .IN4(n385), .Q(n378) );
  OA22X1 U591 ( .IN1(n715), .IN2(n396), .IN3(n376), .IN4(n387), .Q(n377) );
  OA22X1 U592 ( .IN1(n380), .IN2(n385), .IN3(n720), .IN4(n379), .Q(n383) );
  OA22X1 U593 ( .IN1(n381), .IN2(n387), .IN3(n721), .IN4(n396), .Q(n382) );
  NAND3X0 U594 ( .IN1(input_factor_01[22]), .IN2(input_factor_02[22]), .IN3(
        n384), .QN(n390) );
  OA22X1 U595 ( .IN1(n388), .IN2(n387), .IN3(n386), .IN4(n385), .Q(n389) );
  NAND3X0 U596 ( .IN1(n393), .IN2(n392), .IN3(n391), .QN(n395) );
  MUX21X1 U597 ( .IN1(input_factor_01[0]), .IN2(input_factor_02[0]), .S(n415), 
        .Q(N176) );
  MUX21X1 U598 ( .IN1(input_factor_01[1]), .IN2(input_factor_02[1]), .S(n415), 
        .Q(N177) );
  MUX21X1 U599 ( .IN1(input_factor_01[2]), .IN2(input_factor_02[2]), .S(n415), 
        .Q(N178) );
  MUX21X1 U600 ( .IN1(input_factor_01[3]), .IN2(input_factor_02[3]), .S(n415), 
        .Q(N179) );
  MUX21X1 U601 ( .IN1(input_factor_01[4]), .IN2(input_factor_02[4]), .S(n415), 
        .Q(N180) );
  MUX21X1 U602 ( .IN1(input_factor_01[5]), .IN2(input_factor_02[5]), .S(n415), 
        .Q(N181) );
  MUX21X1 U603 ( .IN1(input_factor_01[6]), .IN2(input_factor_02[6]), .S(n415), 
        .Q(N182) );
  MUX21X1 U604 ( .IN1(input_factor_01[7]), .IN2(input_factor_02[7]), .S(n415), 
        .Q(N183) );
  MUX21X1 U605 ( .IN1(input_factor_01[8]), .IN2(input_factor_02[8]), .S(n415), 
        .Q(N184) );
  MUX21X1 U606 ( .IN1(input_factor_01[9]), .IN2(input_factor_02[9]), .S(n415), 
        .Q(N185) );
  MUX21X1 U607 ( .IN1(input_factor_01[10]), .IN2(input_factor_02[10]), .S(n415), .Q(N186) );
  MUX21X1 U608 ( .IN1(input_factor_01[11]), .IN2(input_factor_02[11]), .S(n415), .Q(N187) );
  MUX21X1 U609 ( .IN1(input_factor_01[12]), .IN2(input_factor_02[12]), .S(n415), .Q(N188) );
  MUX21X1 U610 ( .IN1(input_factor_01[13]), .IN2(input_factor_02[13]), .S(n415), .Q(N189) );
  MUX21X1 U611 ( .IN1(input_factor_01[14]), .IN2(input_factor_02[14]), .S(n415), .Q(N190) );
  MUX21X1 U612 ( .IN1(input_factor_01[15]), .IN2(input_factor_02[15]), .S(n415), .Q(N191) );
  MUX21X1 U613 ( .IN1(input_factor_01[16]), .IN2(input_factor_02[16]), .S(n415), .Q(N192) );
  MUX21X1 U614 ( .IN1(input_factor_01[17]), .IN2(input_factor_02[17]), .S(n415), .Q(N193) );
  MUX21X1 U615 ( .IN1(input_factor_01[18]), .IN2(input_factor_02[18]), .S(n415), .Q(N194) );
  MUX21X1 U616 ( .IN1(input_factor_01[19]), .IN2(input_factor_02[19]), .S(n415), .Q(N195) );
  MUX21X1 U617 ( .IN1(input_factor_01[20]), .IN2(input_factor_02[20]), .S(n415), .Q(N196) );
  MUX21X1 U618 ( .IN1(input_factor_01[21]), .IN2(input_factor_02[21]), .S(n415), .Q(N197) );
  MUX21X1 U619 ( .IN1(input_factor_01[22]), .IN2(input_factor_02[22]), .S(n415), .Q(N198) );
  MUX21X1 U620 ( .IN1(add_result[0]), .IN2(sub_result[0]), .S(n526), .Q(n844)
         );
  MUX21X1 U621 ( .IN1(add_result[2]), .IN2(sub_result[2]), .S(n526), .Q(n822)
         );
  MUX21X1 U622 ( .IN1(add_result[3]), .IN2(sub_result[3]), .S(n526), .Q(n814)
         );
  MUX21X1 U623 ( .IN1(add_result[4]), .IN2(sub_result[4]), .S(n526), .Q(n823)
         );
  MUX21X1 U624 ( .IN1(add_result[5]), .IN2(sub_result[5]), .S(n526), .Q(n815)
         );
  MUX21X1 U625 ( .IN1(add_result[6]), .IN2(sub_result[6]), .S(n526), .Q(n790)
         );
  MUX21X1 U626 ( .IN1(add_result[7]), .IN2(sub_result[7]), .S(n526), .Q(n782)
         );
  MUX21X1 U627 ( .IN1(add_result[9]), .IN2(sub_result[9]), .S(n526), .Q(n766)
         );
  MUX21X1 U628 ( .IN1(add_result[10]), .IN2(sub_result[10]), .S(n526), .Q(n758) );
  NOR4X0 U629 ( .IN1(n526), .IN2(add_result[14]), .IN3(add_result[15]), .IN4(
        add_result[13]), .QN(n535) );
  NOR4X0 U630 ( .IN1(sub_result[15]), .IN2(sub_result[14]), .IN3(
        sub_result[13]), .IN4(n17), .QN(n533) );
  NOR2X0 U631 ( .IN1(n535), .IN2(n533), .QN(n401) );
  MUX21X1 U632 ( .IN1(add_result[11]), .IN2(sub_result[11]), .S(n526), .Q(n750) );
  MUX21X1 U633 ( .IN1(add_result[16]), .IN2(sub_result[16]), .S(n16), .Q(n419)
         );
  MUX21X1 U634 ( .IN1(add_result[17]), .IN2(sub_result[17]), .S(n16), .Q(n488)
         );
  MUX21X1 U635 ( .IN1(add_result[20]), .IN2(sub_result[20]), .S(n16), .Q(n422)
         );
  INVX0 U636 ( .INP(n422), .ZN(n515) );
  MUX21X1 U637 ( .IN1(add_result[22]), .IN2(sub_result[22]), .S(n16), .Q(n423)
         );
  INVX0 U638 ( .INP(n423), .ZN(n398) );
  MUX21X1 U639 ( .IN1(add_result[23]), .IN2(sub_result[23]), .S(n16), .Q(n418)
         );
  MUX21X1 U640 ( .IN1(add_result[21]), .IN2(sub_result[21]), .S(n16), .Q(n425)
         );
  NOR2X0 U641 ( .IN1(n426), .IN2(n425), .QN(n427) );
  MUX21X1 U642 ( .IN1(add_result[19]), .IN2(sub_result[19]), .S(n16), .Q(n497)
         );
  NOR2X0 U643 ( .IN1(n399), .IN2(n497), .QN(n424) );
  MUX21X1 U644 ( .IN1(add_result[18]), .IN2(sub_result[18]), .S(n16), .Q(n421)
         );
  NOR2X0 U645 ( .IN1(n488), .IN2(n400), .QN(n420) );
  MUX21X1 U646 ( .IN1(add_result[12]), .IN2(sub_result[12]), .S(n16), .Q(n465)
         );
  NOR4X0 U647 ( .IN1(n401), .IN2(n750), .IN3(n589), .IN4(n465), .QN(n745) );
  MUX21X1 U648 ( .IN1(add_result[8]), .IN2(sub_result[8]), .S(n16), .Q(n774)
         );
  NOR3X0 U649 ( .IN1(n766), .IN2(n586), .IN3(n774), .QN(n540) );
  NOR2X0 U650 ( .IN1(n790), .IN2(n402), .QN(n539) );
  NOR2X0 U651 ( .IN1(n823), .IN2(n403), .QN(n547) );
  NOR2X0 U652 ( .IN1(n822), .IN2(n404), .QN(n541) );
  NAND3X0 U653 ( .IN1(n836), .IN2(n828), .IN3(n541), .QN(n587) );
  NOR4X0 U654 ( .IN1(input_factor_02[4]), .IN2(input_factor_02[5]), .IN3(
        input_factor_02[6]), .IN4(input_factor_02[7]), .QN(n408) );
  NOR4X0 U655 ( .IN1(input_factor_02[0]), .IN2(input_factor_02[1]), .IN3(
        input_factor_02[2]), .IN4(input_factor_02[3]), .QN(n407) );
  NOR4X0 U656 ( .IN1(input_factor_02[12]), .IN2(input_factor_02[13]), .IN3(
        input_factor_02[14]), .IN4(input_factor_02[15]), .QN(n406) );
  NOR4X0 U657 ( .IN1(input_factor_02[8]), .IN2(input_factor_02[9]), .IN3(
        input_factor_02[10]), .IN4(input_factor_02[11]), .QN(n405) );
  NAND4X0 U658 ( .IN1(n408), .IN2(n407), .IN3(n406), .IN4(n405), .QN(n414) );
  NOR4X0 U659 ( .IN1(input_factor_02[26]), .IN2(input_factor_02[27]), .IN3(
        input_factor_02[30]), .IN4(input_factor_02[25]), .QN(n412) );
  NOR4X0 U660 ( .IN1(input_factor_02[29]), .IN2(input_factor_02[23]), .IN3(
        input_factor_02[24]), .IN4(input_factor_02[28]), .QN(n411) );
  NOR4X0 U661 ( .IN1(input_factor_02[19]), .IN2(input_factor_02[20]), .IN3(
        input_factor_02[21]), .IN4(input_factor_02[22]), .QN(n410) );
  NOR4X0 U662 ( .IN1(input_factor_02[31]), .IN2(input_factor_02[16]), .IN3(
        input_factor_02[17]), .IN4(input_factor_02[18]), .QN(n409) );
  NAND4X0 U663 ( .IN1(n412), .IN2(n411), .IN3(n410), .IN4(n409), .QN(n413) );
  AO222X1 U664 ( .IN1(input_factor_01[31]), .IN2(n640), .IN3(
        input_factor_01[31]), .IN4(n416), .IN5(n415), .IN6(input_factor_02[31]), .Q(n417) );
  AND2X1 U665 ( .IN1(n587), .IN2(n417), .Q(N211) );
  MUX21X1 U666 ( .IN1(n844), .IN2(n842), .S(add_sub_result_24_), .Q(N226) );
  MUX21X1 U667 ( .IN1(n842), .IN2(n822), .S(add_sub_result_24_), .Q(N227) );
  MUX21X1 U668 ( .IN1(n822), .IN2(n814), .S(add_sub_result_24_), .Q(N228) );
  MUX21X1 U669 ( .IN1(n814), .IN2(n823), .S(add_sub_result_24_), .Q(N229) );
  MUX21X1 U670 ( .IN1(n823), .IN2(n815), .S(add_sub_result_24_), .Q(N230) );
  MUX21X1 U671 ( .IN1(n815), .IN2(n790), .S(add_sub_result_24_), .Q(N231) );
  MUX21X1 U672 ( .IN1(n790), .IN2(n782), .S(add_sub_result_24_), .Q(N232) );
  MUX21X1 U673 ( .IN1(n782), .IN2(n774), .S(add_sub_result_24_), .Q(N233) );
  MUX21X1 U674 ( .IN1(n774), .IN2(n766), .S(add_sub_result_24_), .Q(N234) );
  MUX21X1 U675 ( .IN1(n766), .IN2(n758), .S(add_sub_result_24_), .Q(N235) );
  MUX21X1 U676 ( .IN1(n758), .IN2(n750), .S(add_sub_result_24_), .Q(N236) );
  MUX21X1 U677 ( .IN1(n750), .IN2(n465), .S(add_sub_result_24_), .Q(N237) );
  MUX21X1 U678 ( .IN1(add_result[13]), .IN2(sub_result[13]), .S(n16), .Q(n470)
         );
  MUX21X1 U679 ( .IN1(n465), .IN2(n470), .S(add_sub_result_24_), .Q(N238) );
  MUX21X1 U680 ( .IN1(add_result[14]), .IN2(sub_result[14]), .S(n16), .Q(n524)
         );
  MUX21X1 U681 ( .IN1(n470), .IN2(n524), .S(add_sub_result_24_), .Q(N239) );
  MUX21X1 U682 ( .IN1(add_result[15]), .IN2(sub_result[15]), .S(n16), .Q(n479)
         );
  MUX21X1 U683 ( .IN1(n524), .IN2(n479), .S(add_sub_result_24_), .Q(N240) );
  MUX21X1 U684 ( .IN1(n479), .IN2(n419), .S(add_sub_result_24_), .Q(N241) );
  MUX21X1 U685 ( .IN1(n419), .IN2(n488), .S(add_sub_result_24_), .Q(N242) );
  MUX21X1 U686 ( .IN1(n488), .IN2(n421), .S(add_sub_result_24_), .Q(N243) );
  MUX21X1 U687 ( .IN1(n421), .IN2(n497), .S(add_sub_result_24_), .Q(N244) );
  MUX21X1 U688 ( .IN1(n497), .IN2(n422), .S(add_sub_result_24_), .Q(N245) );
  MUX21X1 U689 ( .IN1(n422), .IN2(n425), .S(add_sub_result_24_), .Q(N246) );
  MUX21X1 U690 ( .IN1(n425), .IN2(n423), .S(add_sub_result_24_), .Q(N247) );
  MUX21X1 U691 ( .IN1(n423), .IN2(n418), .S(add_sub_result_24_), .Q(N248) );
  NAND4X0 U692 ( .IN1(n519), .IN2(n508), .IN3(n512), .IN4(n510), .QN(N256) );
  INVX0 U693 ( .INP(n425), .ZN(n511) );
  NOR2X0 U694 ( .IN1(n511), .IN2(n426), .QN(n442) );
  NAND4X0 U695 ( .IN1(n519), .IN2(n506), .IN3(n512), .IN4(n514), .QN(N257) );
  NAND3X0 U696 ( .IN1(n427), .IN2(n515), .IN3(n497), .QN(n516) );
  NAND4X0 U697 ( .IN1(n519), .IN2(n508), .IN3(n516), .IN4(n506), .QN(N258) );
  NOR2X0 U698 ( .IN1(n836), .IN2(n510), .QN(N260) );
  INVX0 U699 ( .INP(n510), .ZN(n444) );
  AO22X1 U700 ( .IN1(n444), .IN2(n842), .IN3(n442), .IN4(n844), .Q(N261) );
  INVX0 U701 ( .INP(n512), .ZN(n443) );
  AO222X1 U702 ( .IN1(n844), .IN2(n443), .IN3(n842), .IN4(n442), .IN5(n822), 
        .IN6(n444), .Q(N262) );
  OA22X1 U703 ( .IN1(n828), .IN2(n512), .IN3(n836), .IN4(n516), .Q(n429) );
  OA22X1 U704 ( .IN1(n834), .IN2(n514), .IN3(n832), .IN4(n510), .Q(n428) );
  OA22X1 U705 ( .IN1(n812), .IN2(n510), .IN3(n832), .IN4(n514), .Q(n432) );
  OA22X1 U706 ( .IN1(n828), .IN2(n516), .IN3(n836), .IN4(n508), .Q(n431) );
  NAND3X0 U707 ( .IN1(n432), .IN2(n431), .IN3(n430), .QN(N264) );
  OA22X1 U708 ( .IN1(n802), .IN2(n510), .IN3(n832), .IN4(n512), .Q(n436) );
  OA22X1 U709 ( .IN1(n834), .IN2(n516), .IN3(n828), .IN4(n508), .Q(n435) );
  INVX0 U710 ( .INP(n506), .ZN(n437) );
  NAND4X0 U711 ( .IN1(n436), .IN2(n435), .IN3(n434), .IN4(n433), .QN(N265) );
  OA22X1 U712 ( .IN1(n812), .IN2(n512), .IN3(n832), .IN4(n516), .Q(n441) );
  OA22X1 U713 ( .IN1(n803), .IN2(n510), .IN3(n802), .IN4(n514), .Q(n440) );
  OA22X1 U714 ( .IN1(n834), .IN2(n508), .IN3(n836), .IN4(n519), .Q(n439) );
  NAND4X0 U715 ( .IN1(n441), .IN2(n440), .IN3(n439), .IN4(n438), .QN(N266) );
  NOR4X0 U716 ( .IN1(n444), .IN2(n443), .IN3(n442), .IN4(N258), .QN(n588) );
  OA22X1 U717 ( .IN1(n834), .IN2(n506), .IN3(n832), .IN4(n508), .Q(n448) );
  OA22X1 U718 ( .IN1(n795), .IN2(n510), .IN3(n802), .IN4(n512), .Q(n447) );
  OA22X1 U719 ( .IN1(n803), .IN2(n514), .IN3(n812), .IN4(n516), .Q(n446) );
  OA22X1 U720 ( .IN1(n828), .IN2(n519), .IN3(n836), .IN4(n138), .Q(n445) );
  NAND4X0 U721 ( .IN1(n448), .IN2(n447), .IN3(n446), .IN4(n445), .QN(N267) );
  OA22X1 U722 ( .IN1(n812), .IN2(n508), .IN3(n832), .IN4(n506), .Q(n452) );
  OA22X1 U723 ( .IN1(n787), .IN2(n510), .IN3(n803), .IN4(n512), .Q(n451) );
  OA22X1 U724 ( .IN1(n795), .IN2(n514), .IN3(n802), .IN4(n516), .Q(n450) );
  OA22X1 U725 ( .IN1(n834), .IN2(n519), .IN3(n828), .IN4(n138), .Q(n449) );
  NAND4X0 U726 ( .IN1(n452), .IN2(n451), .IN3(n450), .IN4(n449), .QN(N268) );
  OA22X1 U727 ( .IN1(n802), .IN2(n508), .IN3(n812), .IN4(n506), .Q(n456) );
  OA22X1 U728 ( .IN1(n779), .IN2(n510), .IN3(n795), .IN4(n512), .Q(n455) );
  OA22X1 U729 ( .IN1(n787), .IN2(n514), .IN3(n803), .IN4(n516), .Q(n454) );
  OA22X1 U730 ( .IN1(n834), .IN2(n138), .IN3(n832), .IN4(n519), .Q(n453) );
  NAND4X0 U731 ( .IN1(n456), .IN2(n455), .IN3(n454), .IN4(n453), .QN(N269) );
  OA22X1 U732 ( .IN1(n803), .IN2(n508), .IN3(n802), .IN4(n506), .Q(n460) );
  OA22X1 U733 ( .IN1(n787), .IN2(n512), .IN3(n771), .IN4(n510), .Q(n459) );
  OA22X1 U734 ( .IN1(n779), .IN2(n514), .IN3(n795), .IN4(n516), .Q(n458) );
  OA22X1 U735 ( .IN1(n812), .IN2(n519), .IN3(n832), .IN4(n138), .Q(n457) );
  NAND4X0 U736 ( .IN1(n460), .IN2(n459), .IN3(n458), .IN4(n457), .QN(N270) );
  OA22X1 U737 ( .IN1(n795), .IN2(n508), .IN3(n803), .IN4(n506), .Q(n464) );
  OA22X1 U738 ( .IN1(n763), .IN2(n510), .IN3(n779), .IN4(n512), .Q(n463) );
  OA22X1 U739 ( .IN1(n787), .IN2(n516), .IN3(n771), .IN4(n514), .Q(n462) );
  OA22X1 U740 ( .IN1(n802), .IN2(n519), .IN3(n812), .IN4(n138), .Q(n461) );
  NAND4X0 U741 ( .IN1(n464), .IN2(n463), .IN3(n462), .IN4(n461), .QN(N271) );
  OA22X1 U742 ( .IN1(n787), .IN2(n508), .IN3(n795), .IN4(n506), .Q(n469) );
  OA22X1 U743 ( .IN1(n755), .IN2(n510), .IN3(n771), .IN4(n512), .Q(n468) );
  OA22X1 U744 ( .IN1(n763), .IN2(n514), .IN3(n779), .IN4(n516), .Q(n467) );
  OA22X1 U745 ( .IN1(n803), .IN2(n519), .IN3(n802), .IN4(n138), .Q(n466) );
  NAND4X0 U746 ( .IN1(n469), .IN2(n468), .IN3(n467), .IN4(n466), .QN(N272) );
  OA22X1 U747 ( .IN1(n787), .IN2(n506), .IN3(n779), .IN4(n508), .Q(n474) );
  OA22X1 U748 ( .IN1(n763), .IN2(n512), .IN3(n744), .IN4(n510), .Q(n473) );
  OA22X1 U749 ( .IN1(n755), .IN2(n514), .IN3(n771), .IN4(n516), .Q(n472) );
  OA22X1 U750 ( .IN1(n795), .IN2(n519), .IN3(n803), .IN4(n138), .Q(n471) );
  NAND4X0 U751 ( .IN1(n474), .IN2(n473), .IN3(n472), .IN4(n471), .QN(N273) );
  OA22X1 U752 ( .IN1(n771), .IN2(n508), .IN3(n779), .IN4(n506), .Q(n478) );
  INVX0 U753 ( .INP(n524), .ZN(n518) );
  OA22X1 U754 ( .IN1(n518), .IN2(n510), .IN3(n755), .IN4(n512), .Q(n477) );
  OA22X1 U755 ( .IN1(n763), .IN2(n516), .IN3(n744), .IN4(n514), .Q(n476) );
  OA22X1 U756 ( .IN1(n787), .IN2(n519), .IN3(n795), .IN4(n138), .Q(n475) );
  NAND4X0 U757 ( .IN1(n478), .IN2(n477), .IN3(n476), .IN4(n475), .QN(N274) );
  OA22X1 U758 ( .IN1(n763), .IN2(n508), .IN3(n771), .IN4(n506), .Q(n483) );
  OA22X1 U759 ( .IN1(n590), .IN2(n510), .IN3(n744), .IN4(n512), .Q(n482) );
  OA22X1 U760 ( .IN1(n518), .IN2(n514), .IN3(n755), .IN4(n516), .Q(n481) );
  OA22X1 U761 ( .IN1(n787), .IN2(n138), .IN3(n779), .IN4(n519), .Q(n480) );
  NAND4X0 U762 ( .IN1(n483), .IN2(n482), .IN3(n481), .IN4(n480), .QN(N275) );
  OA22X1 U763 ( .IN1(n755), .IN2(n508), .IN3(n763), .IN4(n506), .Q(n487) );
  OA22X1 U764 ( .IN1(n518), .IN2(n512), .IN3(n507), .IN4(n510), .Q(n486) );
  OA22X1 U765 ( .IN1(n590), .IN2(n514), .IN3(n744), .IN4(n516), .Q(n485) );
  OA22X1 U766 ( .IN1(n771), .IN2(n519), .IN3(n779), .IN4(n138), .Q(n484) );
  NAND4X0 U767 ( .IN1(n487), .IN2(n486), .IN3(n485), .IN4(n484), .QN(N276) );
  OA22X1 U768 ( .IN1(n755), .IN2(n506), .IN3(n744), .IN4(n508), .Q(n492) );
  INVX0 U769 ( .INP(n488), .ZN(n509) );
  OA22X1 U770 ( .IN1(n590), .IN2(n512), .IN3(n509), .IN4(n510), .Q(n491) );
  OA22X1 U771 ( .IN1(n518), .IN2(n516), .IN3(n507), .IN4(n514), .Q(n490) );
  OA22X1 U772 ( .IN1(n763), .IN2(n519), .IN3(n771), .IN4(n138), .Q(n489) );
  NAND4X0 U773 ( .IN1(n492), .IN2(n491), .IN3(n490), .IN4(n489), .QN(N277) );
  OA22X1 U774 ( .IN1(n518), .IN2(n508), .IN3(n744), .IN4(n506), .Q(n496) );
  OA22X1 U775 ( .IN1(n517), .IN2(n510), .IN3(n507), .IN4(n512), .Q(n495) );
  OA22X1 U776 ( .IN1(n590), .IN2(n516), .IN3(n509), .IN4(n514), .Q(n494) );
  OA22X1 U777 ( .IN1(n755), .IN2(n519), .IN3(n763), .IN4(n138), .Q(n493) );
  NAND4X0 U778 ( .IN1(n496), .IN2(n495), .IN3(n494), .IN4(n493), .QN(N278) );
  OA22X1 U779 ( .IN1(n590), .IN2(n508), .IN3(n518), .IN4(n506), .Q(n501) );
  INVX0 U780 ( .INP(n497), .ZN(n513) );
  OA22X1 U781 ( .IN1(n509), .IN2(n512), .IN3(n513), .IN4(n510), .Q(n500) );
  OA22X1 U782 ( .IN1(n517), .IN2(n514), .IN3(n507), .IN4(n516), .Q(n499) );
  OA22X1 U783 ( .IN1(n755), .IN2(n138), .IN3(n744), .IN4(n519), .Q(n498) );
  NAND4X0 U784 ( .IN1(n501), .IN2(n500), .IN3(n499), .IN4(n498), .QN(N279) );
  OA22X1 U785 ( .IN1(n590), .IN2(n506), .IN3(n507), .IN4(n508), .Q(n505) );
  OA22X1 U786 ( .IN1(n517), .IN2(n512), .IN3(n515), .IN4(n510), .Q(n504) );
  OA22X1 U787 ( .IN1(n509), .IN2(n516), .IN3(n513), .IN4(n514), .Q(n503) );
  OA22X1 U788 ( .IN1(n518), .IN2(n519), .IN3(n744), .IN4(n138), .Q(n502) );
  NAND4X0 U789 ( .IN1(n505), .IN2(n504), .IN3(n503), .IN4(n502), .QN(N280) );
  OA22X1 U790 ( .IN1(n509), .IN2(n508), .IN3(n507), .IN4(n506), .Q(n523) );
  OA22X1 U791 ( .IN1(n513), .IN2(n512), .IN3(n511), .IN4(n510), .Q(n522) );
  OA22X1 U792 ( .IN1(n517), .IN2(n516), .IN3(n515), .IN4(n514), .Q(n521) );
  OA22X1 U793 ( .IN1(n590), .IN2(n519), .IN3(n518), .IN4(n138), .Q(n520) );
  NAND4X0 U794 ( .IN1(n523), .IN2(n522), .IN3(n521), .IN4(n520), .QN(N281) );
  NAND3X0 U795 ( .IN1(n524), .IN2(n537), .IN3(n590), .QN(n743) );
  AO22X1 U796 ( .IN1(n535), .IN2(add_result[12]), .IN3(n533), .IN4(
        sub_result[12]), .Q(n525) );
  INVX0 U797 ( .INP(n743), .ZN(n531) );
  NOR3X0 U798 ( .IN1(n526), .IN2(add_result[14]), .IN3(add_result[15]), .QN(
        n528) );
  NOR3X0 U799 ( .IN1(sub_result[14]), .IN2(sub_result[15]), .IN3(n17), .QN(
        n527) );
  AO22X1 U800 ( .IN1(n528), .IN2(add_result[13]), .IN3(n527), .IN4(
        sub_result[13]), .Q(n529) );
  NOR2X0 U801 ( .IN1(n531), .IN2(n530), .QN(N308) );
  INVX0 U802 ( .INP(add_result[12]), .ZN(n534) );
  INVX0 U803 ( .INP(sub_result[12]), .ZN(n532) );
  AO22X1 U804 ( .IN1(n535), .IN2(n534), .IN3(n533), .IN4(n532), .Q(n536) );
  NAND3X0 U805 ( .IN1(n537), .IN2(n750), .IN3(n536), .QN(n837) );
  NAND4X0 U806 ( .IN1(N308), .IN2(n837), .IN3(n820), .IN4(n811), .QN(n804) );
  NAND4X0 U807 ( .IN1(n820), .IN2(n743), .IN3(n749), .IN4(n804), .QN(N306) );
  NAND4X0 U808 ( .IN1(n811), .IN2(n742), .IN3(n749), .IN4(n804), .QN(N307) );
  AO22X1 U809 ( .IN1(n726), .IN2(exponent_factor_12[0]), .IN3(n848), .IN4(
        exponent_factor_21[0]), .Q(N34) );
  NAND3X0 U810 ( .IN1(n832), .IN2(n547), .IN3(n822), .QN(n560) );
  NAND3X0 U811 ( .IN1(n802), .IN2(n539), .IN3(n823), .QN(n555) );
  NAND3X0 U812 ( .IN1(n795), .IN2(n540), .IN3(n790), .QN(n556) );
  NAND3X0 U813 ( .IN1(n834), .IN2(n828), .IN3(n832), .QN(n538) );
  AND2X1 U814 ( .IN1(n555), .IN2(n557), .Q(n542) );
  NAND4X0 U815 ( .IN1(n544), .IN2(n542), .IN3(n556), .IN4(n558), .QN(n543) );
  NAND4X0 U816 ( .IN1(n560), .IN2(n555), .IN3(n556), .IN4(n543), .QN(N346) );
  NAND3X0 U817 ( .IN1(n542), .IN2(n559), .IN3(n543), .QN(N347) );
  NOR2X0 U818 ( .IN1(n836), .IN2(n558), .QN(N349) );
  AO22X1 U819 ( .IN1(n726), .IN2(exponent_factor_12[1]), .IN3(n848), .IN4(
        exponent_factor_21[1]), .Q(N35) );
  OAI22X1 U820 ( .IN1(n828), .IN2(n558), .IN3(n836), .IN4(n556), .QN(N350) );
  OAI222X1 U821 ( .IN1(n557), .IN2(n836), .IN3(n556), .IN4(n828), .IN5(n558), 
        .IN6(n834), .QN(N351) );
  OA22X1 U822 ( .IN1(n834), .IN2(n556), .IN3(n832), .IN4(n558), .Q(n546) );
  OA22X1 U823 ( .IN1(n828), .IN2(n557), .IN3(n836), .IN4(n555), .Q(n545) );
  OA22X1 U824 ( .IN1(n812), .IN2(n558), .IN3(n832), .IN4(n556), .Q(n550) );
  OA22X1 U825 ( .IN1(n834), .IN2(n557), .IN3(n828), .IN4(n555), .Q(n549) );
  AND2X1 U826 ( .IN1(n547), .IN2(n814), .Q(n561) );
  NAND3X0 U827 ( .IN1(n550), .IN2(n549), .IN3(n548), .QN(N353) );
  OA22X1 U828 ( .IN1(n802), .IN2(n558), .IN3(n812), .IN4(n556), .Q(n554) );
  OA22X1 U829 ( .IN1(n834), .IN2(n555), .IN3(n836), .IN4(n560), .Q(n553) );
  OR2X1 U830 ( .IN1(n557), .IN2(n832), .Q(n551) );
  NAND4X0 U831 ( .IN1(n554), .IN2(n553), .IN3(n552), .IN4(n551), .QN(N354) );
  OA22X1 U832 ( .IN1(n802), .IN2(n556), .IN3(n832), .IN4(n555), .Q(n565) );
  OA22X1 U833 ( .IN1(n803), .IN2(n558), .IN3(n812), .IN4(n557), .Q(n564) );
  OA22X1 U834 ( .IN1(n828), .IN2(n560), .IN3(n836), .IN4(n559), .Q(n563) );
  NAND4X0 U835 ( .IN1(n565), .IN2(n564), .IN3(n563), .IN4(n562), .QN(N355) );
  AO22X1 U836 ( .IN1(n726), .IN2(exponent_factor_12[2]), .IN3(n848), .IN4(
        exponent_factor_21[2]), .Q(N36) );
  AO22X1 U837 ( .IN1(n726), .IN2(exponent_factor_12[3]), .IN3(n848), .IN4(
        exponent_factor_21[3]), .Q(N37) );
  AO22X1 U838 ( .IN1(n726), .IN2(exponent_factor_12[4]), .IN3(n848), .IN4(
        exponent_factor_21[4]), .Q(N38) );
  NAND4X0 U839 ( .IN1(n739), .IN2(n568), .IN3(n567), .IN4(n566), .QN(n573) );
  INVX0 U840 ( .INP(input_factor_01[23]), .ZN(n583) );
  NAND4X0 U841 ( .IN1(n583), .IN2(n571), .IN3(n570), .IN4(n569), .QN(n572) );
  NOR2X0 U842 ( .IN1(n573), .IN2(n572), .QN(n582) );
  NOR4X0 U843 ( .IN1(input_factor_01[7]), .IN2(input_factor_01[6]), .IN3(
        input_factor_01[5]), .IN4(input_factor_01[4]), .QN(n581) );
  NOR4X0 U844 ( .IN1(input_factor_01[3]), .IN2(input_factor_01[2]), .IN3(
        input_factor_01[0]), .IN4(input_factor_01[1]), .QN(n580) );
  NAND4X0 U845 ( .IN1(n727), .IN2(n720), .IN3(n714), .IN4(n708), .QN(n578) );
  NAND4X0 U846 ( .IN1(n574), .IN2(n702), .IN3(n696), .IN4(n690), .QN(n577) );
  NAND4X0 U847 ( .IN1(n684), .IN2(n678), .IN3(n672), .IN4(n666), .QN(n576) );
  NAND4X0 U848 ( .IN1(n660), .IN2(n654), .IN3(n648), .IN4(n644), .QN(n575) );
  NOR4X0 U849 ( .IN1(n578), .IN2(n577), .IN3(n576), .IN4(n575), .QN(n579) );
  OA22X1 U850 ( .IN1(n584), .IN2(n729), .IN3(n728), .IN4(n583), .Q(n599) );
  INVX0 U851 ( .INP(n804), .ZN(n585) );
  OA21X1 U852 ( .IN1(n787), .IN2(n586), .IN3(n585), .Q(n592) );
  NAND3X0 U853 ( .IN1(n587), .IN2(n728), .IN3(n729), .QN(n594) );
  OA21X1 U854 ( .IN1(n590), .IN2(n589), .IN3(n588), .Q(n591) );
  AOI22X1 U855 ( .IN1(n732), .IN2(add_output_exponent_w3[0]), .IN3(n731), 
        .IN4(add_output_exponent_w2[0]), .QN(n598) );
  INVX0 U856 ( .INP(n594), .ZN(n593) );
  AND4X1 U857 ( .IN1(n595), .IN2(n593), .IN3(n592), .IN4(n591), .Q(n733) );
  NAND4X0 U858 ( .IN1(n599), .IN2(n598), .IN3(n597), .IN4(n596), .QN(N380) );
  AOI22X1 U859 ( .IN1(input_factor_02[24]), .IN2(n641), .IN3(n640), .IN4(
        input_factor_01[24]), .QN(n603) );
  AOI22X1 U860 ( .IN1(n732), .IN2(add_output_exponent_w3[1]), .IN3(n731), 
        .IN4(add_output_exponent_w2[1]), .QN(n602) );
  NAND4X0 U861 ( .IN1(n603), .IN2(n602), .IN3(n601), .IN4(n600), .QN(N381) );
  AOI22X1 U862 ( .IN1(input_factor_02[25]), .IN2(n641), .IN3(n640), .IN4(
        input_factor_01[25]), .QN(n607) );
  AOI22X1 U863 ( .IN1(n732), .IN2(add_output_exponent_w3[2]), .IN3(n731), 
        .IN4(add_output_exponent_w2[2]), .QN(n606) );
  NAND4X0 U864 ( .IN1(n607), .IN2(n606), .IN3(n605), .IN4(n604), .QN(N382) );
  AOI22X1 U865 ( .IN1(input_factor_02[26]), .IN2(n641), .IN3(n640), .IN4(
        input_factor_01[26]), .QN(n611) );
  AOI22X1 U866 ( .IN1(n732), .IN2(add_output_exponent_w3[3]), .IN3(n731), 
        .IN4(add_output_exponent_w2[3]), .QN(n610) );
  NAND4X0 U867 ( .IN1(n611), .IN2(n610), .IN3(n609), .IN4(n608), .QN(N383) );
  AOI22X1 U868 ( .IN1(input_factor_02[27]), .IN2(n641), .IN3(n640), .IN4(
        input_factor_01[27]), .QN(n615) );
  AOI22X1 U869 ( .IN1(n732), .IN2(add_output_exponent_w3[4]), .IN3(n731), 
        .IN4(add_output_exponent_w2[4]), .QN(n614) );
  NAND4X0 U870 ( .IN1(n615), .IN2(n614), .IN3(n613), .IN4(n612), .QN(N384) );
  AOI22X1 U871 ( .IN1(input_factor_02[28]), .IN2(n641), .IN3(n640), .IN4(
        input_factor_01[28]), .QN(n619) );
  AOI22X1 U872 ( .IN1(n732), .IN2(add_output_exponent_w3[5]), .IN3(n731), 
        .IN4(add_output_exponent_w2[5]), .QN(n618) );
  NAND4X0 U873 ( .IN1(n619), .IN2(n618), .IN3(n617), .IN4(n616), .QN(N385) );
  AOI22X1 U874 ( .IN1(input_factor_02[29]), .IN2(n641), .IN3(n640), .IN4(
        input_factor_01[29]), .QN(n623) );
  AOI22X1 U875 ( .IN1(n732), .IN2(add_output_exponent_w3[6]), .IN3(n731), 
        .IN4(add_output_exponent_w2[6]), .QN(n622) );
  NAND4X0 U876 ( .IN1(n623), .IN2(n622), .IN3(n621), .IN4(n620), .QN(N386) );
  OA22X1 U877 ( .IN1(n740), .IN2(n729), .IN3(n728), .IN4(n739), .Q(n627) );
  AOI22X1 U878 ( .IN1(n732), .IN2(add_output_exponent_w3[7]), .IN3(n731), 
        .IN4(add_output_exponent_w2[7]), .QN(n626) );
  NAND4X0 U879 ( .IN1(n627), .IN2(n626), .IN3(n625), .IN4(n624), .QN(N387) );
  AO222X1 U880 ( .IN1(input_factor_02[0]), .IN2(n641), .IN3(input_factor_01[0]), .IN4(n640), .IN5(n734), .IN6(pre_sig_res_01[0]), .Q(N388) );
  AOI22X1 U881 ( .IN1(n731), .IN2(pre_sig_res_02[1]), .IN3(n734), .IN4(
        pre_sig_res_01[1]), .QN(n629) );
  AOI22X1 U882 ( .IN1(input_factor_02[1]), .IN2(n641), .IN3(n640), .IN4(
        input_factor_01[1]), .QN(n628) );
  AO22X1 U883 ( .IN1(n726), .IN2(exponent_factor_12[5]), .IN3(n848), .IN4(
        exponent_factor_21[5]), .Q(N39) );
  AOI22X1 U884 ( .IN1(n731), .IN2(pre_sig_res_02[2]), .IN3(n734), .IN4(
        pre_sig_res_01[2]), .QN(n631) );
  AOI22X1 U885 ( .IN1(input_factor_02[2]), .IN2(n641), .IN3(n640), .IN4(
        input_factor_01[2]), .QN(n630) );
  AOI22X1 U886 ( .IN1(n731), .IN2(pre_sig_res_02[3]), .IN3(n734), .IN4(
        pre_sig_res_01[3]), .QN(n633) );
  AOI22X1 U887 ( .IN1(input_factor_02[3]), .IN2(n641), .IN3(n640), .IN4(
        input_factor_01[3]), .QN(n632) );
  AOI22X1 U888 ( .IN1(n731), .IN2(pre_sig_res_02[4]), .IN3(n734), .IN4(
        pre_sig_res_01[4]), .QN(n635) );
  AOI22X1 U889 ( .IN1(input_factor_02[4]), .IN2(n641), .IN3(n640), .IN4(
        input_factor_01[4]), .QN(n634) );
  AOI22X1 U890 ( .IN1(n731), .IN2(pre_sig_res_02[5]), .IN3(n734), .IN4(
        pre_sig_res_01[5]), .QN(n637) );
  AOI22X1 U891 ( .IN1(input_factor_02[5]), .IN2(n641), .IN3(n640), .IN4(
        input_factor_01[5]), .QN(n636) );
  AOI22X1 U892 ( .IN1(n731), .IN2(pre_sig_res_02[6]), .IN3(n734), .IN4(
        pre_sig_res_01[6]), .QN(n639) );
  AOI22X1 U893 ( .IN1(input_factor_02[6]), .IN2(n641), .IN3(n640), .IN4(
        input_factor_01[6]), .QN(n638) );
  AOI22X1 U894 ( .IN1(n731), .IN2(pre_sig_res_02[7]), .IN3(n734), .IN4(
        pre_sig_res_01[7]), .QN(n643) );
  AOI22X1 U895 ( .IN1(input_factor_02[7]), .IN2(n641), .IN3(n640), .IN4(
        input_factor_01[7]), .QN(n642) );
  AOI22X1 U896 ( .IN1(n731), .IN2(pre_sig_res_02[8]), .IN3(n734), .IN4(
        pre_sig_res_01[8]), .QN(n647) );
  OA22X1 U897 ( .IN1(n645), .IN2(n729), .IN3(n728), .IN4(n644), .Q(n646) );
  OA22X1 U898 ( .IN1(n649), .IN2(n729), .IN3(n728), .IN4(n648), .Q(n653) );
  NAND4X0 U899 ( .IN1(n653), .IN2(n652), .IN3(n651), .IN4(n650), .QN(N397) );
  OA22X1 U900 ( .IN1(n655), .IN2(n729), .IN3(n728), .IN4(n654), .Q(n659) );
  NAND4X0 U901 ( .IN1(n659), .IN2(n658), .IN3(n657), .IN4(n656), .QN(N398) );
  OA22X1 U902 ( .IN1(n661), .IN2(n729), .IN3(n728), .IN4(n660), .Q(n665) );
  NAND4X0 U903 ( .IN1(n665), .IN2(n664), .IN3(n663), .IN4(n662), .QN(N399) );
  AO22X1 U904 ( .IN1(n726), .IN2(exponent_factor_12[6]), .IN3(n848), .IN4(
        exponent_factor_21[6]), .Q(N40) );
  OA22X1 U905 ( .IN1(n667), .IN2(n729), .IN3(n728), .IN4(n666), .Q(n671) );
  NAND4X0 U906 ( .IN1(n671), .IN2(n670), .IN3(n669), .IN4(n668), .QN(N400) );
  OA22X1 U907 ( .IN1(n673), .IN2(n729), .IN3(n728), .IN4(n672), .Q(n677) );
  NAND4X0 U908 ( .IN1(n677), .IN2(n676), .IN3(n675), .IN4(n674), .QN(N401) );
  OA22X1 U909 ( .IN1(n679), .IN2(n729), .IN3(n728), .IN4(n678), .Q(n683) );
  NAND4X0 U910 ( .IN1(n683), .IN2(n682), .IN3(n681), .IN4(n680), .QN(N402) );
  OA22X1 U911 ( .IN1(n685), .IN2(n729), .IN3(n728), .IN4(n684), .Q(n689) );
  NAND4X0 U912 ( .IN1(n689), .IN2(n688), .IN3(n687), .IN4(n686), .QN(N403) );
  OA22X1 U913 ( .IN1(n691), .IN2(n729), .IN3(n728), .IN4(n690), .Q(n695) );
  AOI22X1 U914 ( .IN1(n732), .IN2(pre_sig_res_03[16]), .IN3(n731), .IN4(
        pre_sig_res_02[16]), .QN(n694) );
  NAND4X0 U915 ( .IN1(n695), .IN2(n694), .IN3(n693), .IN4(n692), .QN(N404) );
  OA22X1 U916 ( .IN1(n697), .IN2(n729), .IN3(n728), .IN4(n696), .Q(n701) );
  AOI22X1 U917 ( .IN1(n732), .IN2(pre_sig_res_03[17]), .IN3(n731), .IN4(
        pre_sig_res_02[17]), .QN(n700) );
  NAND4X0 U918 ( .IN1(n701), .IN2(n700), .IN3(n699), .IN4(n698), .QN(N405) );
  OA22X1 U919 ( .IN1(n703), .IN2(n729), .IN3(n728), .IN4(n702), .Q(n707) );
  AOI22X1 U920 ( .IN1(n732), .IN2(pre_sig_res_03[18]), .IN3(n731), .IN4(
        pre_sig_res_02[18]), .QN(n706) );
  NAND4X0 U921 ( .IN1(n707), .IN2(n706), .IN3(n705), .IN4(n704), .QN(N406) );
  OA22X1 U922 ( .IN1(n709), .IN2(n729), .IN3(n728), .IN4(n708), .Q(n713) );
  AOI22X1 U923 ( .IN1(n732), .IN2(pre_sig_res_03[19]), .IN3(n731), .IN4(
        pre_sig_res_02[19]), .QN(n712) );
  NAND4X0 U924 ( .IN1(n713), .IN2(n712), .IN3(n711), .IN4(n710), .QN(N407) );
  OA22X1 U925 ( .IN1(n715), .IN2(n729), .IN3(n728), .IN4(n714), .Q(n719) );
  AOI22X1 U926 ( .IN1(n732), .IN2(pre_sig_res_03[20]), .IN3(n731), .IN4(
        pre_sig_res_02[20]), .QN(n718) );
  NAND4X0 U927 ( .IN1(n719), .IN2(n718), .IN3(n717), .IN4(n716), .QN(N408) );
  OA22X1 U928 ( .IN1(n721), .IN2(n729), .IN3(n728), .IN4(n720), .Q(n725) );
  AOI22X1 U929 ( .IN1(n732), .IN2(pre_sig_res_03[21]), .IN3(n731), .IN4(
        pre_sig_res_02[21]), .QN(n724) );
  NAND4X0 U930 ( .IN1(n725), .IN2(n724), .IN3(n723), .IN4(n722), .QN(N409) );
  AO22X1 U931 ( .IN1(n726), .IN2(exponent_factor_12[7]), .IN3(n848), .IN4(
        exponent_factor_21[7]), .Q(N41) );
  OA22X1 U932 ( .IN1(n730), .IN2(n729), .IN3(n728), .IN4(n727), .Q(n738) );
  AOI22X1 U933 ( .IN1(n732), .IN2(pre_sig_res_03[22]), .IN3(n731), .IN4(
        pre_sig_res_02[22]), .QN(n737) );
  NAND4X0 U934 ( .IN1(n738), .IN2(n737), .IN3(n736), .IN4(n735), .QN(N410) );
  AO22X1 U935 ( .IN1(larger_exponent[7]), .IN2(n78), .IN3(rst_n), .IN4(n741), 
        .Q(n115) );
  NOR2X0 U936 ( .IN1(n78), .IN2(n742), .QN(n843) );
  NOR2X0 U937 ( .IN1(n743), .IN2(n78), .QN(n845) );
  OA22X1 U938 ( .IN1(n755), .IN2(n833), .IN3(n744), .IN4(n831), .Q(n754) );
  OA22X1 U939 ( .IN1(n771), .IN2(n837), .IN3(n795), .IN4(n804), .Q(n748) );
  INVX0 U940 ( .INP(rst_n), .ZN(n846) );
  NAND3X0 U941 ( .IN1(n746), .IN2(n766), .IN3(n745), .QN(n747) );
  OA22X1 U942 ( .IN1(n78), .IN2(n748), .IN3(n846), .IN4(n747), .Q(n753) );
  NAND4X0 U943 ( .IN1(n754), .IN2(n753), .IN3(n752), .IN4(n751), .QN(n94) );
  OA22X1 U944 ( .IN1(n755), .IN2(n831), .IN3(n763), .IN4(n833), .Q(n762) );
  OA22X1 U945 ( .IN1(n795), .IN2(n811), .IN3(n803), .IN4(n804), .Q(n757) );
  OA22X1 U946 ( .IN1(n787), .IN2(n820), .IN3(n779), .IN4(n837), .Q(n756) );
  AO21X1 U947 ( .IN1(n757), .IN2(n756), .IN3(n78), .Q(n761) );
  NAND4X0 U948 ( .IN1(n762), .IN2(n761), .IN3(n760), .IN4(n759), .QN(n95) );
  OA22X1 U949 ( .IN1(n763), .IN2(n831), .IN3(n771), .IN4(n833), .Q(n770) );
  OA22X1 U950 ( .IN1(n803), .IN2(n811), .IN3(n802), .IN4(n804), .Q(n765) );
  OA22X1 U951 ( .IN1(n787), .IN2(n837), .IN3(n795), .IN4(n820), .Q(n764) );
  AO21X1 U952 ( .IN1(n765), .IN2(n764), .IN3(n78), .Q(n769) );
  NAND4X0 U953 ( .IN1(n770), .IN2(n769), .IN3(n768), .IN4(n767), .QN(n96) );
  OA22X1 U954 ( .IN1(n771), .IN2(n831), .IN3(n779), .IN4(n833), .Q(n778) );
  OA22X1 U955 ( .IN1(n802), .IN2(n811), .IN3(n812), .IN4(n804), .Q(n773) );
  OA22X1 U956 ( .IN1(n795), .IN2(n837), .IN3(n803), .IN4(n820), .Q(n772) );
  AO21X1 U957 ( .IN1(n773), .IN2(n772), .IN3(n78), .Q(n777) );
  NAND4X0 U958 ( .IN1(n778), .IN2(n777), .IN3(n776), .IN4(n775), .QN(n97) );
  OA22X1 U959 ( .IN1(n787), .IN2(n833), .IN3(n779), .IN4(n831), .Q(n786) );
  OA22X1 U960 ( .IN1(n812), .IN2(n811), .IN3(n832), .IN4(n804), .Q(n781) );
  OA22X1 U961 ( .IN1(n803), .IN2(n837), .IN3(n802), .IN4(n820), .Q(n780) );
  AO21X1 U962 ( .IN1(n781), .IN2(n780), .IN3(n78), .Q(n785) );
  NAND4X0 U963 ( .IN1(n786), .IN2(n785), .IN3(n784), .IN4(n783), .QN(n98) );
  OA22X1 U964 ( .IN1(n787), .IN2(n831), .IN3(n795), .IN4(n833), .Q(n794) );
  OA22X1 U965 ( .IN1(n834), .IN2(n804), .IN3(n832), .IN4(n811), .Q(n789) );
  OA22X1 U966 ( .IN1(n802), .IN2(n837), .IN3(n812), .IN4(n820), .Q(n788) );
  AO21X1 U967 ( .IN1(n789), .IN2(n788), .IN3(n78), .Q(n793) );
  NAND4X0 U968 ( .IN1(n794), .IN2(n793), .IN3(n792), .IN4(n791), .QN(n99) );
  OA22X1 U969 ( .IN1(n795), .IN2(n831), .IN3(n803), .IN4(n833), .Q(n801) );
  OA22X1 U970 ( .IN1(n834), .IN2(n811), .IN3(n828), .IN4(n804), .Q(n797) );
  OA22X1 U971 ( .IN1(n812), .IN2(n837), .IN3(n832), .IN4(n820), .Q(n796) );
  AO21X1 U972 ( .IN1(n797), .IN2(n796), .IN3(n78), .Q(n800) );
  NAND4X0 U973 ( .IN1(n801), .IN2(n800), .IN3(n799), .IN4(n798), .QN(n100) );
  OA22X1 U974 ( .IN1(n803), .IN2(n831), .IN3(n802), .IN4(n833), .Q(n810) );
  OA22X1 U975 ( .IN1(n828), .IN2(n811), .IN3(n836), .IN4(n804), .Q(n806) );
  OA22X1 U976 ( .IN1(n834), .IN2(n820), .IN3(n832), .IN4(n837), .Q(n805) );
  AO21X1 U977 ( .IN1(n806), .IN2(n805), .IN3(n78), .Q(n809) );
  NAND4X0 U978 ( .IN1(n810), .IN2(n809), .IN3(n808), .IN4(n807), .QN(n101) );
  OA222X1 U979 ( .IN1(n837), .IN2(n834), .IN3(n811), .IN4(n836), .IN5(n820), 
        .IN6(n828), .Q(n813) );
  OA22X1 U980 ( .IN1(n78), .IN2(n813), .IN3(n812), .IN4(n833), .Q(n819) );
  NAND4X0 U981 ( .IN1(n819), .IN2(n818), .IN3(n817), .IN4(n816), .QN(n102) );
  OA22X1 U982 ( .IN1(n828), .IN2(n837), .IN3(n836), .IN4(n820), .Q(n821) );
  OA22X1 U983 ( .IN1(n832), .IN2(n833), .IN3(n821), .IN4(n846), .Q(n827) );
  NAND4X0 U984 ( .IN1(n827), .IN2(n826), .IN3(n825), .IN4(n824), .QN(n103) );
  AOI22X1 U985 ( .IN1(pre_sig_res_03[11]), .IN2(n846), .IN3(n835), .IN4(n844), 
        .QN(n830) );
  OA22X1 U986 ( .IN1(n834), .IN2(n831), .IN3(n828), .IN4(n833), .Q(n829) );
  OA22X1 U987 ( .IN1(n834), .IN2(n833), .IN3(n832), .IN4(n831), .Q(n841) );
  OR3X1 U988 ( .IN1(n837), .IN2(n846), .IN3(n836), .Q(n839) );
  NAND4X0 U989 ( .IN1(n841), .IN2(n840), .IN3(n839), .IN4(n838), .QN(n105) );
  AO222X1 U990 ( .IN1(n844), .IN2(n843), .IN3(n842), .IN4(n845), .IN5(n846), 
        .IN6(pre_sig_res_03[10]), .Q(n106) );
  AO22X1 U991 ( .IN1(pre_sig_res_03[9]), .IN2(n846), .IN3(n845), .IN4(n844), 
        .Q(n107) );
  AO222X1 U992 ( .IN1(input_factor_02[23]), .IN2(n850), .IN3(
        input_factor_01[23]), .IN4(n849), .IN5(larger_exponent[0]), .IN6(n78), 
        .Q(n108) );
  AO222X1 U993 ( .IN1(input_factor_02[24]), .IN2(n850), .IN3(
        input_factor_01[24]), .IN4(n849), .IN5(n78), .IN6(larger_exponent[1]), 
        .Q(n109) );
  AO222X1 U994 ( .IN1(input_factor_02[25]), .IN2(n850), .IN3(
        input_factor_01[25]), .IN4(n849), .IN5(n78), .IN6(larger_exponent[2]), 
        .Q(n110) );
  AO222X1 U995 ( .IN1(input_factor_02[26]), .IN2(n850), .IN3(
        input_factor_01[26]), .IN4(n849), .IN5(n78), .IN6(larger_exponent[3]), 
        .Q(n111) );
  AO222X1 U996 ( .IN1(input_factor_02[27]), .IN2(n850), .IN3(
        input_factor_01[27]), .IN4(n849), .IN5(n78), .IN6(larger_exponent[4]), 
        .Q(n112) );
  AO222X1 U997 ( .IN1(input_factor_02[28]), .IN2(n850), .IN3(
        input_factor_01[28]), .IN4(n849), .IN5(n78), .IN6(larger_exponent[5]), 
        .Q(n113) );
  AO222X1 U998 ( .IN1(input_factor_02[29]), .IN2(n850), .IN3(
        input_factor_01[29]), .IN4(n849), .IN5(n78), .IN6(larger_exponent[6]), 
        .Q(n114) );
endmodule


module mac ( clk, rst_n, refresh_mac, ena_mac, ena_mac_wait, ena_mul_add, 
        mac_input_01, mac_input_02, mac_output );
  input [31:0] mac_input_01;
  input [31:0] mac_input_02;
  output [31:0] mac_output;
  input clk, rst_n, refresh_mac, ena_mac, ena_mac_wait, ena_mul_add;
  wire   n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n138;
  wire   [31:0] next_mac_input_01;
  wire   [31:0] next_mac_input_02;
  wire   [31:0] weight_input_mul;
  wire   [31:0] next_weight_input_mul;
  wire   [31:0] pre_adder_output;

  floating_point_multiple_0 floating_point_multiple_01 ( .clk(clk), .rst_n(
        rst_n), .input_factor_01(next_mac_input_01), .input_factor_02(
        next_mac_input_02), .output_multiply(weight_input_mul) );
  floating_point_adder_0 floating_point_adder_01 ( .clk(clk), .rst_n(rst_n), 
        .input_factor_01(next_weight_input_mul), .input_factor_02(mac_output), 
        .output_adder(pre_adder_output) );
  DFFARX1 next_mac_input_01_reg_31_ ( .D(n137), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_01[31]) );
  DFFARX1 next_mac_input_01_reg_30_ ( .D(n136), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_01[30]) );
  DFFARX1 next_mac_input_01_reg_29_ ( .D(n135), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_01[29]) );
  DFFARX1 next_mac_input_01_reg_28_ ( .D(n134), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_01[28]) );
  DFFARX1 next_mac_input_01_reg_27_ ( .D(n133), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_01[27]) );
  DFFARX1 next_mac_input_01_reg_26_ ( .D(n132), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_01[26]) );
  DFFARX1 next_mac_input_01_reg_25_ ( .D(n131), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_01[25]) );
  DFFARX1 next_mac_input_01_reg_24_ ( .D(n130), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_01[24]) );
  DFFARX1 next_mac_input_01_reg_23_ ( .D(n129), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_01[23]) );
  DFFARX1 next_mac_input_01_reg_22_ ( .D(n128), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_01[22]) );
  DFFARX1 next_mac_input_01_reg_21_ ( .D(n127), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_01[21]) );
  DFFARX1 next_mac_input_01_reg_20_ ( .D(n126), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_01[20]) );
  DFFARX1 next_mac_input_01_reg_19_ ( .D(n125), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_01[19]) );
  DFFARX1 next_mac_input_01_reg_18_ ( .D(n124), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_01[18]) );
  DFFARX1 next_mac_input_01_reg_17_ ( .D(n123), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_01[17]) );
  DFFARX1 next_mac_input_01_reg_16_ ( .D(n122), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_01[16]) );
  DFFARX1 next_mac_input_01_reg_15_ ( .D(n121), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_01[15]) );
  DFFARX1 next_mac_input_01_reg_14_ ( .D(n120), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_01[14]) );
  DFFARX1 next_mac_input_01_reg_13_ ( .D(n119), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_01[13]) );
  DFFARX1 next_mac_input_01_reg_12_ ( .D(n118), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_01[12]) );
  DFFARX1 next_mac_input_01_reg_11_ ( .D(n117), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_01[11]) );
  DFFARX1 next_mac_input_01_reg_10_ ( .D(n116), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_01[10]) );
  DFFARX1 next_mac_input_01_reg_9_ ( .D(n115), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_01[9]) );
  DFFARX1 next_mac_input_01_reg_8_ ( .D(n114), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_01[8]) );
  DFFARX1 next_mac_input_01_reg_7_ ( .D(n113), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_01[7]) );
  DFFARX1 next_mac_input_01_reg_6_ ( .D(n112), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_01[6]) );
  DFFARX1 next_mac_input_01_reg_5_ ( .D(n111), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_01[5]) );
  DFFARX1 next_mac_input_01_reg_4_ ( .D(n110), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_01[4]) );
  DFFARX1 next_mac_input_01_reg_3_ ( .D(n109), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_01[3]) );
  DFFARX1 next_mac_input_01_reg_2_ ( .D(n108), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_01[2]) );
  DFFARX1 next_mac_input_01_reg_1_ ( .D(n107), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_01[1]) );
  DFFARX1 next_mac_input_01_reg_0_ ( .D(n106), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_01[0]) );
  DFFARX1 next_mac_input_02_reg_31_ ( .D(n105), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_02[31]) );
  DFFARX1 next_mac_input_02_reg_30_ ( .D(n104), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_02[30]) );
  DFFARX1 next_mac_input_02_reg_29_ ( .D(n103), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_02[29]) );
  DFFARX1 next_mac_input_02_reg_28_ ( .D(n102), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_02[28]) );
  DFFARX1 next_mac_input_02_reg_27_ ( .D(n101), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_02[27]) );
  DFFARX1 next_mac_input_02_reg_26_ ( .D(n100), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_02[26]) );
  DFFARX1 next_mac_input_02_reg_25_ ( .D(n99), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_02[25]) );
  DFFARX1 next_mac_input_02_reg_24_ ( .D(n98), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_02[24]) );
  DFFARX1 next_mac_input_02_reg_23_ ( .D(n97), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_02[23]) );
  DFFARX1 next_mac_input_02_reg_22_ ( .D(n96), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_02[22]) );
  DFFARX1 next_mac_input_02_reg_21_ ( .D(n95), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_02[21]) );
  DFFARX1 next_mac_input_02_reg_20_ ( .D(n94), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_02[20]) );
  DFFARX1 next_mac_input_02_reg_19_ ( .D(n93), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_02[19]) );
  DFFARX1 next_mac_input_02_reg_18_ ( .D(n92), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_02[18]) );
  DFFARX1 next_mac_input_02_reg_17_ ( .D(n91), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_02[17]) );
  DFFARX1 next_mac_input_02_reg_16_ ( .D(n90), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_02[16]) );
  DFFARX1 next_mac_input_02_reg_15_ ( .D(n89), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_02[15]) );
  DFFARX1 next_mac_input_02_reg_14_ ( .D(n88), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_02[14]) );
  DFFARX1 next_mac_input_02_reg_13_ ( .D(n87), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_02[13]) );
  DFFARX1 next_mac_input_02_reg_12_ ( .D(n86), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_02[12]) );
  DFFARX1 next_mac_input_02_reg_11_ ( .D(n85), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_02[11]) );
  DFFARX1 next_mac_input_02_reg_10_ ( .D(n84), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_02[10]) );
  DFFARX1 next_mac_input_02_reg_9_ ( .D(n83), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_02[9]) );
  DFFARX1 next_mac_input_02_reg_8_ ( .D(n82), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_02[8]) );
  DFFARX1 next_mac_input_02_reg_7_ ( .D(n81), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_02[7]) );
  DFFARX1 next_mac_input_02_reg_6_ ( .D(n80), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_02[6]) );
  DFFARX1 next_mac_input_02_reg_5_ ( .D(n79), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_02[5]) );
  DFFARX1 next_mac_input_02_reg_4_ ( .D(n78), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_02[4]) );
  DFFARX1 next_mac_input_02_reg_3_ ( .D(n77), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_02[3]) );
  DFFARX1 next_mac_input_02_reg_2_ ( .D(n76), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_02[2]) );
  DFFARX1 next_mac_input_02_reg_1_ ( .D(n75), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_02[1]) );
  DFFARX1 next_mac_input_02_reg_0_ ( .D(n74), .CLK(clk), .RSTB(rst_n), .Q(
        next_mac_input_02[0]) );
  DFFARX1 next_weight_input_mul_reg_31_ ( .D(n73), .CLK(clk), .RSTB(rst_n), 
        .Q(next_weight_input_mul[31]) );
  DFFARX1 next_weight_input_mul_reg_30_ ( .D(n72), .CLK(clk), .RSTB(rst_n), 
        .Q(next_weight_input_mul[30]) );
  DFFARX1 next_weight_input_mul_reg_29_ ( .D(n71), .CLK(clk), .RSTB(rst_n), 
        .Q(next_weight_input_mul[29]) );
  DFFARX1 next_weight_input_mul_reg_28_ ( .D(n70), .CLK(clk), .RSTB(rst_n), 
        .Q(next_weight_input_mul[28]) );
  DFFARX1 next_weight_input_mul_reg_27_ ( .D(n69), .CLK(clk), .RSTB(rst_n), 
        .Q(next_weight_input_mul[27]) );
  DFFARX1 next_weight_input_mul_reg_26_ ( .D(n68), .CLK(clk), .RSTB(rst_n), 
        .Q(next_weight_input_mul[26]) );
  DFFARX1 next_weight_input_mul_reg_25_ ( .D(n67), .CLK(clk), .RSTB(rst_n), 
        .Q(next_weight_input_mul[25]) );
  DFFARX1 next_weight_input_mul_reg_24_ ( .D(n66), .CLK(clk), .RSTB(rst_n), 
        .Q(next_weight_input_mul[24]) );
  DFFARX1 next_weight_input_mul_reg_23_ ( .D(n65), .CLK(clk), .RSTB(rst_n), 
        .Q(next_weight_input_mul[23]) );
  DFFARX1 next_weight_input_mul_reg_22_ ( .D(n64), .CLK(clk), .RSTB(rst_n), 
        .Q(next_weight_input_mul[22]) );
  DFFARX1 next_weight_input_mul_reg_21_ ( .D(n63), .CLK(clk), .RSTB(rst_n), 
        .Q(next_weight_input_mul[21]) );
  DFFARX1 next_weight_input_mul_reg_20_ ( .D(n62), .CLK(clk), .RSTB(rst_n), 
        .Q(next_weight_input_mul[20]) );
  DFFARX1 next_weight_input_mul_reg_19_ ( .D(n61), .CLK(clk), .RSTB(rst_n), 
        .Q(next_weight_input_mul[19]) );
  DFFARX1 next_weight_input_mul_reg_18_ ( .D(n60), .CLK(clk), .RSTB(rst_n), 
        .Q(next_weight_input_mul[18]) );
  DFFARX1 next_weight_input_mul_reg_17_ ( .D(n59), .CLK(clk), .RSTB(rst_n), 
        .Q(next_weight_input_mul[17]) );
  DFFARX1 next_weight_input_mul_reg_16_ ( .D(n58), .CLK(clk), .RSTB(rst_n), 
        .Q(next_weight_input_mul[16]) );
  DFFARX1 next_weight_input_mul_reg_15_ ( .D(n57), .CLK(clk), .RSTB(rst_n), 
        .Q(next_weight_input_mul[15]) );
  DFFARX1 next_weight_input_mul_reg_14_ ( .D(n56), .CLK(clk), .RSTB(rst_n), 
        .Q(next_weight_input_mul[14]) );
  DFFARX1 next_weight_input_mul_reg_13_ ( .D(n55), .CLK(clk), .RSTB(rst_n), 
        .Q(next_weight_input_mul[13]) );
  DFFARX1 next_weight_input_mul_reg_12_ ( .D(n54), .CLK(clk), .RSTB(rst_n), 
        .Q(next_weight_input_mul[12]) );
  DFFARX1 next_weight_input_mul_reg_11_ ( .D(n53), .CLK(clk), .RSTB(rst_n), 
        .Q(next_weight_input_mul[11]) );
  DFFARX1 next_weight_input_mul_reg_10_ ( .D(n52), .CLK(clk), .RSTB(rst_n), 
        .Q(next_weight_input_mul[10]) );
  DFFARX1 next_weight_input_mul_reg_9_ ( .D(n51), .CLK(clk), .RSTB(rst_n), .Q(
        next_weight_input_mul[9]) );
  DFFARX1 next_weight_input_mul_reg_8_ ( .D(n50), .CLK(clk), .RSTB(rst_n), .Q(
        next_weight_input_mul[8]) );
  DFFARX1 next_weight_input_mul_reg_7_ ( .D(n49), .CLK(clk), .RSTB(rst_n), .Q(
        next_weight_input_mul[7]) );
  DFFARX1 next_weight_input_mul_reg_6_ ( .D(n48), .CLK(clk), .RSTB(rst_n), .Q(
        next_weight_input_mul[6]) );
  DFFARX1 next_weight_input_mul_reg_5_ ( .D(n47), .CLK(clk), .RSTB(rst_n), .Q(
        next_weight_input_mul[5]) );
  DFFARX1 next_weight_input_mul_reg_4_ ( .D(n46), .CLK(clk), .RSTB(rst_n), .Q(
        next_weight_input_mul[4]) );
  DFFARX1 next_weight_input_mul_reg_3_ ( .D(n45), .CLK(clk), .RSTB(rst_n), .Q(
        next_weight_input_mul[3]) );
  DFFARX1 next_weight_input_mul_reg_2_ ( .D(n44), .CLK(clk), .RSTB(rst_n), .Q(
        next_weight_input_mul[2]) );
  DFFARX1 next_weight_input_mul_reg_1_ ( .D(n43), .CLK(clk), .RSTB(rst_n), .Q(
        next_weight_input_mul[1]) );
  DFFARX1 next_weight_input_mul_reg_0_ ( .D(n42), .CLK(clk), .RSTB(rst_n), .Q(
        next_weight_input_mul[0]) );
  DFFARX1 next_adder_output_reg_0_ ( .D(n41), .CLK(clk), .RSTB(rst_n), .Q(
        mac_output[0]) );
  DFFARX1 next_adder_output_reg_1_ ( .D(n40), .CLK(clk), .RSTB(rst_n), .Q(
        mac_output[1]) );
  DFFARX1 next_adder_output_reg_2_ ( .D(n39), .CLK(clk), .RSTB(rst_n), .Q(
        mac_output[2]) );
  DFFARX1 next_adder_output_reg_3_ ( .D(n38), .CLK(clk), .RSTB(rst_n), .Q(
        mac_output[3]) );
  DFFARX1 next_adder_output_reg_4_ ( .D(n37), .CLK(clk), .RSTB(rst_n), .Q(
        mac_output[4]) );
  DFFARX1 next_adder_output_reg_5_ ( .D(n36), .CLK(clk), .RSTB(rst_n), .Q(
        mac_output[5]) );
  DFFARX1 next_adder_output_reg_6_ ( .D(n35), .CLK(clk), .RSTB(rst_n), .Q(
        mac_output[6]) );
  DFFARX1 next_adder_output_reg_7_ ( .D(n34), .CLK(clk), .RSTB(rst_n), .Q(
        mac_output[7]) );
  DFFARX1 next_adder_output_reg_8_ ( .D(n33), .CLK(clk), .RSTB(rst_n), .Q(
        mac_output[8]) );
  DFFARX1 next_adder_output_reg_9_ ( .D(n32), .CLK(clk), .RSTB(rst_n), .Q(
        mac_output[9]) );
  DFFARX1 next_adder_output_reg_10_ ( .D(n31), .CLK(clk), .RSTB(rst_n), .Q(
        mac_output[10]) );
  DFFARX1 next_adder_output_reg_11_ ( .D(n30), .CLK(clk), .RSTB(rst_n), .Q(
        mac_output[11]) );
  DFFARX1 next_adder_output_reg_12_ ( .D(n29), .CLK(clk), .RSTB(rst_n), .Q(
        mac_output[12]) );
  DFFARX1 next_adder_output_reg_13_ ( .D(n28), .CLK(clk), .RSTB(rst_n), .Q(
        mac_output[13]) );
  DFFARX1 next_adder_output_reg_14_ ( .D(n27), .CLK(clk), .RSTB(rst_n), .Q(
        mac_output[14]) );
  DFFARX1 next_adder_output_reg_15_ ( .D(n26), .CLK(clk), .RSTB(rst_n), .Q(
        mac_output[15]) );
  DFFARX1 next_adder_output_reg_16_ ( .D(n25), .CLK(clk), .RSTB(rst_n), .Q(
        mac_output[16]) );
  DFFARX1 next_adder_output_reg_17_ ( .D(n24), .CLK(clk), .RSTB(rst_n), .Q(
        mac_output[17]) );
  DFFARX1 next_adder_output_reg_18_ ( .D(n23), .CLK(clk), .RSTB(rst_n), .Q(
        mac_output[18]) );
  DFFARX1 next_adder_output_reg_19_ ( .D(n22), .CLK(clk), .RSTB(rst_n), .Q(
        mac_output[19]) );
  DFFARX1 next_adder_output_reg_20_ ( .D(n21), .CLK(clk), .RSTB(rst_n), .Q(
        mac_output[20]) );
  DFFARX1 next_adder_output_reg_21_ ( .D(n20), .CLK(clk), .RSTB(rst_n), .Q(
        mac_output[21]) );
  DFFARX1 next_adder_output_reg_22_ ( .D(n19), .CLK(clk), .RSTB(rst_n), .Q(
        mac_output[22]) );
  DFFARX1 next_adder_output_reg_23_ ( .D(n18), .CLK(clk), .RSTB(rst_n), .Q(
        mac_output[23]) );
  DFFARX1 next_adder_output_reg_24_ ( .D(n17), .CLK(clk), .RSTB(rst_n), .Q(
        mac_output[24]) );
  DFFARX1 next_adder_output_reg_25_ ( .D(n16), .CLK(clk), .RSTB(rst_n), .Q(
        mac_output[25]) );
  DFFARX1 next_adder_output_reg_26_ ( .D(n15), .CLK(clk), .RSTB(rst_n), .Q(
        mac_output[26]) );
  DFFARX1 next_adder_output_reg_27_ ( .D(n14), .CLK(clk), .RSTB(rst_n), .Q(
        mac_output[27]) );
  DFFARX1 next_adder_output_reg_28_ ( .D(n13), .CLK(clk), .RSTB(rst_n), .Q(
        mac_output[28]) );
  DFFARX1 next_adder_output_reg_29_ ( .D(n12), .CLK(clk), .RSTB(rst_n), .Q(
        mac_output[29]) );
  DFFARX1 next_adder_output_reg_30_ ( .D(n11), .CLK(clk), .RSTB(rst_n), .Q(
        mac_output[30]) );
  DFFARX1 next_adder_output_reg_31_ ( .D(n10), .CLK(clk), .RSTB(rst_n), .Q(
        mac_output[31]) );
  NOR2X0 U2 ( .IN1(n8), .IN2(ena_mul_add), .QN(n2) );
  INVX0 U3 ( .INP(n4), .ZN(n3) );
  NOR2X0 U4 ( .IN1(ena_mul_add), .IN2(n5), .QN(n6) );
  INVX0 U5 ( .INP(ena_mac), .ZN(n5) );
  AND2X1 U6 ( .IN1(ena_mac), .IN2(ena_mul_add), .Q(n7) );
  NOR2X0 U7 ( .IN1(refresh_mac), .IN2(n138), .QN(n1) );
  NOR2X0 U8 ( .IN1(refresh_mac), .IN2(n9), .QN(n138) );
  OA21X1 U9 ( .IN1(ena_mac_wait), .IN2(ena_mac), .IN3(ena_mul_add), .Q(n9) );
  NOR2X0 U10 ( .IN1(ena_mac_wait), .IN2(ena_mac), .QN(n8) );
  INVX0 U11 ( .INP(n6), .ZN(n4) );
  AO22X1 U12 ( .IN1(n7), .IN2(mac_input_01[31]), .IN3(n3), .IN4(
        next_mac_input_01[31]), .Q(n137) );
  AO22X1 U13 ( .IN1(n7), .IN2(mac_input_01[30]), .IN3(n3), .IN4(
        next_mac_input_01[30]), .Q(n136) );
  AO22X1 U14 ( .IN1(n7), .IN2(mac_input_01[29]), .IN3(n3), .IN4(
        next_mac_input_01[29]), .Q(n135) );
  AO22X1 U15 ( .IN1(n7), .IN2(mac_input_01[28]), .IN3(n3), .IN4(
        next_mac_input_01[28]), .Q(n134) );
  AO22X1 U16 ( .IN1(n7), .IN2(mac_input_01[27]), .IN3(n3), .IN4(
        next_mac_input_01[27]), .Q(n133) );
  AO22X1 U17 ( .IN1(n7), .IN2(mac_input_01[26]), .IN3(n3), .IN4(
        next_mac_input_01[26]), .Q(n132) );
  AO22X1 U18 ( .IN1(n7), .IN2(mac_input_01[25]), .IN3(n3), .IN4(
        next_mac_input_01[25]), .Q(n131) );
  AO22X1 U19 ( .IN1(n7), .IN2(mac_input_01[24]), .IN3(n3), .IN4(
        next_mac_input_01[24]), .Q(n130) );
  AO22X1 U20 ( .IN1(n7), .IN2(mac_input_01[23]), .IN3(n3), .IN4(
        next_mac_input_01[23]), .Q(n129) );
  AO22X1 U21 ( .IN1(n7), .IN2(mac_input_01[22]), .IN3(n3), .IN4(
        next_mac_input_01[22]), .Q(n128) );
  AO22X1 U22 ( .IN1(n7), .IN2(mac_input_01[21]), .IN3(n3), .IN4(
        next_mac_input_01[21]), .Q(n127) );
  AO22X1 U23 ( .IN1(n7), .IN2(mac_input_01[20]), .IN3(n3), .IN4(
        next_mac_input_01[20]), .Q(n126) );
  AO22X1 U24 ( .IN1(n7), .IN2(mac_input_01[19]), .IN3(n6), .IN4(
        next_mac_input_01[19]), .Q(n125) );
  AO22X1 U25 ( .IN1(n7), .IN2(mac_input_01[18]), .IN3(n6), .IN4(
        next_mac_input_01[18]), .Q(n124) );
  AO22X1 U26 ( .IN1(n7), .IN2(mac_input_01[17]), .IN3(n6), .IN4(
        next_mac_input_01[17]), .Q(n123) );
  AO22X1 U27 ( .IN1(n7), .IN2(mac_input_01[16]), .IN3(n6), .IN4(
        next_mac_input_01[16]), .Q(n122) );
  AO22X1 U28 ( .IN1(n7), .IN2(mac_input_01[15]), .IN3(n6), .IN4(
        next_mac_input_01[15]), .Q(n121) );
  AO22X1 U29 ( .IN1(n7), .IN2(mac_input_01[14]), .IN3(n6), .IN4(
        next_mac_input_01[14]), .Q(n120) );
  AO22X1 U30 ( .IN1(n7), .IN2(mac_input_01[13]), .IN3(n6), .IN4(
        next_mac_input_01[13]), .Q(n119) );
  AO22X1 U31 ( .IN1(n7), .IN2(mac_input_01[12]), .IN3(n6), .IN4(
        next_mac_input_01[12]), .Q(n118) );
  AO22X1 U32 ( .IN1(n7), .IN2(mac_input_01[11]), .IN3(n3), .IN4(
        next_mac_input_01[11]), .Q(n117) );
  AO22X1 U33 ( .IN1(n7), .IN2(mac_input_01[10]), .IN3(n6), .IN4(
        next_mac_input_01[10]), .Q(n116) );
  AO22X1 U34 ( .IN1(n7), .IN2(mac_input_01[9]), .IN3(n3), .IN4(
        next_mac_input_01[9]), .Q(n115) );
  AO22X1 U35 ( .IN1(n7), .IN2(mac_input_01[8]), .IN3(n3), .IN4(
        next_mac_input_01[8]), .Q(n114) );
  AO22X1 U36 ( .IN1(n7), .IN2(mac_input_01[7]), .IN3(n6), .IN4(
        next_mac_input_01[7]), .Q(n113) );
  AO22X1 U37 ( .IN1(n7), .IN2(mac_input_01[6]), .IN3(n6), .IN4(
        next_mac_input_01[6]), .Q(n112) );
  AO22X1 U38 ( .IN1(n7), .IN2(mac_input_01[5]), .IN3(n6), .IN4(
        next_mac_input_01[5]), .Q(n111) );
  AO22X1 U39 ( .IN1(n7), .IN2(mac_input_01[4]), .IN3(n6), .IN4(
        next_mac_input_01[4]), .Q(n110) );
  AO22X1 U40 ( .IN1(n7), .IN2(mac_input_01[3]), .IN3(n6), .IN4(
        next_mac_input_01[3]), .Q(n109) );
  AO22X1 U41 ( .IN1(n7), .IN2(mac_input_01[2]), .IN3(n6), .IN4(
        next_mac_input_01[2]), .Q(n108) );
  AO22X1 U42 ( .IN1(n7), .IN2(mac_input_01[1]), .IN3(n6), .IN4(
        next_mac_input_01[1]), .Q(n107) );
  AO22X1 U43 ( .IN1(n7), .IN2(mac_input_01[0]), .IN3(n6), .IN4(
        next_mac_input_01[0]), .Q(n106) );
  AO22X1 U44 ( .IN1(n7), .IN2(mac_input_02[31]), .IN3(n6), .IN4(
        next_mac_input_02[31]), .Q(n105) );
  AO22X1 U45 ( .IN1(n7), .IN2(mac_input_02[30]), .IN3(n6), .IN4(
        next_mac_input_02[30]), .Q(n104) );
  AO22X1 U46 ( .IN1(n7), .IN2(mac_input_02[29]), .IN3(n6), .IN4(
        next_mac_input_02[29]), .Q(n103) );
  AO22X1 U47 ( .IN1(n7), .IN2(mac_input_02[28]), .IN3(n6), .IN4(
        next_mac_input_02[28]), .Q(n102) );
  AO22X1 U48 ( .IN1(n7), .IN2(mac_input_02[27]), .IN3(n6), .IN4(
        next_mac_input_02[27]), .Q(n101) );
  AO22X1 U49 ( .IN1(n7), .IN2(mac_input_02[26]), .IN3(n6), .IN4(
        next_mac_input_02[26]), .Q(n100) );
  AO22X1 U50 ( .IN1(n7), .IN2(mac_input_02[25]), .IN3(n6), .IN4(
        next_mac_input_02[25]), .Q(n99) );
  AO22X1 U51 ( .IN1(n7), .IN2(mac_input_02[24]), .IN3(n6), .IN4(
        next_mac_input_02[24]), .Q(n98) );
  AO22X1 U52 ( .IN1(n7), .IN2(mac_input_02[23]), .IN3(n6), .IN4(
        next_mac_input_02[23]), .Q(n97) );
  AO22X1 U53 ( .IN1(n7), .IN2(mac_input_02[22]), .IN3(n6), .IN4(
        next_mac_input_02[22]), .Q(n96) );
  AO22X1 U54 ( .IN1(n7), .IN2(mac_input_02[21]), .IN3(n6), .IN4(
        next_mac_input_02[21]), .Q(n95) );
  AO22X1 U55 ( .IN1(n7), .IN2(mac_input_02[20]), .IN3(n6), .IN4(
        next_mac_input_02[20]), .Q(n94) );
  AO22X1 U56 ( .IN1(n7), .IN2(mac_input_02[19]), .IN3(n6), .IN4(
        next_mac_input_02[19]), .Q(n93) );
  AO22X1 U57 ( .IN1(n7), .IN2(mac_input_02[18]), .IN3(n6), .IN4(
        next_mac_input_02[18]), .Q(n92) );
  AO22X1 U58 ( .IN1(n7), .IN2(mac_input_02[17]), .IN3(n6), .IN4(
        next_mac_input_02[17]), .Q(n91) );
  AO22X1 U59 ( .IN1(n7), .IN2(mac_input_02[16]), .IN3(n6), .IN4(
        next_mac_input_02[16]), .Q(n90) );
  AO22X1 U60 ( .IN1(n7), .IN2(mac_input_02[15]), .IN3(n6), .IN4(
        next_mac_input_02[15]), .Q(n89) );
  AO22X1 U61 ( .IN1(n7), .IN2(mac_input_02[14]), .IN3(n6), .IN4(
        next_mac_input_02[14]), .Q(n88) );
  AO22X1 U62 ( .IN1(n7), .IN2(mac_input_02[13]), .IN3(n6), .IN4(
        next_mac_input_02[13]), .Q(n87) );
  AO22X1 U63 ( .IN1(n7), .IN2(mac_input_02[12]), .IN3(n6), .IN4(
        next_mac_input_02[12]), .Q(n86) );
  AO22X1 U64 ( .IN1(n7), .IN2(mac_input_02[11]), .IN3(n6), .IN4(
        next_mac_input_02[11]), .Q(n85) );
  AO22X1 U65 ( .IN1(n7), .IN2(mac_input_02[10]), .IN3(n6), .IN4(
        next_mac_input_02[10]), .Q(n84) );
  AO22X1 U66 ( .IN1(n7), .IN2(mac_input_02[9]), .IN3(n6), .IN4(
        next_mac_input_02[9]), .Q(n83) );
  AO22X1 U67 ( .IN1(n7), .IN2(mac_input_02[8]), .IN3(n6), .IN4(
        next_mac_input_02[8]), .Q(n82) );
  AO22X1 U68 ( .IN1(n7), .IN2(mac_input_02[7]), .IN3(n6), .IN4(
        next_mac_input_02[7]), .Q(n81) );
  AO22X1 U69 ( .IN1(n7), .IN2(mac_input_02[6]), .IN3(n6), .IN4(
        next_mac_input_02[6]), .Q(n80) );
  AO22X1 U70 ( .IN1(n7), .IN2(mac_input_02[5]), .IN3(n6), .IN4(
        next_mac_input_02[5]), .Q(n79) );
  AO22X1 U71 ( .IN1(n7), .IN2(mac_input_02[4]), .IN3(n6), .IN4(
        next_mac_input_02[4]), .Q(n78) );
  AO22X1 U72 ( .IN1(n7), .IN2(mac_input_02[3]), .IN3(n6), .IN4(
        next_mac_input_02[3]), .Q(n77) );
  AO22X1 U73 ( .IN1(n7), .IN2(mac_input_02[2]), .IN3(n6), .IN4(
        next_mac_input_02[2]), .Q(n76) );
  AO22X1 U74 ( .IN1(n7), .IN2(mac_input_02[1]), .IN3(n6), .IN4(
        next_mac_input_02[1]), .Q(n75) );
  AO22X1 U75 ( .IN1(n7), .IN2(mac_input_02[0]), .IN3(n6), .IN4(
        next_mac_input_02[0]), .Q(n74) );
  AO22X1 U76 ( .IN1(n9), .IN2(weight_input_mul[31]), .IN3(n2), .IN4(
        next_weight_input_mul[31]), .Q(n73) );
  AO22X1 U77 ( .IN1(n9), .IN2(weight_input_mul[30]), .IN3(n2), .IN4(
        next_weight_input_mul[30]), .Q(n72) );
  AO22X1 U78 ( .IN1(n9), .IN2(weight_input_mul[29]), .IN3(n2), .IN4(
        next_weight_input_mul[29]), .Q(n71) );
  AO22X1 U79 ( .IN1(n9), .IN2(weight_input_mul[28]), .IN3(n2), .IN4(
        next_weight_input_mul[28]), .Q(n70) );
  AO22X1 U80 ( .IN1(n9), .IN2(weight_input_mul[27]), .IN3(n2), .IN4(
        next_weight_input_mul[27]), .Q(n69) );
  AO22X1 U81 ( .IN1(n9), .IN2(weight_input_mul[26]), .IN3(n2), .IN4(
        next_weight_input_mul[26]), .Q(n68) );
  AO22X1 U82 ( .IN1(n9), .IN2(weight_input_mul[25]), .IN3(n2), .IN4(
        next_weight_input_mul[25]), .Q(n67) );
  AO22X1 U83 ( .IN1(n9), .IN2(weight_input_mul[24]), .IN3(n2), .IN4(
        next_weight_input_mul[24]), .Q(n66) );
  AO22X1 U84 ( .IN1(n9), .IN2(weight_input_mul[23]), .IN3(n2), .IN4(
        next_weight_input_mul[23]), .Q(n65) );
  AO22X1 U85 ( .IN1(n9), .IN2(weight_input_mul[22]), .IN3(n2), .IN4(
        next_weight_input_mul[22]), .Q(n64) );
  AO22X1 U86 ( .IN1(n9), .IN2(weight_input_mul[21]), .IN3(n2), .IN4(
        next_weight_input_mul[21]), .Q(n63) );
  AO22X1 U87 ( .IN1(n9), .IN2(weight_input_mul[20]), .IN3(n2), .IN4(
        next_weight_input_mul[20]), .Q(n62) );
  AO22X1 U88 ( .IN1(n9), .IN2(weight_input_mul[19]), .IN3(n2), .IN4(
        next_weight_input_mul[19]), .Q(n61) );
  AO22X1 U89 ( .IN1(n9), .IN2(weight_input_mul[18]), .IN3(n2), .IN4(
        next_weight_input_mul[18]), .Q(n60) );
  AO22X1 U90 ( .IN1(n9), .IN2(weight_input_mul[17]), .IN3(n2), .IN4(
        next_weight_input_mul[17]), .Q(n59) );
  AO22X1 U91 ( .IN1(n9), .IN2(weight_input_mul[16]), .IN3(n2), .IN4(
        next_weight_input_mul[16]), .Q(n58) );
  AO22X1 U92 ( .IN1(n9), .IN2(weight_input_mul[15]), .IN3(n2), .IN4(
        next_weight_input_mul[15]), .Q(n57) );
  AO22X1 U93 ( .IN1(n9), .IN2(weight_input_mul[14]), .IN3(n2), .IN4(
        next_weight_input_mul[14]), .Q(n56) );
  AO22X1 U94 ( .IN1(n9), .IN2(weight_input_mul[13]), .IN3(n2), .IN4(
        next_weight_input_mul[13]), .Q(n55) );
  AO22X1 U95 ( .IN1(n9), .IN2(weight_input_mul[12]), .IN3(n2), .IN4(
        next_weight_input_mul[12]), .Q(n54) );
  AO22X1 U96 ( .IN1(n9), .IN2(weight_input_mul[11]), .IN3(n2), .IN4(
        next_weight_input_mul[11]), .Q(n53) );
  AO22X1 U97 ( .IN1(n9), .IN2(weight_input_mul[10]), .IN3(n2), .IN4(
        next_weight_input_mul[10]), .Q(n52) );
  AO22X1 U98 ( .IN1(n9), .IN2(weight_input_mul[9]), .IN3(n2), .IN4(
        next_weight_input_mul[9]), .Q(n51) );
  AO22X1 U99 ( .IN1(n9), .IN2(weight_input_mul[8]), .IN3(n2), .IN4(
        next_weight_input_mul[8]), .Q(n50) );
  AO22X1 U100 ( .IN1(n9), .IN2(weight_input_mul[7]), .IN3(n2), .IN4(
        next_weight_input_mul[7]), .Q(n49) );
  AO22X1 U101 ( .IN1(n9), .IN2(weight_input_mul[6]), .IN3(n2), .IN4(
        next_weight_input_mul[6]), .Q(n48) );
  AO22X1 U102 ( .IN1(n9), .IN2(weight_input_mul[5]), .IN3(n2), .IN4(
        next_weight_input_mul[5]), .Q(n47) );
  AO22X1 U103 ( .IN1(n9), .IN2(weight_input_mul[4]), .IN3(n2), .IN4(
        next_weight_input_mul[4]), .Q(n46) );
  AO22X1 U104 ( .IN1(n9), .IN2(weight_input_mul[3]), .IN3(n2), .IN4(
        next_weight_input_mul[3]), .Q(n45) );
  AO22X1 U105 ( .IN1(n9), .IN2(weight_input_mul[2]), .IN3(n2), .IN4(
        next_weight_input_mul[2]), .Q(n44) );
  AO22X1 U106 ( .IN1(n9), .IN2(weight_input_mul[1]), .IN3(n2), .IN4(
        next_weight_input_mul[1]), .Q(n43) );
  AO22X1 U107 ( .IN1(n9), .IN2(weight_input_mul[0]), .IN3(n2), .IN4(
        next_weight_input_mul[0]), .Q(n42) );
  AO22X1 U108 ( .IN1(n138), .IN2(mac_output[0]), .IN3(n1), .IN4(
        pre_adder_output[0]), .Q(n41) );
  AO22X1 U109 ( .IN1(n138), .IN2(mac_output[1]), .IN3(n1), .IN4(
        pre_adder_output[1]), .Q(n40) );
  AO22X1 U110 ( .IN1(n138), .IN2(mac_output[2]), .IN3(n1), .IN4(
        pre_adder_output[2]), .Q(n39) );
  AO22X1 U111 ( .IN1(n138), .IN2(mac_output[3]), .IN3(n1), .IN4(
        pre_adder_output[3]), .Q(n38) );
  AO22X1 U112 ( .IN1(n138), .IN2(mac_output[4]), .IN3(n1), .IN4(
        pre_adder_output[4]), .Q(n37) );
  AO22X1 U113 ( .IN1(n138), .IN2(mac_output[5]), .IN3(n1), .IN4(
        pre_adder_output[5]), .Q(n36) );
  AO22X1 U114 ( .IN1(n138), .IN2(mac_output[6]), .IN3(n1), .IN4(
        pre_adder_output[6]), .Q(n35) );
  AO22X1 U115 ( .IN1(n138), .IN2(mac_output[7]), .IN3(n1), .IN4(
        pre_adder_output[7]), .Q(n34) );
  AO22X1 U116 ( .IN1(n138), .IN2(mac_output[8]), .IN3(n1), .IN4(
        pre_adder_output[8]), .Q(n33) );
  AO22X1 U117 ( .IN1(n138), .IN2(mac_output[9]), .IN3(n1), .IN4(
        pre_adder_output[9]), .Q(n32) );
  AO22X1 U118 ( .IN1(n138), .IN2(mac_output[10]), .IN3(n1), .IN4(
        pre_adder_output[10]), .Q(n31) );
  AO22X1 U119 ( .IN1(n138), .IN2(mac_output[11]), .IN3(n1), .IN4(
        pre_adder_output[11]), .Q(n30) );
  AO22X1 U120 ( .IN1(n138), .IN2(mac_output[12]), .IN3(n1), .IN4(
        pre_adder_output[12]), .Q(n29) );
  AO22X1 U121 ( .IN1(n138), .IN2(mac_output[13]), .IN3(n1), .IN4(
        pre_adder_output[13]), .Q(n28) );
  AO22X1 U122 ( .IN1(n138), .IN2(mac_output[14]), .IN3(n1), .IN4(
        pre_adder_output[14]), .Q(n27) );
  AO22X1 U123 ( .IN1(n138), .IN2(mac_output[15]), .IN3(n1), .IN4(
        pre_adder_output[15]), .Q(n26) );
  AO22X1 U124 ( .IN1(n138), .IN2(mac_output[16]), .IN3(n1), .IN4(
        pre_adder_output[16]), .Q(n25) );
  AO22X1 U125 ( .IN1(n138), .IN2(mac_output[17]), .IN3(n1), .IN4(
        pre_adder_output[17]), .Q(n24) );
  AO22X1 U126 ( .IN1(n138), .IN2(mac_output[18]), .IN3(n1), .IN4(
        pre_adder_output[18]), .Q(n23) );
  AO22X1 U127 ( .IN1(n138), .IN2(mac_output[19]), .IN3(n1), .IN4(
        pre_adder_output[19]), .Q(n22) );
  AO22X1 U128 ( .IN1(n138), .IN2(mac_output[20]), .IN3(n1), .IN4(
        pre_adder_output[20]), .Q(n21) );
  AO22X1 U129 ( .IN1(n138), .IN2(mac_output[21]), .IN3(n1), .IN4(
        pre_adder_output[21]), .Q(n20) );
  AO22X1 U130 ( .IN1(n138), .IN2(mac_output[22]), .IN3(n1), .IN4(
        pre_adder_output[22]), .Q(n19) );
  AO22X1 U131 ( .IN1(n138), .IN2(mac_output[23]), .IN3(n1), .IN4(
        pre_adder_output[23]), .Q(n18) );
  AO22X1 U132 ( .IN1(n138), .IN2(mac_output[24]), .IN3(n1), .IN4(
        pre_adder_output[24]), .Q(n17) );
  AO22X1 U133 ( .IN1(n138), .IN2(mac_output[25]), .IN3(n1), .IN4(
        pre_adder_output[25]), .Q(n16) );
  AO22X1 U134 ( .IN1(n138), .IN2(mac_output[26]), .IN3(n1), .IN4(
        pre_adder_output[26]), .Q(n15) );
  AO22X1 U135 ( .IN1(n138), .IN2(mac_output[27]), .IN3(n1), .IN4(
        pre_adder_output[27]), .Q(n14) );
  AO22X1 U136 ( .IN1(n138), .IN2(mac_output[28]), .IN3(n1), .IN4(
        pre_adder_output[28]), .Q(n13) );
  AO22X1 U137 ( .IN1(n138), .IN2(mac_output[29]), .IN3(n1), .IN4(
        pre_adder_output[29]), .Q(n12) );
  AO22X1 U138 ( .IN1(n138), .IN2(mac_output[30]), .IN3(n1), .IN4(
        pre_adder_output[30]), .Q(n11) );
  AO22X1 U139 ( .IN1(n138), .IN2(mac_output[31]), .IN3(n1), .IN4(
        pre_adder_output[31]), .Q(n10) );
endmodule


module linear_function ( clk, rst_n, linear_input, linear_output );
  input [31:0] linear_input;
  output [31:0] linear_output;
  input clk, rst_n;
  wire   N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54,
         N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68,
         N69, N70, n1, n2, n3;

  DFFARX1 linear_output_reg_31_ ( .D(linear_input[31]), .CLK(clk), .RSTB(rst_n), .Q(linear_output[31]) );
  DFFARX1 linear_output_reg_29_ ( .D(N70), .CLK(clk), .RSTB(rst_n), .Q(
        linear_output[29]) );
  DFFARX1 linear_output_reg_28_ ( .D(N69), .CLK(clk), .RSTB(rst_n), .Q(
        linear_output[28]) );
  DFFARX1 linear_output_reg_27_ ( .D(N68), .CLK(clk), .RSTB(rst_n), .Q(
        linear_output[27]) );
  DFFARX1 linear_output_reg_26_ ( .D(N67), .CLK(clk), .RSTB(rst_n), .Q(
        linear_output[26]) );
  DFFARX1 linear_output_reg_25_ ( .D(N66), .CLK(clk), .RSTB(rst_n), .Q(
        linear_output[25]) );
  DFFARX1 linear_output_reg_24_ ( .D(N65), .CLK(clk), .RSTB(rst_n), .Q(
        linear_output[24]) );
  DFFARX1 linear_output_reg_23_ ( .D(N64), .CLK(clk), .RSTB(rst_n), .Q(
        linear_output[23]) );
  DFFARX1 linear_output_reg_22_ ( .D(N63), .CLK(clk), .RSTB(rst_n), .Q(
        linear_output[22]) );
  DFFARX1 linear_output_reg_21_ ( .D(N62), .CLK(clk), .RSTB(rst_n), .Q(
        linear_output[21]) );
  DFFARX1 linear_output_reg_20_ ( .D(N61), .CLK(clk), .RSTB(rst_n), .Q(
        linear_output[20]) );
  DFFARX1 linear_output_reg_19_ ( .D(N60), .CLK(clk), .RSTB(rst_n), .Q(
        linear_output[19]) );
  DFFARX1 linear_output_reg_18_ ( .D(N59), .CLK(clk), .RSTB(rst_n), .Q(
        linear_output[18]) );
  DFFARX1 linear_output_reg_17_ ( .D(N58), .CLK(clk), .RSTB(rst_n), .Q(
        linear_output[17]) );
  DFFARX1 linear_output_reg_16_ ( .D(N57), .CLK(clk), .RSTB(rst_n), .Q(
        linear_output[16]) );
  DFFARX1 linear_output_reg_15_ ( .D(N56), .CLK(clk), .RSTB(rst_n), .Q(
        linear_output[15]) );
  DFFARX1 linear_output_reg_14_ ( .D(N55), .CLK(clk), .RSTB(rst_n), .Q(
        linear_output[14]) );
  DFFARX1 linear_output_reg_13_ ( .D(N54), .CLK(clk), .RSTB(rst_n), .Q(
        linear_output[13]) );
  DFFARX1 linear_output_reg_12_ ( .D(N53), .CLK(clk), .RSTB(rst_n), .Q(
        linear_output[12]) );
  DFFARX1 linear_output_reg_11_ ( .D(N52), .CLK(clk), .RSTB(rst_n), .Q(
        linear_output[11]) );
  DFFARX1 linear_output_reg_10_ ( .D(N51), .CLK(clk), .RSTB(rst_n), .Q(
        linear_output[10]) );
  DFFARX1 linear_output_reg_9_ ( .D(N50), .CLK(clk), .RSTB(rst_n), .Q(
        linear_output[9]) );
  DFFARX1 linear_output_reg_8_ ( .D(N49), .CLK(clk), .RSTB(rst_n), .Q(
        linear_output[8]) );
  DFFARX1 linear_output_reg_7_ ( .D(N48), .CLK(clk), .RSTB(rst_n), .Q(
        linear_output[7]) );
  DFFARX1 linear_output_reg_6_ ( .D(N47), .CLK(clk), .RSTB(rst_n), .Q(
        linear_output[6]) );
  DFFARX1 linear_output_reg_5_ ( .D(N46), .CLK(clk), .RSTB(rst_n), .Q(
        linear_output[5]) );
  DFFARX1 linear_output_reg_4_ ( .D(N45), .CLK(clk), .RSTB(rst_n), .Q(
        linear_output[4]) );
  DFFARX1 linear_output_reg_3_ ( .D(N44), .CLK(clk), .RSTB(rst_n), .Q(
        linear_output[3]) );
  DFFARX1 linear_output_reg_2_ ( .D(N43), .CLK(clk), .RSTB(rst_n), .Q(
        linear_output[2]) );
  DFFARX1 linear_output_reg_1_ ( .D(N42), .CLK(clk), .RSTB(rst_n), .Q(
        linear_output[1]) );
  DFFARX1 linear_output_reg_0_ ( .D(N41), .CLK(clk), .RSTB(rst_n), .Q(
        linear_output[0]) );
  NOR2X0 U3 ( .IN1(linear_input[30]), .IN2(n2), .QN(n3) );
  AND4X1 U4 ( .IN1(linear_input[23]), .IN2(linear_input[26]), .IN3(
        linear_input[25]), .IN4(linear_input[27]), .Q(n1) );
  AND4X1 U5 ( .IN1(linear_input[24]), .IN2(linear_input[29]), .IN3(
        linear_input[28]), .IN4(n1), .Q(n2) );
  AND2X1 U6 ( .IN1(n3), .IN2(linear_input[0]), .Q(N41) );
  AND2X1 U7 ( .IN1(n3), .IN2(linear_input[1]), .Q(N42) );
  AND2X1 U8 ( .IN1(n3), .IN2(linear_input[2]), .Q(N43) );
  AND2X1 U9 ( .IN1(n3), .IN2(linear_input[3]), .Q(N44) );
  AND2X1 U10 ( .IN1(n3), .IN2(linear_input[4]), .Q(N45) );
  AND2X1 U11 ( .IN1(n3), .IN2(linear_input[5]), .Q(N46) );
  AND2X1 U12 ( .IN1(n3), .IN2(linear_input[6]), .Q(N47) );
  AND2X1 U13 ( .IN1(n3), .IN2(linear_input[7]), .Q(N48) );
  AND2X1 U14 ( .IN1(n3), .IN2(linear_input[8]), .Q(N49) );
  AND2X1 U15 ( .IN1(n3), .IN2(linear_input[9]), .Q(N50) );
  AND2X1 U16 ( .IN1(n3), .IN2(linear_input[10]), .Q(N51) );
  AND2X1 U17 ( .IN1(n3), .IN2(linear_input[11]), .Q(N52) );
  AND2X1 U18 ( .IN1(n3), .IN2(linear_input[12]), .Q(N53) );
  AND2X1 U19 ( .IN1(n3), .IN2(linear_input[13]), .Q(N54) );
  AND2X1 U20 ( .IN1(n3), .IN2(linear_input[14]), .Q(N55) );
  AND2X1 U21 ( .IN1(n3), .IN2(linear_input[15]), .Q(N56) );
  AND2X1 U22 ( .IN1(n3), .IN2(linear_input[16]), .Q(N57) );
  AND2X1 U23 ( .IN1(n3), .IN2(linear_input[17]), .Q(N58) );
  AND2X1 U24 ( .IN1(n3), .IN2(linear_input[18]), .Q(N59) );
  AND2X1 U25 ( .IN1(n3), .IN2(linear_input[19]), .Q(N60) );
  AND2X1 U26 ( .IN1(n3), .IN2(linear_input[20]), .Q(N61) );
  AND2X1 U27 ( .IN1(n3), .IN2(linear_input[21]), .Q(N62) );
  AND2X1 U28 ( .IN1(n3), .IN2(linear_input[22]), .Q(N63) );
  OR2X1 U29 ( .IN1(linear_input[30]), .IN2(linear_input[23]), .Q(N64) );
  OR2X1 U30 ( .IN1(linear_input[30]), .IN2(linear_input[24]), .Q(N65) );
  OR2X1 U31 ( .IN1(linear_input[30]), .IN2(linear_input[25]), .Q(N66) );
  OR2X1 U32 ( .IN1(linear_input[30]), .IN2(linear_input[26]), .Q(N67) );
  OR2X1 U33 ( .IN1(linear_input[30]), .IN2(linear_input[27]), .Q(N68) );
  OR2X1 U34 ( .IN1(linear_input[30]), .IN2(linear_input[28]), .Q(N69) );
  OR2X1 U35 ( .IN1(linear_input[30]), .IN2(linear_input[29]), .Q(N70) );
endmodule


module step_function ( clk, rst_n, step_input, step_output );
  input [31:0] step_input;
  output [31:0] step_output;
  input clk, rst_n;


  DFFASX1 step_output_reg_23_ ( .D(step_input[31]), .CLK(clk), .SETB(rst_n), 
        .QN(step_output[23]) );
endmodule


module sigmoid_floating_point_compare ( clk, rst_n, factor_input, factor_a, 
        factor_b, factor_c, factor_d );
  input [31:0] factor_input;
  output [31:0] factor_a;
  output [31:0] factor_b;
  output [31:0] factor_c;
  output [31:0] factor_d;
  input clk, rst_n;
  wire   N55, N56, N57, N58, N151, N154, N155, N156, N157, N158, N159, N161,
         N162, N163, N165, N166, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n93, n94, n95, n96, n133, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n90, n91, n92, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177;
  wire   [2:0] case_num;

  DFFARX1 case_num_reg_3_ ( .D(N58), .CLK(clk), .RSTB(rst_n), .Q(n4), .QN(n95)
         );
  DFFARX1 case_num_reg_2_ ( .D(N57), .CLK(clk), .RSTB(rst_n), .Q(case_num[2]), 
        .QN(n3) );
  DFFARX1 case_num_reg_1_ ( .D(N56), .CLK(clk), .RSTB(rst_n), .Q(case_num[1]), 
        .QN(n2) );
  DFFARX1 case_num_reg_0_ ( .D(N55), .CLK(clk), .RSTB(rst_n), .Q(case_num[0]), 
        .QN(n1) );
  DFFARX1 factor_a_reg_31_ ( .D(N163), .CLK(clk), .RSTB(rst_n), .Q(
        factor_a[31]) );
  DFFARX1 factor_a_reg_29_ ( .D(N165), .CLK(clk), .RSTB(rst_n), .Q(
        factor_a[29]) );
  DFFARX1 factor_a_reg_28_ ( .D(N165), .CLK(clk), .RSTB(rst_n), .Q(
        factor_a[28]) );
  DFFARX1 factor_a_reg_27_ ( .D(N165), .CLK(clk), .RSTB(rst_n), .Q(
        factor_a[27]) );
  DFFASX1 factor_a_reg_26_ ( .D(n133), .CLK(clk), .SETB(rst_n), .QN(
        factor_a[26]) );
  DFFARX1 factor_a_reg_25_ ( .D(N151), .CLK(clk), .RSTB(rst_n), .Q(
        factor_a[25]) );
  DFFARX1 factor_a_reg_24_ ( .D(N161), .CLK(clk), .RSTB(rst_n), .Q(
        factor_a[24]) );
  DFFARX1 factor_a_reg_23_ ( .D(N154), .CLK(clk), .RSTB(rst_n), .Q(
        factor_a[23]) );
  DFFARX1 factor_a_reg_22_ ( .D(N163), .CLK(clk), .RSTB(rst_n), .Q(
        factor_a[22]) );
  DFFARX1 factor_a_reg_21_ ( .D(N162), .CLK(clk), .RSTB(rst_n), .Q(
        factor_a[21]) );
  DFFARX1 factor_a_reg_20_ ( .D(N161), .CLK(clk), .RSTB(rst_n), .Q(
        factor_a[20]) );
  DFFASX1 factor_a_reg_19_ ( .D(n93), .CLK(clk), .SETB(rst_n), .QN(
        factor_a[19]) );
  DFFARX1 factor_a_reg_18_ ( .D(N159), .CLK(clk), .RSTB(rst_n), .Q(
        factor_a[18]) );
  DFFARX1 factor_a_reg_17_ ( .D(N156), .CLK(clk), .RSTB(rst_n), .Q(
        factor_a[17]) );
  DFFARX1 factor_a_reg_16_ ( .D(N157), .CLK(clk), .RSTB(rst_n), .Q(
        factor_a[16]) );
  DFFARX1 factor_a_reg_15_ ( .D(N157), .CLK(clk), .RSTB(rst_n), .Q(
        factor_a[15]) );
  DFFARX1 factor_a_reg_14_ ( .D(N158), .CLK(clk), .RSTB(rst_n), .Q(
        factor_a[14]) );
  DFFASX1 factor_a_reg_12_ ( .D(n94), .CLK(clk), .SETB(rst_n), .QN(
        factor_a[12]) );
  DFFARX1 factor_a_reg_11_ ( .D(N154), .CLK(clk), .RSTB(rst_n), .Q(
        factor_a[11]) );
  DFFARX1 factor_a_reg_10_ ( .D(N157), .CLK(clk), .RSTB(rst_n), .Q(
        factor_a[10]) );
  DFFARX1 factor_a_reg_9_ ( .D(N156), .CLK(clk), .RSTB(rst_n), .Q(factor_a[9])
         );
  DFFARX1 factor_a_reg_8_ ( .D(N155), .CLK(clk), .RSTB(rst_n), .Q(factor_a[8])
         );
  DFFARX1 factor_a_reg_7_ ( .D(N154), .CLK(clk), .RSTB(rst_n), .Q(factor_a[7])
         );
  DFFARX1 factor_a_reg_5_ ( .D(N154), .CLK(clk), .RSTB(rst_n), .Q(factor_a[5])
         );
  DFFASX1 factor_a_reg_4_ ( .D(n94), .CLK(clk), .SETB(rst_n), .QN(factor_a[4])
         );
  DFFASX1 factor_a_reg_3_ ( .D(n96), .CLK(clk), .SETB(rst_n), .QN(factor_a[3])
         );
  DFFARX1 factor_a_reg_2_ ( .D(N165), .CLK(clk), .RSTB(rst_n), .Q(factor_a[2])
         );
  DFFARX1 factor_a_reg_1_ ( .D(N151), .CLK(clk), .RSTB(rst_n), .Q(factor_a[1])
         );
  DFFARX1 factor_a_reg_0_ ( .D(N151), .CLK(clk), .RSTB(rst_n), .Q(factor_a[0])
         );
  DFFARX1 factor_b_reg_31_ ( .D(N166), .CLK(clk), .RSTB(rst_n), .Q(
        factor_b[31]) );
  DFFARX1 factor_b_reg_29_ ( .D(N165), .CLK(clk), .RSTB(rst_n), .Q(
        factor_b[29]) );
  DFFARX1 factor_b_reg_28_ ( .D(N165), .CLK(clk), .RSTB(rst_n), .Q(
        factor_b[28]) );
  DFFARX1 factor_b_reg_27_ ( .D(N165), .CLK(clk), .RSTB(rst_n), .Q(
        factor_b[27]) );
  DFFARX1 factor_b_reg_26_ ( .D(N154), .CLK(clk), .RSTB(rst_n), .Q(
        factor_b[26]) );
  DFFASX1 factor_b_reg_25_ ( .D(n133), .CLK(clk), .SETB(rst_n), .QN(
        factor_b[25]) );
  DFFARX1 factor_b_reg_24_ ( .D(N162), .CLK(clk), .RSTB(rst_n), .Q(
        factor_b[24]) );
  DFFARX1 factor_b_reg_23_ ( .D(N155), .CLK(clk), .RSTB(rst_n), .Q(
        factor_b[23]) );
  DFFARX1 factor_b_reg_21_ ( .D(N158), .CLK(clk), .RSTB(rst_n), .Q(
        factor_b[21]) );
  DFFASX1 factor_b_reg_20_ ( .D(n94), .CLK(clk), .SETB(rst_n), .QN(
        factor_b[20]) );
  DFFARX1 factor_b_reg_17_ ( .D(N165), .CLK(clk), .RSTB(rst_n), .Q(
        factor_b[17]) );
  DFFARX1 factor_b_reg_16_ ( .D(N156), .CLK(clk), .RSTB(rst_n), .Q(
        factor_b[16]) );
  DFFARX1 factor_b_reg_15_ ( .D(N158), .CLK(clk), .RSTB(rst_n), .Q(
        factor_b[15]) );
  DFFASX1 factor_b_reg_14_ ( .D(n133), .CLK(clk), .SETB(rst_n), .QN(
        factor_b[14]) );
  DFFARX1 factor_b_reg_13_ ( .D(N158), .CLK(clk), .RSTB(rst_n), .Q(
        factor_b[13]) );
  DFFASX1 factor_b_reg_12_ ( .D(n94), .CLK(clk), .SETB(rst_n), .QN(
        factor_b[12]) );
  DFFARX1 factor_b_reg_11_ ( .D(N154), .CLK(clk), .RSTB(rst_n), .Q(
        factor_b[11]) );
  DFFARX1 factor_b_reg_10_ ( .D(N162), .CLK(clk), .RSTB(rst_n), .Q(
        factor_b[10]) );
  DFFARX1 factor_b_reg_9_ ( .D(N163), .CLK(clk), .RSTB(rst_n), .Q(factor_b[9])
         );
  DFFASX1 factor_b_reg_8_ ( .D(n96), .CLK(clk), .SETB(rst_n), .QN(factor_b[8])
         );
  DFFASX1 factor_b_reg_7_ ( .D(n96), .CLK(clk), .SETB(rst_n), .QN(factor_b[7])
         );
  DFFARX1 factor_b_reg_6_ ( .D(N151), .CLK(clk), .RSTB(rst_n), .Q(factor_b[6])
         );
  DFFARX1 factor_b_reg_5_ ( .D(N156), .CLK(clk), .RSTB(rst_n), .Q(factor_b[5])
         );
  DFFASX1 factor_b_reg_4_ ( .D(n96), .CLK(clk), .SETB(rst_n), .QN(factor_b[4])
         );
  DFFARX1 factor_b_reg_3_ ( .D(N156), .CLK(clk), .RSTB(rst_n), .Q(factor_b[3])
         );
  DFFARX1 factor_b_reg_2_ ( .D(N154), .CLK(clk), .RSTB(rst_n), .Q(factor_b[2])
         );
  DFFARX1 factor_b_reg_1_ ( .D(N156), .CLK(clk), .RSTB(rst_n), .Q(factor_b[1])
         );
  DFFASX1 factor_b_reg_0_ ( .D(n96), .CLK(clk), .SETB(rst_n), .QN(factor_b[0])
         );
  DFFX1 factor_c_reg_31_ ( .D(n89), .CLK(clk), .Q(factor_c[31]) );
  DFFX1 factor_c_reg_29_ ( .D(n88), .CLK(clk), .Q(factor_c[29]) );
  DFFX1 factor_c_reg_28_ ( .D(n87), .CLK(clk), .Q(factor_c[28]) );
  DFFX1 factor_c_reg_27_ ( .D(n86), .CLK(clk), .Q(factor_c[27]) );
  DFFX1 factor_c_reg_26_ ( .D(n85), .CLK(clk), .Q(factor_c[26]) );
  DFFX1 factor_c_reg_25_ ( .D(n84), .CLK(clk), .Q(factor_c[25]) );
  DFFX1 factor_c_reg_24_ ( .D(n83), .CLK(clk), .Q(factor_c[24]) );
  DFFX1 factor_c_reg_23_ ( .D(n82), .CLK(clk), .Q(factor_c[23]) );
  DFFX1 factor_c_reg_22_ ( .D(n81), .CLK(clk), .Q(factor_c[22]) );
  DFFX1 factor_c_reg_21_ ( .D(n80), .CLK(clk), .Q(factor_c[21]) );
  DFFX1 factor_c_reg_19_ ( .D(n79), .CLK(clk), .Q(factor_c[19]) );
  DFFX1 factor_c_reg_18_ ( .D(n78), .CLK(clk), .Q(factor_c[18]) );
  DFFX1 factor_c_reg_17_ ( .D(n77), .CLK(clk), .Q(factor_c[17]) );
  DFFX1 factor_c_reg_16_ ( .D(n76), .CLK(clk), .Q(factor_c[16]) );
  DFFX1 factor_c_reg_15_ ( .D(n75), .CLK(clk), .Q(factor_c[15]) );
  DFFX1 factor_c_reg_14_ ( .D(n74), .CLK(clk), .Q(factor_c[14]) );
  DFFX1 factor_c_reg_13_ ( .D(n73), .CLK(clk), .Q(factor_c[13]) );
  DFFX1 factor_c_reg_11_ ( .D(n72), .CLK(clk), .Q(factor_c[11]) );
  DFFX1 factor_c_reg_10_ ( .D(n71), .CLK(clk), .Q(factor_c[10]) );
  DFFX1 factor_c_reg_9_ ( .D(n70), .CLK(clk), .Q(factor_c[9]) );
  DFFX1 factor_c_reg_8_ ( .D(n69), .CLK(clk), .Q(factor_c[8]) );
  DFFX1 factor_c_reg_7_ ( .D(n68), .CLK(clk), .Q(factor_c[7]) );
  DFFX1 factor_c_reg_6_ ( .D(n67), .CLK(clk), .Q(factor_c[6]) );
  DFFX1 factor_c_reg_5_ ( .D(n66), .CLK(clk), .Q(factor_c[5]) );
  DFFX1 factor_c_reg_4_ ( .D(n65), .CLK(clk), .Q(factor_c[4]) );
  DFFX1 factor_c_reg_3_ ( .D(n64), .CLK(clk), .Q(factor_c[3]) );
  DFFX1 factor_c_reg_2_ ( .D(n63), .CLK(clk), .Q(factor_c[2]) );
  DFFX1 factor_c_reg_0_ ( .D(n62), .CLK(clk), .Q(factor_c[0]) );
  DFFX1 factor_d_reg_31_ ( .D(n61), .CLK(clk), .Q(factor_d[31]) );
  DFFX1 factor_d_reg_29_ ( .D(n60), .CLK(clk), .Q(factor_d[29]) );
  DFFX1 factor_d_reg_28_ ( .D(n59), .CLK(clk), .Q(factor_d[28]) );
  DFFX1 factor_d_reg_27_ ( .D(n58), .CLK(clk), .Q(factor_d[27]) );
  DFFX1 factor_d_reg_26_ ( .D(n57), .CLK(clk), .Q(factor_d[26]) );
  DFFX1 factor_d_reg_25_ ( .D(n56), .CLK(clk), .Q(factor_d[25]) );
  DFFX1 factor_d_reg_24_ ( .D(n55), .CLK(clk), .Q(factor_d[24]) );
  DFFX1 factor_d_reg_23_ ( .D(n54), .CLK(clk), .Q(factor_d[23]) );
  DFFX1 factor_d_reg_22_ ( .D(n53), .CLK(clk), .Q(factor_d[22]) );
  DFFX1 factor_d_reg_21_ ( .D(n52), .CLK(clk), .Q(factor_d[21]) );
  DFFX1 factor_d_reg_20_ ( .D(n51), .CLK(clk), .Q(factor_d[20]) );
  DFFX1 factor_d_reg_19_ ( .D(n50), .CLK(clk), .Q(factor_d[19]) );
  DFFX1 factor_d_reg_18_ ( .D(n49), .CLK(clk), .Q(factor_d[18]) );
  DFFX1 factor_d_reg_17_ ( .D(n48), .CLK(clk), .Q(factor_d[17]) );
  DFFX1 factor_d_reg_16_ ( .D(n47), .CLK(clk), .Q(factor_d[16]) );
  DFFX1 factor_d_reg_15_ ( .D(n46), .CLK(clk), .Q(factor_d[15]) );
  DFFX1 factor_d_reg_13_ ( .D(n45), .CLK(clk), .Q(factor_d[13]) );
  DFFX1 factor_d_reg_12_ ( .D(n44), .CLK(clk), .Q(factor_d[12]) );
  DFFX1 factor_d_reg_11_ ( .D(n43), .CLK(clk), .Q(factor_d[11]) );
  DFFX1 factor_d_reg_10_ ( .D(n42), .CLK(clk), .Q(factor_d[10]) );
  DFFX1 factor_d_reg_9_ ( .D(n41), .CLK(clk), .Q(factor_d[9]) );
  DFFX1 factor_d_reg_8_ ( .D(n40), .CLK(clk), .Q(factor_d[8]) );
  DFFX1 factor_d_reg_7_ ( .D(n39), .CLK(clk), .Q(factor_d[7]) );
  DFFX1 factor_d_reg_6_ ( .D(n38), .CLK(clk), .Q(factor_d[6]) );
  DFFX1 factor_d_reg_5_ ( .D(n37), .CLK(clk), .Q(factor_d[5]) );
  DFFX1 factor_d_reg_4_ ( .D(n36), .CLK(clk), .Q(factor_d[4]) );
  DFFX1 factor_d_reg_3_ ( .D(n35), .CLK(clk), .Q(factor_d[3]) );
  DFFX1 factor_d_reg_2_ ( .D(n34), .CLK(clk), .Q(factor_d[2]) );
  DFFX1 factor_d_reg_1_ ( .D(n33), .CLK(clk), .Q(factor_d[1]) );
  DFFX1 factor_d_reg_0_ ( .D(n32), .CLK(clk), .Q(factor_d[0]) );
  INVX1 U3 ( .INP(rst_n), .ZN(n31) );
  NAND2X0 U4 ( .IN1(n9), .IN2(n10), .QN(n108) );
  NAND2X0 U5 ( .IN1(n19), .IN2(n163), .QN(n20) );
  NAND2X0 U6 ( .IN1(n174), .IN2(n176), .QN(n19) );
  NAND2X0 U7 ( .IN1(n169), .IN2(n157), .QN(n163) );
  NAND2X0 U8 ( .IN1(case_num[2]), .IN2(n157), .QN(n166) );
  NAND2X0 U9 ( .IN1(n124), .IN2(n15), .QN(n126) );
  NAND2X0 U10 ( .IN1(n7), .IN2(n8), .QN(n113) );
  NAND2X0 U11 ( .IN1(n106), .IN2(n139), .QN(n145) );
  NAND2X0 U12 ( .IN1(n11), .IN2(n12), .QN(n33) );
  NAND2X0 U13 ( .IN1(n31), .IN2(factor_d[1]), .QN(n12) );
  NAND2X0 U14 ( .IN1(n5), .IN2(n6), .QN(n39) );
  NAND2X0 U15 ( .IN1(n31), .IN2(factor_d[7]), .QN(n6) );
  NAND2X0 U16 ( .IN1(n156), .IN2(n158), .QN(n41) );
  NAND2X0 U17 ( .IN1(n159), .IN2(n158), .QN(n45) );
  NAND2X0 U18 ( .IN1(n161), .IN2(n160), .QN(n46) );
  NAND2X0 U19 ( .IN1(n31), .IN2(factor_d[15]), .QN(n161) );
  NAND2X0 U20 ( .IN1(n31), .IN2(factor_d[16]), .QN(n22) );
  NAND2X0 U21 ( .IN1(n162), .IN2(n163), .QN(n48) );
  NAND2X0 U22 ( .IN1(n164), .IN2(n163), .QN(n49) );
  NAND2X0 U23 ( .IN1(n31), .IN2(factor_d[18]), .QN(n164) );
  NAND2X0 U24 ( .IN1(n165), .IN2(n166), .QN(n51) );
  NAND2X0 U25 ( .IN1(n31), .IN2(factor_d[20]), .QN(n165) );
  NAND2X0 U26 ( .IN1(n167), .IN2(n166), .QN(n52) );
  NAND2X0 U27 ( .IN1(n31), .IN2(factor_d[21]), .QN(n167) );
  NAND2X0 U28 ( .IN1(n173), .IN2(n149), .QN(N155) );
  NAND2X0 U29 ( .IN1(N151), .IN2(n18), .QN(n94) );
  NAND2X0 U30 ( .IN1(n93), .IN2(n133), .QN(N158) );
  NAND2X0 U31 ( .IN1(n146), .IN2(n133), .QN(N156) );
  NAND2X0 U32 ( .IN1(n23), .IN2(n133), .QN(N159) );
  NAND2X0 U33 ( .IN1(n94), .IN2(n133), .QN(N162) );
  NAND2X0 U34 ( .IN1(n173), .IN2(n96), .QN(N154) );
  NAND2X0 U35 ( .IN1(n94), .IN2(n96), .QN(N161) );
  NAND2X0 U36 ( .IN1(n151), .IN2(n150), .QN(N165) );
  NAND2X0 U37 ( .IN1(n96), .IN2(n133), .QN(N163) );
  NAND2X0 U38 ( .IN1(n145), .IN2(n144), .QN(N57) );
  NAND2X0 U39 ( .IN1(factor_input[22]), .IN2(n105), .QN(n139) );
  INVX0 U40 ( .INP(n146), .ZN(N157) );
  NOR2X0 U41 ( .IN1(n31), .IN2(n94), .QN(n175) );
  NOR2X0 U42 ( .IN1(n96), .IN2(n31), .QN(n177) );
  INVX0 U43 ( .INP(n153), .ZN(n96) );
  NOR2X0 U44 ( .IN1(n1), .IN2(n147), .QN(n153) );
  NAND2X0 U45 ( .IN1(n95), .IN2(case_num[1]), .QN(n173) );
  NAND2X0 U46 ( .IN1(factor_input[20]), .IN2(n112), .QN(n8) );
  NAND2X0 U47 ( .IN1(factor_input[7]), .IN2(n107), .QN(n10) );
  NOR2X0 U48 ( .IN1(factor_input[9]), .IN2(factor_input[8]), .QN(n9) );
  NOR2X0 U49 ( .IN1(factor_input[22]), .IN2(factor_input[21]), .QN(n7) );
  NOR2X0 U50 ( .IN1(n154), .IN2(n175), .QN(n11) );
  NOR2X0 U51 ( .IN1(n155), .IN2(n154), .QN(n5) );
  INVX0 U52 ( .INP(factor_input[6]), .ZN(n13) );
  INVX0 U53 ( .INP(factor_input[9]), .ZN(n14) );
  INVX0 U54 ( .INP(factor_input[18]), .ZN(n15) );
  INVX0 U55 ( .INP(factor_input[23]), .ZN(n16) );
  INVX0 U56 ( .INP(factor_input[30]), .ZN(n17) );
  NOR2X0 U57 ( .IN1(n31), .IN2(n173), .QN(n157) );
  NOR2X0 U58 ( .IN1(n1), .IN2(n166), .QN(n154) );
  INVX0 U59 ( .INP(n173), .ZN(N151) );
  MUX21X1 U60 ( .IN1(n1), .IN2(case_num[0]), .S(n3), .Q(n18) );
  NOR2X0 U61 ( .IN1(n18), .IN2(n173), .QN(n174) );
  INVX0 U62 ( .INP(n31), .ZN(n176) );
  NOR2X0 U63 ( .IN1(case_num[2]), .IN2(n1), .QN(n169) );
  AO21X1 U64 ( .IN1(n31), .IN2(factor_d[2]), .IN3(n20), .Q(n34) );
  AO21X1 U65 ( .IN1(n31), .IN2(factor_d[12]), .IN3(n20), .Q(n44) );
  INVX0 U66 ( .INP(n175), .ZN(n21) );
  NAND2X0 U67 ( .IN1(n157), .IN2(n1), .QN(n160) );
  NAND3X0 U68 ( .IN1(n22), .IN2(n21), .IN3(n160), .QN(n47) );
  INVX0 U69 ( .INP(n174), .ZN(n93) );
  NAND3X0 U70 ( .IN1(n95), .IN2(case_num[2]), .IN3(n2), .QN(n133) );
  NAND3X0 U71 ( .IN1(n3), .IN2(n2), .IN3(n95), .QN(n147) );
  NOR2X0 U72 ( .IN1(n174), .IN2(n153), .QN(n146) );
  INVX0 U73 ( .INP(N161), .ZN(n23) );
  NAND2X0 U74 ( .IN1(case_num[0]), .IN2(n95), .QN(n150) );
  OAI22X1 U75 ( .IN1(case_num[1]), .IN2(n150), .IN3(n3), .IN4(n173), .QN(N166)
         );
  OR4X1 U76 ( .IN1(factor_input[24]), .IN2(factor_input[25]), .IN3(
        factor_input[26]), .IN4(factor_input[27]), .Q(n24) );
  NOR3X0 U77 ( .IN1(factor_input[28]), .IN2(factor_input[29]), .IN3(n24), .QN(
        n92) );
  NOR2X0 U78 ( .IN1(n17), .IN2(n92), .QN(n141) );
  INVX0 U79 ( .INP(n141), .ZN(n97) );
  AND3X1 U80 ( .IN1(factor_input[2]), .IN2(factor_input[1]), .IN3(
        factor_input[0]), .Q(n25) );
  NOR4X0 U81 ( .IN1(factor_input[4]), .IN2(factor_input[3]), .IN3(
        factor_input[5]), .IN4(n25), .QN(n26) );
  NAND2X0 U82 ( .IN1(factor_input[7]), .IN2(factor_input[6]), .QN(n116) );
  NOR2X0 U83 ( .IN1(n26), .IN2(n116), .QN(n28) );
  OR4X1 U84 ( .IN1(factor_input[13]), .IN2(factor_input[11]), .IN3(
        factor_input[10]), .IN4(factor_input[14]), .Q(n27) );
  AO221X1 U85 ( .IN1(factor_input[9]), .IN2(factor_input[8]), .IN3(
        factor_input[9]), .IN4(n28), .IN5(n27), .Q(n29) );
  OR3X1 U86 ( .IN1(factor_input[13]), .IN2(factor_input[12]), .IN3(
        factor_input[14]), .Q(n110) );
  AND3X1 U87 ( .IN1(factor_input[15]), .IN2(n29), .IN3(n110), .Q(n30) );
  OA21X1 U88 ( .IN1(factor_input[16]), .IN2(n30), .IN3(factor_input[17]), .Q(
        n90) );
  AO21X1 U89 ( .IN1(factor_input[18]), .IN2(n90), .IN3(factor_input[19]), .Q(
        n91) );
  NAND4X0 U90 ( .IN1(factor_input[20]), .IN2(factor_input[22]), .IN3(
        factor_input[21]), .IN4(n91), .QN(n127) );
  AND2X1 U91 ( .IN1(n92), .IN2(factor_input[30]), .Q(n136) );
  NAND2X0 U92 ( .IN1(n136), .IN2(factor_input[23]), .QN(n140) );
  NOR2X0 U93 ( .IN1(n140), .IN2(factor_input[31]), .QN(n106) );
  INVX0 U94 ( .INP(n106), .ZN(n138) );
  OA22X1 U95 ( .IN1(factor_input[31]), .IN2(n97), .IN3(n127), .IN4(n138), .Q(
        n137) );
  NOR2X0 U96 ( .IN1(factor_input[7]), .IN2(factor_input[8]), .QN(n100) );
  NAND4X0 U97 ( .IN1(factor_input[4]), .IN2(factor_input[3]), .IN3(
        factor_input[5]), .IN4(factor_input[2]), .QN(n117) );
  INVX0 U98 ( .INP(n117), .ZN(n98) );
  NAND2X0 U99 ( .IN1(n98), .IN2(factor_input[1]), .QN(n99) );
  NAND4X0 U100 ( .IN1(n100), .IN2(n14), .IN3(n99), .IN4(n13), .QN(n101) );
  OA221X1 U101 ( .IN1(factor_input[11]), .IN2(factor_input[10]), .IN3(
        factor_input[11]), .IN4(n101), .IN5(factor_input[12]), .Q(n102) );
  OR2X1 U102 ( .IN1(factor_input[15]), .IN2(factor_input[14]), .Q(n122) );
  OR4X1 U103 ( .IN1(factor_input[16]), .IN2(factor_input[13]), .IN3(n102), 
        .IN4(n122), .Q(n103) );
  OA221X1 U104 ( .IN1(factor_input[18]), .IN2(factor_input[17]), .IN3(
        factor_input[18]), .IN4(n103), .IN5(factor_input[19]), .Q(n104) );
  OR3X1 U105 ( .IN1(n104), .IN2(factor_input[20]), .IN3(factor_input[21]), .Q(
        n105) );
  NAND4X0 U106 ( .IN1(factor_input[24]), .IN2(factor_input[25]), .IN3(
        factor_input[26]), .IN4(factor_input[27]), .QN(n115) );
  AO221X1 U107 ( .IN1(factor_input[5]), .IN2(factor_input[4]), .IN3(
        factor_input[5]), .IN4(factor_input[3]), .IN5(factor_input[6]), .Q(
        n107) );
  AND3X1 U108 ( .IN1(factor_input[10]), .IN2(factor_input[11]), .IN3(n108), 
        .Q(n109) );
  OR4X1 U109 ( .IN1(n110), .IN2(factor_input[17]), .IN3(factor_input[16]), 
        .IN4(n109), .Q(n111) );
  AO221X1 U110 ( .IN1(factor_input[18]), .IN2(factor_input[15]), .IN3(
        factor_input[18]), .IN4(n111), .IN5(factor_input[19]), .Q(n112) );
  NAND3X0 U111 ( .IN1(factor_input[29]), .IN2(factor_input[28]), .IN3(n113), 
        .QN(n114) );
  NOR4X0 U112 ( .IN1(factor_input[30]), .IN2(n16), .IN3(n115), .IN4(n114), 
        .QN(n135) );
  OA21X1 U113 ( .IN1(factor_input[9]), .IN2(factor_input[10]), .IN3(
        factor_input[11]), .Q(n121) );
  NOR2X0 U114 ( .IN1(n117), .IN2(n116), .QN(n118) );
  AO221X1 U115 ( .IN1(n118), .IN2(factor_input[1]), .IN3(n118), .IN4(
        factor_input[0]), .IN5(factor_input[10]), .Q(n120) );
  OR3X1 U116 ( .IN1(factor_input[13]), .IN2(factor_input[12]), .IN3(
        factor_input[15]), .Q(n119) );
  AO221X1 U117 ( .IN1(n121), .IN2(factor_input[8]), .IN3(n121), .IN4(n120), 
        .IN5(n119), .Q(n123) );
  NAND4X0 U118 ( .IN1(factor_input[16]), .IN2(factor_input[17]), .IN3(n123), 
        .IN4(n122), .QN(n124) );
  AND3X1 U119 ( .IN1(factor_input[22]), .IN2(factor_input[20]), .IN3(
        factor_input[21]), .Q(n125) );
  NAND3X0 U120 ( .IN1(n126), .IN2(n125), .IN3(factor_input[19]), .QN(n131) );
  INVX0 U121 ( .INP(n127), .ZN(n128) );
  NOR2X0 U122 ( .IN1(n128), .IN2(n139), .QN(n129) );
  OA221X1 U123 ( .IN1(factor_input[23]), .IN2(n131), .IN3(n16), .IN4(n129), 
        .IN5(n136), .Q(n130) );
  OAI21X1 U124 ( .IN1(n135), .IN2(n130), .IN3(factor_input[31]), .QN(n134) );
  OR2X1 U125 ( .IN1(n136), .IN2(n135), .Q(n143) );
  AO221X1 U126 ( .IN1(n143), .IN2(factor_input[23]), .IN3(n143), .IN4(n131), 
        .IN5(factor_input[31]), .Q(n132) );
  NAND4X0 U127 ( .IN1(n137), .IN2(n145), .IN3(n134), .IN4(n132), .QN(N55) );
  AO221X1 U128 ( .IN1(n136), .IN2(n139), .IN3(n136), .IN4(n16), .IN5(n135), 
        .Q(N56) );
  OAI21X1 U129 ( .IN1(n139), .IN2(n138), .IN3(n137), .QN(N58) );
  INVX0 U130 ( .INP(n140), .ZN(n142) );
  AO221X1 U131 ( .IN1(n143), .IN2(factor_input[31]), .IN3(n143), .IN4(n142), 
        .IN5(n141), .Q(n144) );
  MUX21X1 U132 ( .IN1(factor_d[4]), .IN2(N161), .S(n176), .Q(n36) );
  MUX21X1 U133 ( .IN1(factor_d[5]), .IN2(N157), .S(n176), .Q(n37) );
  MUX21X1 U134 ( .IN1(factor_d[19]), .IN2(N157), .S(n176), .Q(n50) );
  MUX21X1 U135 ( .IN1(factor_d[25]), .IN2(n147), .S(n176), .Q(n56) );
  OA21X1 U136 ( .IN1(case_num[0]), .IN2(n147), .IN3(n176), .Q(n148) );
  AO21X1 U137 ( .IN1(n31), .IN2(factor_d[26]), .IN3(n148), .Q(n57) );
  AO21X1 U138 ( .IN1(n31), .IN2(factor_d[27]), .IN3(n148), .Q(n58) );
  AO21X1 U139 ( .IN1(n31), .IN2(factor_d[28]), .IN3(n148), .Q(n59) );
  AO21X1 U140 ( .IN1(n31), .IN2(factor_d[29]), .IN3(n148), .Q(n60) );
  MUX21X1 U141 ( .IN1(factor_c[0]), .IN2(N161), .S(n176), .Q(n62) );
  MUX21X1 U142 ( .IN1(factor_c[5]), .IN2(N157), .S(n176), .Q(n66) );
  MUX21X1 U143 ( .IN1(factor_c[8]), .IN2(N157), .S(n176), .Q(n69) );
  MUX21X1 U144 ( .IN1(factor_c[11]), .IN2(N157), .S(n176), .Q(n72) );
  MUX21X1 U145 ( .IN1(factor_c[13]), .IN2(N161), .S(n176), .Q(n73) );
  MUX21X1 U146 ( .IN1(factor_c[14]), .IN2(N161), .S(n176), .Q(n74) );
  MUX21X1 U147 ( .IN1(factor_c[15]), .IN2(N157), .S(n176), .Q(n75) );
  MUX21X1 U148 ( .IN1(factor_c[18]), .IN2(N161), .S(n176), .Q(n78) );
  NAND2X0 U149 ( .IN1(case_num[2]), .IN2(n95), .QN(n149) );
  MUX21X1 U150 ( .IN1(factor_c[25]), .IN2(N155), .S(n176), .Q(n84) );
  INVX0 U151 ( .INP(N155), .ZN(n151) );
  MUX21X1 U152 ( .IN1(factor_c[26]), .IN2(N165), .S(n176), .Q(n85) );
  MUX21X1 U153 ( .IN1(factor_c[27]), .IN2(N165), .S(n176), .Q(n86) );
  MUX21X1 U154 ( .IN1(factor_c[28]), .IN2(N165), .S(n176), .Q(n87) );
  MUX21X1 U155 ( .IN1(factor_c[29]), .IN2(N165), .S(n176), .Q(n88) );
  INVX0 U156 ( .INP(n177), .ZN(n158) );
  OAI21X1 U157 ( .IN1(case_num[0]), .IN2(n166), .IN3(n158), .QN(n168) );
  AO21X1 U158 ( .IN1(n31), .IN2(factor_d[0]), .IN3(n168), .Q(n32) );
  AO21X1 U159 ( .IN1(n31), .IN2(factor_d[3]), .IN3(n154), .Q(n35) );
  AO22X1 U160 ( .IN1(n31), .IN2(factor_d[6]), .IN3(rst_n), .IN4(N161), .Q(n152) );
  OR2X1 U161 ( .IN1(n154), .IN2(n152), .Q(n38) );
  AND2X1 U162 ( .IN1(n153), .IN2(rst_n), .Q(n155) );
  AO21X1 U163 ( .IN1(n31), .IN2(factor_d[8]), .IN3(n175), .Q(n40) );
  AOI22X1 U164 ( .IN1(n31), .IN2(factor_d[9]), .IN3(n157), .IN4(n3), .QN(n156)
         );
  MUX21X1 U165 ( .IN1(factor_d[10]), .IN2(n174), .S(n176), .Q(n42) );
  AO21X1 U166 ( .IN1(n31), .IN2(factor_d[11]), .IN3(n175), .Q(n43) );
  AOI22X1 U167 ( .IN1(n31), .IN2(factor_d[13]), .IN3(case_num[0]), .IN4(n157), 
        .QN(n159) );
  AOI22X1 U168 ( .IN1(n31), .IN2(factor_d[17]), .IN3(rst_n), .IN4(N157), .QN(
        n162) );
  AO21X1 U169 ( .IN1(n31), .IN2(factor_d[22]), .IN3(n168), .Q(n53) );
  AO221X1 U170 ( .IN1(case_num[1]), .IN2(n1), .IN3(n2), .IN4(n169), .IN5(n4), 
        .Q(n170) );
  MUX21X1 U171 ( .IN1(factor_d[23]), .IN2(n170), .S(n176), .Q(n54) );
  NAND2X0 U172 ( .IN1(case_num[2]), .IN2(n2), .QN(n171) );
  NAND3X0 U173 ( .IN1(n171), .IN2(n1), .IN3(n95), .QN(n172) );
  MUX21X1 U174 ( .IN1(factor_d[24]), .IN2(n172), .S(n176), .Q(n55) );
  AO21X1 U175 ( .IN1(n31), .IN2(factor_d[31]), .IN3(n177), .Q(n61) );
  MUX21X1 U176 ( .IN1(factor_c[2]), .IN2(N154), .S(n176), .Q(n63) );
  AO21X1 U177 ( .IN1(n31), .IN2(factor_c[3]), .IN3(n175), .Q(n64) );
  AO21X1 U178 ( .IN1(n31), .IN2(factor_c[4]), .IN3(n175), .Q(n65) );
  AO21X1 U179 ( .IN1(n31), .IN2(factor_c[6]), .IN3(n177), .Q(n67) );
  AO21X1 U180 ( .IN1(n31), .IN2(factor_c[7]), .IN3(n175), .Q(n68) );
  MUX21X1 U181 ( .IN1(factor_c[9]), .IN2(N154), .S(n176), .Q(n70) );
  AO21X1 U182 ( .IN1(n31), .IN2(factor_c[10]), .IN3(n175), .Q(n71) );
  MUX21X1 U183 ( .IN1(factor_c[16]), .IN2(n174), .S(n176), .Q(n76) );
  AO21X1 U184 ( .IN1(n31), .IN2(factor_c[17]), .IN3(n175), .Q(n77) );
  AO21X1 U185 ( .IN1(n31), .IN2(factor_c[19]), .IN3(n177), .Q(n79) );
  AO21X1 U186 ( .IN1(n31), .IN2(factor_c[21]), .IN3(n175), .Q(n80) );
  AO21X1 U187 ( .IN1(n31), .IN2(factor_c[22]), .IN3(n177), .Q(n81) );
  MUX21X1 U188 ( .IN1(factor_c[23]), .IN2(N162), .S(n176), .Q(n82) );
  AO21X1 U189 ( .IN1(n31), .IN2(factor_c[24]), .IN3(n177), .Q(n83) );
  AO21X1 U190 ( .IN1(n31), .IN2(factor_c[31]), .IN3(n177), .Q(n89) );
endmodule


module add_369 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_370 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_371 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_372 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_373 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_374 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_375 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_376 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_377 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_378 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_379 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_380 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_381 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_382 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_383 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_384 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_385 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_386 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_387 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_388 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_389 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_390 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_391 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_392 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(b), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(b), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module adder24_7 ( clk, rst_n, a, b, cin, out );
  input [23:0] a;
  input [23:0] b;
  output [24:0] out;
  input clk, rst_n, cin;
  wire   c_tmp;
  wire   [24:0] s;
  wire   [22:0] c;

  add_392 add_01 ( .s(s[0]), .a(a[0]), .b(b[0]), .ci(1'b0), .co(c[0]) );
  add_391 add_02 ( .s(s[1]), .a(a[1]), .b(b[1]), .ci(c[0]), .co(c[1]) );
  add_390 add_03 ( .s(s[2]), .a(a[2]), .b(b[2]), .ci(c[1]), .co(c[2]) );
  add_389 add_04 ( .s(s[3]), .a(a[3]), .b(b[3]), .ci(c[2]), .co(c[3]) );
  add_388 add_05 ( .s(s[4]), .a(a[4]), .b(b[4]), .ci(c[3]), .co(c[4]) );
  add_387 add_06 ( .s(s[5]), .a(a[5]), .b(b[5]), .ci(c[4]), .co(c[5]) );
  add_386 add_07 ( .s(s[6]), .a(a[6]), .b(b[6]), .ci(c[5]), .co(c[6]) );
  add_385 add_08 ( .s(s[7]), .a(a[7]), .b(b[7]), .ci(c[6]), .co(c[7]) );
  add_384 add_09 ( .s(s[8]), .a(a[8]), .b(b[8]), .ci(c[7]), .co(c[8]) );
  add_383 add_10 ( .s(s[9]), .a(a[9]), .b(b[9]), .ci(c[8]), .co(c[9]) );
  add_382 add_11 ( .s(s[10]), .a(a[10]), .b(b[10]), .ci(c[9]), .co(c[10]) );
  add_381 add_12 ( .s(s[11]), .a(a[11]), .b(b[11]), .ci(c_tmp), .co(c[11]) );
  add_380 add_13 ( .s(s[12]), .a(a[12]), .b(b[12]), .ci(c[11]), .co(c[12]) );
  add_379 add_14 ( .s(s[13]), .a(a[13]), .b(b[13]), .ci(c[12]), .co(c[13]) );
  add_378 add_15 ( .s(s[14]), .a(a[14]), .b(b[14]), .ci(c[13]), .co(c[14]) );
  add_377 add_16 ( .s(s[15]), .a(a[15]), .b(b[15]), .ci(c[14]), .co(c[15]) );
  add_376 add_17 ( .s(s[16]), .a(a[16]), .b(b[16]), .ci(c[15]), .co(c[16]) );
  add_375 add_18 ( .s(s[17]), .a(a[17]), .b(b[17]), .ci(c[16]), .co(c[17]) );
  add_374 add_19 ( .s(s[18]), .a(a[18]), .b(b[18]), .ci(c[17]), .co(c[18]) );
  add_373 add_20 ( .s(s[19]), .a(a[19]), .b(b[19]), .ci(c[18]), .co(c[19]) );
  add_372 add_21 ( .s(s[20]), .a(a[20]), .b(b[20]), .ci(c[19]), .co(c[20]) );
  add_371 add_22 ( .s(s[21]), .a(a[21]), .b(b[21]), .ci(c[20]), .co(c[21]) );
  add_370 add_23 ( .s(s[22]), .a(a[22]), .b(b[22]), .ci(c[21]), .co(c[22]) );
  add_369 add_24 ( .s(s[23]), .a(a[23]), .b(b[23]), .ci(c[22]), .co(s[24]) );
  DFFARX1 out_reg_10_ ( .D(s[10]), .CLK(clk), .RSTB(rst_n), .Q(out[10]) );
  DFFARX1 out_reg_9_ ( .D(s[9]), .CLK(clk), .RSTB(rst_n), .Q(out[9]) );
  DFFARX1 out_reg_8_ ( .D(s[8]), .CLK(clk), .RSTB(rst_n), .Q(out[8]) );
  DFFARX1 out_reg_7_ ( .D(s[7]), .CLK(clk), .RSTB(rst_n), .Q(out[7]) );
  DFFARX1 out_reg_6_ ( .D(s[6]), .CLK(clk), .RSTB(rst_n), .Q(out[6]) );
  DFFARX1 out_reg_5_ ( .D(s[5]), .CLK(clk), .RSTB(rst_n), .Q(out[5]) );
  DFFARX1 out_reg_4_ ( .D(s[4]), .CLK(clk), .RSTB(rst_n), .Q(out[4]) );
  DFFARX1 out_reg_3_ ( .D(s[3]), .CLK(clk), .RSTB(rst_n), .Q(out[3]) );
  DFFARX1 out_reg_2_ ( .D(s[2]), .CLK(clk), .RSTB(rst_n), .Q(out[2]) );
  DFFARX1 out_reg_1_ ( .D(s[1]), .CLK(clk), .RSTB(rst_n), .Q(out[1]) );
  DFFARX1 out_reg_0_ ( .D(s[0]), .CLK(clk), .RSTB(rst_n), .Q(out[0]) );
  DFFARX1 c_tmp_reg ( .D(c[10]), .CLK(clk), .RSTB(rst_n), .Q(c_tmp) );
  DFFARX1 out_reg_24_ ( .D(s[24]), .CLK(clk), .RSTB(rst_n), .Q(out[24]) );
  DFFARX1 out_reg_23_ ( .D(s[23]), .CLK(clk), .RSTB(rst_n), .Q(out[23]) );
  DFFARX1 out_reg_22_ ( .D(s[22]), .CLK(clk), .RSTB(rst_n), .Q(out[22]) );
  DFFARX1 out_reg_21_ ( .D(s[21]), .CLK(clk), .RSTB(rst_n), .Q(out[21]) );
  DFFARX1 out_reg_20_ ( .D(s[20]), .CLK(clk), .RSTB(rst_n), .Q(out[20]) );
  DFFARX1 out_reg_19_ ( .D(s[19]), .CLK(clk), .RSTB(rst_n), .Q(out[19]) );
  DFFARX1 out_reg_18_ ( .D(s[18]), .CLK(clk), .RSTB(rst_n), .Q(out[18]) );
  DFFARX1 out_reg_17_ ( .D(s[17]), .CLK(clk), .RSTB(rst_n), .Q(out[17]) );
  DFFARX1 out_reg_16_ ( .D(s[16]), .CLK(clk), .RSTB(rst_n), .Q(out[16]) );
  DFFARX1 out_reg_15_ ( .D(s[15]), .CLK(clk), .RSTB(rst_n), .Q(out[15]) );
  DFFARX1 out_reg_14_ ( .D(s[14]), .CLK(clk), .RSTB(rst_n), .Q(out[14]) );
  DFFARX1 out_reg_13_ ( .D(s[13]), .CLK(clk), .RSTB(rst_n), .Q(out[13]) );
  DFFARX1 out_reg_12_ ( .D(s[12]), .CLK(clk), .RSTB(rst_n), .Q(out[12]) );
  DFFARX1 out_reg_11_ ( .D(s[11]), .CLK(clk), .RSTB(rst_n), .Q(out[11]) );
endmodule


module add_393 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_394 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_395 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_396 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_397 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_398 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_399 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_400 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_401 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_402 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_403 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_404 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_405 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_406 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_407 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_408 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_409 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_410 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_411 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_412 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_413 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_414 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_415 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_416 ( s, a, ci, co, b_BAR );
  input a, ci, b_BAR;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(b_BAR), .IN2(n1), .QN(co) );
  INVX0 U2 ( .INP(a), .ZN(n1) );
  MUX21X1 U3 ( .IN1(a), .IN2(n1), .S(b_BAR), .Q(s) );
endmodule


module adder24_8 ( clk, rst_n, a, b, cin, out );
  input [23:0] a;
  input [23:0] b;
  output [24:0] out;
  input clk, rst_n, cin;
  wire   c_tmp, n_1_net_, n_2_net_, n_3_net_, n_4_net_, n_5_net_, n_6_net_,
         n_7_net_, n_8_net_, n_9_net_, n_10_net_, n_11_net_, n_12_net_,
         n_13_net_, n_14_net_, n_15_net_, n_16_net_, n_17_net_, n_18_net_,
         n_19_net_, n_20_net_, n_21_net_, n_22_net_, n_23_net_;
  wire   [24:0] s;
  wire   [23:0] c;

  add_416 add_01 ( .s(s[0]), .a(a[0]), .ci(1'b1), .co(c[0]), .b_BAR(b[0]) );
  add_415 add_02 ( .s(s[1]), .a(a[1]), .b(n_1_net_), .ci(c[0]), .co(c[1]) );
  add_414 add_03 ( .s(s[2]), .a(a[2]), .b(n_2_net_), .ci(c[1]), .co(c[2]) );
  add_413 add_04 ( .s(s[3]), .a(a[3]), .b(n_3_net_), .ci(c[2]), .co(c[3]) );
  add_412 add_05 ( .s(s[4]), .a(a[4]), .b(n_4_net_), .ci(c[3]), .co(c[4]) );
  add_411 add_06 ( .s(s[5]), .a(a[5]), .b(n_5_net_), .ci(c[4]), .co(c[5]) );
  add_410 add_07 ( .s(s[6]), .a(a[6]), .b(n_6_net_), .ci(c[5]), .co(c[6]) );
  add_409 add_08 ( .s(s[7]), .a(a[7]), .b(n_7_net_), .ci(c[6]), .co(c[7]) );
  add_408 add_09 ( .s(s[8]), .a(a[8]), .b(n_8_net_), .ci(c[7]), .co(c[8]) );
  add_407 add_10 ( .s(s[9]), .a(a[9]), .b(n_9_net_), .ci(c[8]), .co(c[9]) );
  add_406 add_11 ( .s(s[10]), .a(a[10]), .b(n_10_net_), .ci(c[9]), .co(c[10])
         );
  add_405 add_12 ( .s(s[11]), .a(a[11]), .b(n_11_net_), .ci(c_tmp), .co(c[11])
         );
  add_404 add_13 ( .s(s[12]), .a(a[12]), .b(n_12_net_), .ci(c[11]), .co(c[12])
         );
  add_403 add_14 ( .s(s[13]), .a(a[13]), .b(n_13_net_), .ci(c[12]), .co(c[13])
         );
  add_402 add_15 ( .s(s[14]), .a(a[14]), .b(n_14_net_), .ci(c[13]), .co(c[14])
         );
  add_401 add_16 ( .s(s[15]), .a(a[15]), .b(n_15_net_), .ci(c[14]), .co(c[15])
         );
  add_400 add_17 ( .s(s[16]), .a(a[16]), .b(n_16_net_), .ci(c[15]), .co(c[16])
         );
  add_399 add_18 ( .s(s[17]), .a(a[17]), .b(n_17_net_), .ci(c[16]), .co(c[17])
         );
  add_398 add_19 ( .s(s[18]), .a(a[18]), .b(n_18_net_), .ci(c[17]), .co(c[18])
         );
  add_397 add_20 ( .s(s[19]), .a(a[19]), .b(n_19_net_), .ci(c[18]), .co(c[19])
         );
  add_396 add_21 ( .s(s[20]), .a(a[20]), .b(n_20_net_), .ci(c[19]), .co(c[20])
         );
  add_395 add_22 ( .s(s[21]), .a(a[21]), .b(n_21_net_), .ci(c[20]), .co(c[21])
         );
  add_394 add_23 ( .s(s[22]), .a(a[22]), .b(n_22_net_), .ci(c[21]), .co(c[22])
         );
  add_393 add_24 ( .s(s[23]), .a(a[23]), .b(n_23_net_), .ci(c[22]), .co(c[23])
         );
  DFFARX1 out_reg_10_ ( .D(s[10]), .CLK(clk), .RSTB(rst_n), .Q(out[10]) );
  DFFARX1 out_reg_9_ ( .D(s[9]), .CLK(clk), .RSTB(rst_n), .Q(out[9]) );
  DFFARX1 out_reg_8_ ( .D(s[8]), .CLK(clk), .RSTB(rst_n), .Q(out[8]) );
  DFFARX1 out_reg_7_ ( .D(s[7]), .CLK(clk), .RSTB(rst_n), .Q(out[7]) );
  DFFARX1 out_reg_6_ ( .D(s[6]), .CLK(clk), .RSTB(rst_n), .Q(out[6]) );
  DFFARX1 out_reg_5_ ( .D(s[5]), .CLK(clk), .RSTB(rst_n), .Q(out[5]) );
  DFFARX1 out_reg_4_ ( .D(s[4]), .CLK(clk), .RSTB(rst_n), .Q(out[4]) );
  DFFARX1 out_reg_3_ ( .D(s[3]), .CLK(clk), .RSTB(rst_n), .Q(out[3]) );
  DFFARX1 out_reg_2_ ( .D(s[2]), .CLK(clk), .RSTB(rst_n), .Q(out[2]) );
  DFFARX1 out_reg_1_ ( .D(s[1]), .CLK(clk), .RSTB(rst_n), .Q(out[1]) );
  DFFARX1 out_reg_0_ ( .D(s[0]), .CLK(clk), .RSTB(rst_n), .Q(out[0]) );
  DFFARX1 c_tmp_reg ( .D(c[10]), .CLK(clk), .RSTB(rst_n), .Q(c_tmp) );
  DFFARX1 out_reg_24_ ( .D(s[24]), .CLK(clk), .RSTB(rst_n), .Q(out[24]) );
  DFFARX1 out_reg_23_ ( .D(s[23]), .CLK(clk), .RSTB(rst_n), .Q(out[23]) );
  DFFARX1 out_reg_22_ ( .D(s[22]), .CLK(clk), .RSTB(rst_n), .Q(out[22]) );
  DFFARX1 out_reg_21_ ( .D(s[21]), .CLK(clk), .RSTB(rst_n), .Q(out[21]) );
  DFFARX1 out_reg_20_ ( .D(s[20]), .CLK(clk), .RSTB(rst_n), .Q(out[20]) );
  DFFARX1 out_reg_19_ ( .D(s[19]), .CLK(clk), .RSTB(rst_n), .Q(out[19]) );
  DFFARX1 out_reg_18_ ( .D(s[18]), .CLK(clk), .RSTB(rst_n), .Q(out[18]) );
  DFFARX1 out_reg_17_ ( .D(s[17]), .CLK(clk), .RSTB(rst_n), .Q(out[17]) );
  DFFARX1 out_reg_16_ ( .D(s[16]), .CLK(clk), .RSTB(rst_n), .Q(out[16]) );
  DFFARX1 out_reg_15_ ( .D(s[15]), .CLK(clk), .RSTB(rst_n), .Q(out[15]) );
  DFFARX1 out_reg_14_ ( .D(s[14]), .CLK(clk), .RSTB(rst_n), .Q(out[14]) );
  DFFARX1 out_reg_13_ ( .D(s[13]), .CLK(clk), .RSTB(rst_n), .Q(out[13]) );
  DFFARX1 out_reg_12_ ( .D(s[12]), .CLK(clk), .RSTB(rst_n), .Q(out[12]) );
  DFFARX1 out_reg_11_ ( .D(s[11]), .CLK(clk), .RSTB(rst_n), .Q(out[11]) );
  INVX0 U3 ( .INP(b[1]), .ZN(n_1_net_) );
  INVX0 U4 ( .INP(b[2]), .ZN(n_2_net_) );
  INVX0 U5 ( .INP(b[3]), .ZN(n_3_net_) );
  INVX0 U6 ( .INP(b[4]), .ZN(n_4_net_) );
  INVX0 U7 ( .INP(b[5]), .ZN(n_5_net_) );
  INVX0 U8 ( .INP(b[6]), .ZN(n_6_net_) );
  INVX0 U9 ( .INP(b[7]), .ZN(n_7_net_) );
  INVX0 U10 ( .INP(b[8]), .ZN(n_8_net_) );
  INVX0 U11 ( .INP(b[9]), .ZN(n_9_net_) );
  INVX0 U12 ( .INP(b[10]), .ZN(n_10_net_) );
  INVX0 U13 ( .INP(c[23]), .ZN(s[24]) );
  INVX0 U14 ( .INP(b[11]), .ZN(n_11_net_) );
  INVX0 U15 ( .INP(b[12]), .ZN(n_12_net_) );
  INVX0 U16 ( .INP(b[13]), .ZN(n_13_net_) );
  INVX0 U17 ( .INP(b[14]), .ZN(n_14_net_) );
  INVX0 U18 ( .INP(b[15]), .ZN(n_15_net_) );
  INVX0 U19 ( .INP(b[16]), .ZN(n_16_net_) );
  INVX0 U20 ( .INP(b[17]), .ZN(n_17_net_) );
  INVX0 U21 ( .INP(b[18]), .ZN(n_18_net_) );
  INVX0 U22 ( .INP(b[19]), .ZN(n_19_net_) );
  INVX0 U23 ( .INP(b[20]), .ZN(n_20_net_) );
  INVX0 U24 ( .INP(b[21]), .ZN(n_21_net_) );
  INVX0 U25 ( .INP(b[22]), .ZN(n_22_net_) );
  INVX0 U26 ( .INP(b[23]), .ZN(n_23_net_) );
endmodule


module add_337 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  XNOR2X1 U1 ( .IN1(ci), .IN2(a), .Q(s) );
endmodule


module add_338 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_339 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_340 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_341 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_342 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_343 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_344 ( s, a, ci, co, b_BAR );
  input a, ci, b_BAR;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(b_BAR), .IN2(n1), .QN(co) );
  INVX0 U2 ( .INP(a), .ZN(n1) );
  MUX21X1 U3 ( .IN1(a), .IN2(n1), .S(b_BAR), .Q(s) );
endmodule


module adder8_25 ( out, a, b, cin );
  output [7:0] out;
  input [7:0] a;
  input [7:0] b;
  input cin;
  wire   n_1_net_, n_2_net_, n_4_net_;
  wire   [6:0] c;

  add_344 add_01 ( .s(out[0]), .a(a[0]), .ci(1'b1), .co(c[0]), .b_BAR(b[0]) );
  add_343 add_02 ( .s(out[1]), .a(a[1]), .b(n_1_net_), .ci(c[0]), .co(c[1]) );
  add_342 add_03 ( .s(out[2]), .a(a[2]), .b(n_2_net_), .ci(c[1]), .co(c[2]) );
  add_341 add_04 ( .s(out[3]), .a(a[3]), .b(1'b1), .ci(c[2]), .co(c[3]) );
  add_340 add_05 ( .s(out[4]), .a(a[4]), .b(n_4_net_), .ci(c[3]), .co(c[4]) );
  add_339 add_06 ( .s(out[5]), .a(a[5]), .b(1'b1), .ci(c[4]), .co(c[5]) );
  add_338 add_07 ( .s(out[6]), .a(a[6]), .b(1'b1), .ci(c[5]), .co(c[6]) );
  add_337 add_08 ( .s(out[7]), .a(a[7]), .b(1'b1), .ci(c[6]) );
  INVX0 U1 ( .INP(b[1]), .ZN(n_1_net_) );
  INVX0 U2 ( .INP(b[2]), .ZN(n_2_net_) );
  INVX0 U3 ( .INP(b[4]), .ZN(n_4_net_) );
endmodule


module add_345 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  XNOR2X1 U1 ( .IN1(ci), .IN2(a), .Q(s) );
endmodule


module add_346 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_347 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_348 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_349 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_350 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_351 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_352 ( s, a, ci, co, b_BAR );
  input a, ci, b_BAR;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(b_BAR), .IN2(n1), .QN(co) );
  INVX0 U2 ( .INP(a), .ZN(n1) );
  MUX21X1 U3 ( .IN1(a), .IN2(n1), .S(b_BAR), .Q(s) );
endmodule


module adder8_26 ( out, a, b, cin );
  output [7:0] out;
  input [7:0] a;
  input [7:0] b;
  input cin;
  wire   n_1_net_, n_2_net_, n_3_net_;
  wire   [6:0] c;

  add_352 add_01 ( .s(out[0]), .a(a[0]), .ci(1'b1), .co(c[0]), .b_BAR(b[0]) );
  add_351 add_02 ( .s(out[1]), .a(a[1]), .b(n_1_net_), .ci(c[0]), .co(c[1]) );
  add_350 add_03 ( .s(out[2]), .a(a[2]), .b(n_2_net_), .ci(c[1]), .co(c[2]) );
  add_349 add_04 ( .s(out[3]), .a(a[3]), .b(n_3_net_), .ci(c[2]), .co(c[3]) );
  add_348 add_05 ( .s(out[4]), .a(a[4]), .b(1'b1), .ci(c[3]), .co(c[4]) );
  add_347 add_06 ( .s(out[5]), .a(a[5]), .b(1'b1), .ci(c[4]), .co(c[5]) );
  add_346 add_07 ( .s(out[6]), .a(a[6]), .b(1'b1), .ci(c[5]), .co(c[6]) );
  add_345 add_08 ( .s(out[7]), .a(a[7]), .b(1'b1), .ci(c[6]) );
  INVX0 U1 ( .INP(b[1]), .ZN(n_1_net_) );
  INVX0 U2 ( .INP(b[2]), .ZN(n_2_net_) );
  INVX0 U3 ( .INP(b[3]), .ZN(n_3_net_) );
endmodule


module add_353 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  XNOR2X1 U1 ( .IN1(ci), .IN2(a), .Q(s) );
endmodule


module add_354 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_355 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_356 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_357 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_358 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_359 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_360 ( s, a, ci, co, b_BAR );
  input a, ci, b_BAR;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(b_BAR), .IN2(n1), .QN(co) );
  INVX0 U2 ( .INP(a), .ZN(n1) );
  MUX21X1 U3 ( .IN1(a), .IN2(n1), .S(b_BAR), .Q(s) );
endmodule


module adder8_27 ( out, a, b, cin );
  output [7:0] out;
  input [7:0] a;
  input [7:0] b;
  input cin;
  wire   n_1_net_, n_2_net_, n_3_net_;
  wire   [6:0] c;

  add_360 add_01 ( .s(out[0]), .a(a[0]), .ci(1'b1), .co(c[0]), .b_BAR(b[0]) );
  add_359 add_02 ( .s(out[1]), .a(a[1]), .b(n_1_net_), .ci(c[0]), .co(c[1]) );
  add_358 add_03 ( .s(out[2]), .a(a[2]), .b(n_2_net_), .ci(c[1]), .co(c[2]) );
  add_357 add_04 ( .s(out[3]), .a(a[3]), .b(n_3_net_), .ci(c[2]), .co(c[3]) );
  add_356 add_05 ( .s(out[4]), .a(a[4]), .b(1'b1), .ci(c[3]), .co(c[4]) );
  add_355 add_06 ( .s(out[5]), .a(a[5]), .b(1'b1), .ci(c[4]), .co(c[5]) );
  add_354 add_07 ( .s(out[6]), .a(a[6]), .b(1'b1), .ci(c[5]), .co(c[6]) );
  add_353 add_08 ( .s(out[7]), .a(a[7]), .b(1'b1), .ci(c[6]) );
  INVX0 U1 ( .INP(b[1]), .ZN(n_1_net_) );
  INVX0 U2 ( .INP(b[2]), .ZN(n_2_net_) );
  INVX0 U3 ( .INP(b[3]), .ZN(n_3_net_) );
endmodule


module add_361 ( s, a, b, co, ci_BAR );
  input a, b, ci_BAR;
  output s, co;


  XNOR2X1 U1 ( .IN1(a), .IN2(ci_BAR), .Q(s) );
endmodule


module add_362 ( s, a, b, ci, co_BAR );
  input a, b, ci;
  output s, co_BAR;


  NAND2X0 U1 ( .IN1(ci), .IN2(a), .QN(co_BAR) );
  OA21X1 U2 ( .IN1(ci), .IN2(a), .IN3(co_BAR), .Q(s) );
endmodule


module add_363 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_364 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_365 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_366 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_367 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_368 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(b), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(b), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module adder8_28 ( out, a, b, cin );
  output [7:0] out;
  input [7:0] a;
  input [7:0] b;
  input cin;

  wire   [6:0] c;

  add_368 add_01 ( .s(out[0]), .a(a[0]), .b(b[0]), .ci(1'b0), .co(c[0]) );
  add_367 add_02 ( .s(out[1]), .a(a[1]), .b(1'b0), .ci(c[0]), .co(c[1]) );
  add_366 add_03 ( .s(out[2]), .a(a[2]), .b(1'b0), .ci(c[1]), .co(c[2]) );
  add_365 add_04 ( .s(out[3]), .a(a[3]), .b(1'b0), .ci(c[2]), .co(c[3]) );
  add_364 add_05 ( .s(out[4]), .a(a[4]), .b(1'b0), .ci(c[3]), .co(c[4]) );
  add_363 add_06 ( .s(out[5]), .a(a[5]), .b(1'b0), .ci(c[4]), .co(c[5]) );
  add_362 add_07 ( .s(out[6]), .a(a[6]), .b(1'b0), .ci(c[5]), .co_BAR(c[6]) );
  add_361 add_08 ( .s(out[7]), .a(a[7]), .b(1'b0), .ci_BAR(c[6]) );
endmodule


module add_417 ( s, a, ci, co, b_BAR );
  input a, ci, b_BAR;
  output s, co;


  XNOR2X1 U1 ( .IN1(ci), .IN2(a), .Q(s) );
endmodule


module add_418 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_419 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_420 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_421 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_422 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_423 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_424 ( s, a, ci, co, b_BAR );
  input a, ci, b_BAR;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(b_BAR), .IN2(n1), .QN(co) );
  INVX0 U2 ( .INP(a), .ZN(n1) );
  MUX21X1 U3 ( .IN1(a), .IN2(n1), .S(b_BAR), .Q(s) );
endmodule


module adder8_29 ( out, a, b, cin );
  output [7:0] out;
  input [7:0] a;
  input [7:0] b;
  input cin;
  wire   n_1_net_, n_2_net_, n_3_net_, n_4_net_, n_5_net_, n_6_net_;
  wire   [6:0] c;

  add_424 add_01 ( .s(out[0]), .a(a[0]), .ci(1'b1), .co(c[0]), .b_BAR(b[0]) );
  add_423 add_02 ( .s(out[1]), .a(a[1]), .b(n_1_net_), .ci(c[0]), .co(c[1]) );
  add_422 add_03 ( .s(out[2]), .a(a[2]), .b(n_2_net_), .ci(c[1]), .co(c[2]) );
  add_421 add_04 ( .s(out[3]), .a(a[3]), .b(n_3_net_), .ci(c[2]), .co(c[3]) );
  add_420 add_05 ( .s(out[4]), .a(a[4]), .b(n_4_net_), .ci(c[3]), .co(c[4]) );
  add_419 add_06 ( .s(out[5]), .a(a[5]), .b(n_5_net_), .ci(c[4]), .co(c[5]) );
  add_418 add_07 ( .s(out[6]), .a(a[6]), .b(n_6_net_), .ci(c[5]), .co(c[6]) );
  add_417 add_08 ( .s(out[7]), .a(a[7]), .ci(c[6]), .b_BAR(1'b0) );
  INVX0 U1 ( .INP(b[4]), .ZN(n_4_net_) );
  INVX0 U2 ( .INP(b[5]), .ZN(n_5_net_) );
  INVX0 U3 ( .INP(b[6]), .ZN(n_6_net_) );
  INVX0 U4 ( .INP(b[1]), .ZN(n_1_net_) );
  INVX0 U5 ( .INP(b[2]), .ZN(n_2_net_) );
  INVX0 U6 ( .INP(b[3]), .ZN(n_3_net_) );
endmodule


module add_425 ( s, a, ci, co, b_BAR );
  input a, ci, b_BAR;
  output s, co;


  XNOR2X1 U1 ( .IN1(b_BAR), .IN2(ci), .Q(s) );
endmodule


module add_426 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_427 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_428 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_429 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_430 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_431 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_432 ( s, a, ci, co, b_BAR );
  input a, ci, b_BAR;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(b_BAR), .IN2(n1), .QN(co) );
  INVX0 U2 ( .INP(a), .ZN(n1) );
  MUX21X1 U3 ( .IN1(a), .IN2(n1), .S(b_BAR), .Q(s) );
endmodule


module adder8_30 ( out, a, b, cin );
  output [7:0] out;
  input [7:0] a;
  input [7:0] b;
  input cin;
  wire   n_1_net_, n_2_net_, n_3_net_, n_4_net_, n_5_net_, n_6_net_;
  wire   [6:0] c;

  add_432 add_01 ( .s(out[0]), .a(a[0]), .ci(1'b1), .co(c[0]), .b_BAR(b[0]) );
  add_431 add_02 ( .s(out[1]), .a(a[1]), .b(n_1_net_), .ci(c[0]), .co(c[1]) );
  add_430 add_03 ( .s(out[2]), .a(a[2]), .b(n_2_net_), .ci(c[1]), .co(c[2]) );
  add_429 add_04 ( .s(out[3]), .a(a[3]), .b(n_3_net_), .ci(c[2]), .co(c[3]) );
  add_428 add_05 ( .s(out[4]), .a(a[4]), .b(n_4_net_), .ci(c[3]), .co(c[4]) );
  add_427 add_06 ( .s(out[5]), .a(a[5]), .b(n_5_net_), .ci(c[4]), .co(c[5]) );
  add_426 add_07 ( .s(out[6]), .a(a[6]), .b(n_6_net_), .ci(c[5]), .co(c[6]) );
  add_425 add_08 ( .s(out[7]), .a(1'b0), .ci(c[6]), .b_BAR(b[7]) );
  INVX0 U1 ( .INP(b[4]), .ZN(n_4_net_) );
  INVX0 U2 ( .INP(b[5]), .ZN(n_5_net_) );
  INVX0 U3 ( .INP(b[6]), .ZN(n_6_net_) );
  INVX0 U4 ( .INP(b[1]), .ZN(n_1_net_) );
  INVX0 U5 ( .INP(b[2]), .ZN(n_2_net_) );
  INVX0 U6 ( .INP(b[3]), .ZN(n_3_net_) );
endmodule


module floating_point_adder_4 ( clk, rst_n, input_factor_01, input_factor_02, 
        output_adder );
  input [31:0] input_factor_01;
  input [31:0] input_factor_02;
  output [31:0] output_adder;
  input clk, rst_n;
  wire   N34, N35, N36, N37, N38, N39, N40, N41, N152, N153, N154, N155, N156,
         N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, N167,
         N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178,
         N179, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189,
         N190, N191, N192, N193, N194, N195, N196, N197, N198,
         add_sub_result_24_, N211, shift_temp_01_0_, N226, N227, N228, N229,
         N230, N231, N232, N233, N234, N235, N236, N237, N238, N239, N240,
         N241, N242, N243, N244, N245, N246, N247, N248, N256, N257, N258,
         N260, N261, N262, N263, N264, N265, N266, N267, N268, N269, N270,
         N271, N272, N273, N274, N275, N276, N277, N278, N279, N280, N281,
         N306, N307, N308, N346, N347, N348, N349, N350, N351, N352, N353,
         N354, N355, N380, N381, N382, N383, N384, N385, N386, N387, N388,
         N389, N390, N391, N392, N393, N394, N395, N396, N397, N398, N399,
         N400, N401, N402, N403, N404, N405, N406, N407, N408, N409, N410, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861;
  wire   [7:0] exp_diff_value;
  wire   [7:0] exponent_factor_21;
  wire   [7:0] exponent_factor_12;
  wire   [23:0] shift_smaller_factor;
  wire   [22:0] larger_factor;
  wire   [7:0] larger_exponent;
  wire   [24:0] add_result;
  wire   [24:0] sub_result;
  wire   [22:0] pre_sig_res_01;
  wire   [3:0] shift_temp_02;
  wire   [22:1] pre_sig_res_02;
  wire   [2:0] shift_temp_03;
  wire   [22:9] pre_sig_res_03;
  wire   [4:0] shift_temp_04;
  wire   [22:16] pre_sig_res_04;
  wire   [7:0] add_output_exponent_w1;
  wire   [7:0] add_output_exponent_w2;
  wire   [7:0] add_output_exponent_w3;
  wire   [7:0] add_output_exponent_w4;

  adder8_30 adder8_01 ( .out(exponent_factor_21), .a({1'b0, 
        input_factor_02[29:23]}), .b(input_factor_01[30:23]), .cin(1'b1) );
  adder8_29 adder8_02 ( .out(exponent_factor_12), .a(input_factor_01[30:23]), 
        .b({1'b0, input_factor_02[29:23]}), .cin(1'b1) );
  adder24_8 adder24_01 ( .clk(clk), .rst_n(rst_n), .a({shift_temp_04[4], 
        larger_factor}), .b(shift_smaller_factor), .cin(1'b1), .out(sub_result) );
  adder24_7 adder24_02 ( .clk(clk), .rst_n(rst_n), .a({shift_temp_04[4], 
        larger_factor}), .b(shift_smaller_factor), .cin(1'b0), .out(add_result) );
  adder8_28 adder8_03 ( .out(add_output_exponent_w1), .a(larger_exponent), .b(
        {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, shift_temp_01_0_}), .cin(
        1'b0) );
  adder8_27 adder8_04 ( .out(add_output_exponent_w2), .a(larger_exponent), .b(
        {1'b0, 1'b0, 1'b0, 1'b0, shift_temp_02}), .cin(1'b1) );
  adder8_26 adder8_05 ( .out(add_output_exponent_w3), .a(larger_exponent), .b(
        {1'b0, 1'b0, 1'b0, 1'b0, shift_temp_04[4], shift_temp_03}), .cin(1'b1)
         );
  adder8_25 adder8_06 ( .out(add_output_exponent_w4), .a(larger_exponent), .b(
        {1'b0, 1'b0, 1'b0, shift_temp_04[4], 1'b0, shift_temp_04[2:0]}), .cin(
        1'b1) );
  DFFARX1 exp_diff_value_reg_7_ ( .D(N41), .CLK(clk), .RSTB(rst_n), .Q(
        exp_diff_value[7]) );
  DFFARX1 exp_diff_value_reg_6_ ( .D(N40), .CLK(clk), .RSTB(rst_n), .Q(
        exp_diff_value[6]) );
  DFFARX1 exp_diff_value_reg_5_ ( .D(N39), .CLK(clk), .RSTB(rst_n), .Q(
        exp_diff_value[5]) );
  DFFARX1 exp_diff_value_reg_4_ ( .D(N38), .CLK(clk), .RSTB(rst_n), .Q(
        exp_diff_value[4]) );
  DFFARX1 exp_diff_value_reg_3_ ( .D(N37), .CLK(clk), .RSTB(rst_n), .Q(
        exp_diff_value[3]), .QN(n2) );
  DFFARX1 exp_diff_value_reg_2_ ( .D(N36), .CLK(clk), .RSTB(rst_n), .Q(
        exp_diff_value[2]), .QN(n1) );
  DFFARX1 exp_diff_value_reg_1_ ( .D(N35), .CLK(clk), .RSTB(rst_n), .Q(
        exp_diff_value[1]), .QN(n6) );
  DFFARX1 exp_diff_value_reg_0_ ( .D(N34), .CLK(clk), .RSTB(rst_n), .Q(
        exp_diff_value[0]), .QN(n3) );
  DFFARX1 larger_factor_reg_22_ ( .D(N198), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[22]) );
  DFFARX1 larger_factor_reg_21_ ( .D(N197), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[21]) );
  DFFARX1 larger_factor_reg_20_ ( .D(N196), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[20]) );
  DFFARX1 larger_factor_reg_19_ ( .D(N195), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[19]) );
  DFFARX1 larger_factor_reg_18_ ( .D(N194), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[18]) );
  DFFARX1 larger_factor_reg_17_ ( .D(N193), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[17]) );
  DFFARX1 larger_factor_reg_16_ ( .D(N192), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[16]) );
  DFFARX1 larger_factor_reg_15_ ( .D(N191), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[15]) );
  DFFARX1 larger_factor_reg_14_ ( .D(N190), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[14]) );
  DFFARX1 larger_factor_reg_13_ ( .D(N189), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[13]) );
  DFFARX1 larger_factor_reg_12_ ( .D(N188), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[12]) );
  DFFARX1 larger_factor_reg_11_ ( .D(N187), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[11]) );
  DFFARX1 larger_factor_reg_10_ ( .D(N186), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[10]) );
  DFFARX1 larger_factor_reg_9_ ( .D(N185), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[9]) );
  DFFARX1 larger_factor_reg_8_ ( .D(N184), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[8]) );
  DFFARX1 larger_factor_reg_7_ ( .D(N183), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[7]) );
  DFFARX1 larger_factor_reg_6_ ( .D(N182), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[6]) );
  DFFARX1 larger_factor_reg_5_ ( .D(N181), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[5]) );
  DFFARX1 larger_factor_reg_4_ ( .D(N180), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[4]) );
  DFFARX1 larger_factor_reg_3_ ( .D(N179), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[3]) );
  DFFARX1 larger_factor_reg_2_ ( .D(N178), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[2]) );
  DFFARX1 larger_factor_reg_1_ ( .D(N177), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[1]) );
  DFFARX1 larger_factor_reg_0_ ( .D(N176), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[0]) );
  DFFARX1 shift_smaller_factor_reg_23_ ( .D(N175), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[23]) );
  DFFARX1 shift_smaller_factor_reg_22_ ( .D(N174), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[22]) );
  DFFARX1 shift_smaller_factor_reg_21_ ( .D(N173), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[21]) );
  DFFARX1 shift_smaller_factor_reg_20_ ( .D(N172), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[20]) );
  DFFARX1 shift_smaller_factor_reg_19_ ( .D(N171), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[19]) );
  DFFARX1 shift_smaller_factor_reg_18_ ( .D(N170), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[18]) );
  DFFARX1 shift_smaller_factor_reg_17_ ( .D(N169), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[17]) );
  DFFARX1 shift_smaller_factor_reg_16_ ( .D(N168), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[16]) );
  DFFARX1 shift_smaller_factor_reg_15_ ( .D(N167), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[15]) );
  DFFARX1 shift_smaller_factor_reg_14_ ( .D(N166), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[14]) );
  DFFARX1 shift_smaller_factor_reg_13_ ( .D(N165), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[13]) );
  DFFARX1 shift_smaller_factor_reg_12_ ( .D(N164), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[12]) );
  DFFARX1 shift_smaller_factor_reg_11_ ( .D(N163), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[11]) );
  DFFARX1 shift_smaller_factor_reg_10_ ( .D(N162), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[10]) );
  DFFARX1 shift_smaller_factor_reg_9_ ( .D(N161), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[9]) );
  DFFARX1 shift_smaller_factor_reg_8_ ( .D(N160), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[8]) );
  DFFARX1 shift_smaller_factor_reg_7_ ( .D(N159), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[7]) );
  DFFARX1 shift_smaller_factor_reg_6_ ( .D(N158), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[6]) );
  DFFARX1 shift_smaller_factor_reg_5_ ( .D(N157), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[5]) );
  DFFARX1 shift_smaller_factor_reg_4_ ( .D(N156), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[4]) );
  DFFARX1 shift_smaller_factor_reg_3_ ( .D(N155), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[3]) );
  DFFARX1 shift_smaller_factor_reg_2_ ( .D(N154), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[2]) );
  DFFARX1 shift_smaller_factor_reg_1_ ( .D(N153), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[1]) );
  DFFARX1 shift_smaller_factor_reg_0_ ( .D(N152), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[0]) );
  DFFX1 larger_exponent_reg_7_ ( .D(n839), .CLK(clk), .Q(larger_exponent[7])
         );
  DFFX1 larger_exponent_reg_6_ ( .D(n840), .CLK(clk), .Q(larger_exponent[6])
         );
  DFFX1 larger_exponent_reg_5_ ( .D(n841), .CLK(clk), .Q(larger_exponent[5])
         );
  DFFX1 larger_exponent_reg_4_ ( .D(n842), .CLK(clk), .Q(larger_exponent[4])
         );
  DFFX1 larger_exponent_reg_3_ ( .D(n843), .CLK(clk), .Q(larger_exponent[3])
         );
  DFFX1 larger_exponent_reg_2_ ( .D(n844), .CLK(clk), .Q(larger_exponent[2])
         );
  DFFX1 larger_exponent_reg_1_ ( .D(n845), .CLK(clk), .Q(larger_exponent[1])
         );
  DFFX1 larger_exponent_reg_0_ ( .D(n846), .CLK(clk), .Q(larger_exponent[0])
         );
  DFFARX1 shift_temp_04_reg_4_ ( .D(1'b1), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_04[4]) );
  DFFARX1 shift_temp_01_reg_0_ ( .D(add_sub_result_24_), .CLK(clk), .RSTB(
        rst_n), .Q(shift_temp_01_0_) );
  DFFARX1 pre_sig_res_02_reg_1_ ( .D(N260), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[1]) );
  DFFARX1 pre_sig_res_02_reg_2_ ( .D(N261), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[2]) );
  DFFARX1 pre_sig_res_02_reg_3_ ( .D(N262), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[3]) );
  DFFARX1 pre_sig_res_02_reg_4_ ( .D(N263), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[4]) );
  DFFARX1 pre_sig_res_02_reg_5_ ( .D(N264), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[5]) );
  DFFARX1 pre_sig_res_02_reg_6_ ( .D(N265), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[6]) );
  DFFARX1 pre_sig_res_02_reg_7_ ( .D(N266), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[7]) );
  DFFARX1 shift_temp_02_reg_2_ ( .D(N258), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_02[2]) );
  DFFASX1 shift_temp_02_reg_3_ ( .D(n838), .CLK(clk), .SETB(rst_n), .QN(
        shift_temp_02[3]) );
  DFFARX1 pre_sig_res_02_reg_8_ ( .D(N267), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[8]) );
  DFFARX1 pre_sig_res_02_reg_9_ ( .D(N268), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[9]) );
  DFFARX1 pre_sig_res_02_reg_10_ ( .D(N269), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[10]) );
  DFFARX1 pre_sig_res_02_reg_11_ ( .D(N270), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[11]) );
  DFFARX1 pre_sig_res_02_reg_12_ ( .D(N271), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[12]) );
  DFFARX1 pre_sig_res_02_reg_13_ ( .D(N272), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[13]) );
  DFFARX1 pre_sig_res_02_reg_14_ ( .D(N273), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[14]) );
  DFFARX1 pre_sig_res_02_reg_15_ ( .D(N274), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[15]) );
  DFFARX1 pre_sig_res_02_reg_16_ ( .D(N275), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[16]) );
  DFFARX1 pre_sig_res_02_reg_17_ ( .D(N276), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[17]) );
  DFFARX1 pre_sig_res_02_reg_18_ ( .D(N277), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[18]) );
  DFFARX1 pre_sig_res_02_reg_19_ ( .D(N278), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[19]) );
  DFFARX1 pre_sig_res_02_reg_20_ ( .D(N279), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[20]) );
  DFFARX1 pre_sig_res_02_reg_21_ ( .D(N280), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[21]) );
  DFFARX1 pre_sig_res_02_reg_22_ ( .D(N281), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[22]) );
  DFFARX1 shift_temp_02_reg_1_ ( .D(N257), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_02[1]) );
  DFFARX1 shift_temp_02_reg_0_ ( .D(N256), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_02[0]) );
  DFFX1 pre_sig_res_03_reg_9_ ( .D(n847), .CLK(clk), .Q(pre_sig_res_03[9]) );
  DFFX1 pre_sig_res_03_reg_10_ ( .D(n848), .CLK(clk), .Q(pre_sig_res_03[10])
         );
  DFFX1 pre_sig_res_03_reg_12_ ( .D(n849), .CLK(clk), .Q(pre_sig_res_03[12])
         );
  DFFX1 pre_sig_res_03_reg_11_ ( .D(n850), .CLK(clk), .Q(pre_sig_res_03[11])
         );
  DFFX1 pre_sig_res_03_reg_13_ ( .D(n851), .CLK(clk), .Q(pre_sig_res_03[13])
         );
  DFFX1 pre_sig_res_03_reg_14_ ( .D(n852), .CLK(clk), .Q(pre_sig_res_03[14])
         );
  DFFARX1 shift_temp_03_reg_2_ ( .D(N308), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_03[2]) );
  DFFARX1 shift_temp_03_reg_0_ ( .D(N306), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_03[0]) );
  DFFARX1 shift_temp_03_reg_1_ ( .D(N307), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_03[1]) );
  DFFX1 pre_sig_res_03_reg_15_ ( .D(n853), .CLK(clk), .Q(pre_sig_res_03[15])
         );
  DFFX1 pre_sig_res_03_reg_16_ ( .D(n854), .CLK(clk), .Q(pre_sig_res_03[16])
         );
  DFFX1 pre_sig_res_03_reg_17_ ( .D(n855), .CLK(clk), .Q(pre_sig_res_03[17])
         );
  DFFX1 pre_sig_res_03_reg_18_ ( .D(n856), .CLK(clk), .Q(pre_sig_res_03[18])
         );
  DFFX1 pre_sig_res_03_reg_19_ ( .D(n857), .CLK(clk), .Q(pre_sig_res_03[19])
         );
  DFFX1 pre_sig_res_03_reg_20_ ( .D(n858), .CLK(clk), .Q(pre_sig_res_03[20])
         );
  DFFX1 pre_sig_res_03_reg_21_ ( .D(n859), .CLK(clk), .Q(pre_sig_res_03[21])
         );
  DFFX1 pre_sig_res_03_reg_22_ ( .D(n860), .CLK(clk), .Q(pre_sig_res_03[22])
         );
  DFFARX1 pre_sig_res_04_reg_16_ ( .D(N349), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_04[16]) );
  DFFARX1 pre_sig_res_04_reg_17_ ( .D(N350), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_04[17]) );
  DFFARX1 pre_sig_res_04_reg_18_ ( .D(N351), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_04[18]) );
  DFFARX1 pre_sig_res_04_reg_19_ ( .D(N352), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_04[19]) );
  DFFARX1 pre_sig_res_04_reg_20_ ( .D(N353), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_04[20]) );
  DFFARX1 pre_sig_res_04_reg_21_ ( .D(N354), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_04[21]) );
  DFFARX1 pre_sig_res_04_reg_22_ ( .D(N355), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_04[22]) );
  DFFARX1 add_output_sign_reg ( .D(N211), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[31]) );
  DFFARX1 pre_sig_res_01_reg_0_ ( .D(N226), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[0]) );
  DFFARX1 pre_sig_res_01_reg_1_ ( .D(N227), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[1]) );
  DFFARX1 pre_sig_res_01_reg_2_ ( .D(N228), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[2]) );
  DFFARX1 pre_sig_res_01_reg_3_ ( .D(N229), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[3]) );
  DFFARX1 pre_sig_res_01_reg_4_ ( .D(N230), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[4]) );
  DFFARX1 pre_sig_res_01_reg_5_ ( .D(N231), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[5]) );
  DFFARX1 pre_sig_res_01_reg_6_ ( .D(N232), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[6]) );
  DFFARX1 pre_sig_res_01_reg_7_ ( .D(N233), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[7]) );
  DFFARX1 pre_sig_res_01_reg_8_ ( .D(N234), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[8]) );
  DFFARX1 pre_sig_res_01_reg_9_ ( .D(N235), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[9]) );
  DFFARX1 pre_sig_res_01_reg_10_ ( .D(N236), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[10]) );
  DFFARX1 pre_sig_res_01_reg_11_ ( .D(N237), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[11]) );
  DFFARX1 pre_sig_res_01_reg_12_ ( .D(N238), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[12]) );
  DFFARX1 pre_sig_res_01_reg_13_ ( .D(N239), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[13]) );
  DFFARX1 pre_sig_res_01_reg_14_ ( .D(N240), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[14]) );
  DFFARX1 pre_sig_res_01_reg_15_ ( .D(N241), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[15]) );
  DFFARX1 pre_sig_res_01_reg_16_ ( .D(N242), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[16]) );
  DFFARX1 pre_sig_res_01_reg_17_ ( .D(N243), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[17]) );
  DFFARX1 pre_sig_res_01_reg_18_ ( .D(N244), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[18]) );
  DFFARX1 pre_sig_res_01_reg_19_ ( .D(N245), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[19]) );
  DFFARX1 pre_sig_res_01_reg_20_ ( .D(N246), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[20]) );
  DFFARX1 pre_sig_res_01_reg_21_ ( .D(N247), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[21]) );
  DFFARX1 pre_sig_res_01_reg_22_ ( .D(N248), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[22]) );
  DFFARX1 shift_temp_04_reg_2_ ( .D(N348), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_04[2]) );
  DFFARX1 shift_temp_04_reg_1_ ( .D(N347), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_04[1]) );
  DFFARX1 shift_temp_04_reg_0_ ( .D(N346), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_04[0]) );
  DFFARX1 add_output_exponent_reg_7_ ( .D(N387), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[30]) );
  DFFARX1 add_output_exponent_reg_6_ ( .D(N386), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[29]) );
  DFFARX1 add_output_exponent_reg_5_ ( .D(N385), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[28]) );
  DFFARX1 add_output_exponent_reg_4_ ( .D(N384), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[27]) );
  DFFARX1 add_output_exponent_reg_3_ ( .D(N383), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[26]) );
  DFFARX1 add_output_exponent_reg_2_ ( .D(N382), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[25]) );
  DFFARX1 add_output_exponent_reg_1_ ( .D(N381), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[24]) );
  DFFARX1 add_output_exponent_reg_0_ ( .D(N380), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[23]) );
  DFFARX1 add_output_significands_reg_22_ ( .D(N410), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[22]) );
  DFFARX1 add_output_significands_reg_21_ ( .D(N409), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[21]) );
  DFFARX1 add_output_significands_reg_20_ ( .D(N408), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[20]) );
  DFFARX1 add_output_significands_reg_19_ ( .D(N407), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[19]) );
  DFFARX1 add_output_significands_reg_18_ ( .D(N406), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[18]) );
  DFFARX1 add_output_significands_reg_17_ ( .D(N405), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[17]) );
  DFFARX1 add_output_significands_reg_16_ ( .D(N404), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[16]) );
  DFFARX1 add_output_significands_reg_15_ ( .D(N403), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[15]) );
  DFFARX1 add_output_significands_reg_14_ ( .D(N402), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[14]) );
  DFFARX1 add_output_significands_reg_13_ ( .D(N401), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[13]) );
  DFFARX1 add_output_significands_reg_12_ ( .D(N400), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[12]) );
  DFFARX1 add_output_significands_reg_11_ ( .D(N399), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[11]) );
  DFFARX1 add_output_significands_reg_10_ ( .D(N398), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[10]) );
  DFFARX1 add_output_significands_reg_9_ ( .D(N397), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[9]) );
  DFFARX1 add_output_significands_reg_8_ ( .D(N396), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[8]) );
  DFFARX1 add_output_significands_reg_7_ ( .D(N395), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[7]) );
  DFFARX1 add_output_significands_reg_6_ ( .D(N394), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[6]) );
  DFFARX1 add_output_significands_reg_5_ ( .D(N393), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[5]) );
  DFFARX1 add_output_significands_reg_4_ ( .D(N392), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[4]) );
  DFFARX1 add_output_significands_reg_3_ ( .D(N391), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[3]) );
  DFFARX1 add_output_significands_reg_2_ ( .D(N390), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[2]) );
  DFFARX1 add_output_significands_reg_1_ ( .D(N389), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[1]) );
  DFFARX1 add_output_significands_reg_0_ ( .D(N388), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[0]) );
  INVX1 U5 ( .INP(rst_n), .ZN(n861) );
  NAND2X0 U3 ( .IN1(input_factor_02[13]), .IN2(n665), .QN(n58) );
  NAND2X0 U4 ( .IN1(n484), .IN2(n397), .QN(n564) );
  NAND2X0 U6 ( .IN1(input_factor_02[24]), .IN2(n548), .QN(n32) );
  NAND2X0 U7 ( .IN1(input_factor_01[27]), .IN2(n590), .QN(n28) );
  NAND2X0 U8 ( .IN1(input_factor_01[26]), .IN2(n584), .QN(n29) );
  NAND2X0 U9 ( .IN1(input_factor_01[28]), .IN2(n596), .QN(n39) );
  NAND2X0 U10 ( .IN1(input_factor_02[28]), .IN2(n595), .QN(n43) );
  NAND2X0 U11 ( .IN1(n818), .IN2(n524), .QN(n382) );
  NAND2X0 U12 ( .IN1(n788), .IN2(n516), .QN(n381) );
  NAND2X0 U13 ( .IN1(n781), .IN2(n517), .QN(n380) );
  NAND2X0 U14 ( .IN1(n757), .IN2(n731), .QN(n561) );
  NAND2X0 U15 ( .IN1(n401), .IN2(n494), .QN(n378) );
  NAND2X0 U16 ( .IN1(n492), .IN2(n404), .QN(n377) );
  NAND2X0 U17 ( .IN1(n376), .IN2(n570), .QN(n403) );
  NAND2X0 U18 ( .IN1(n80), .IN2(n79), .QN(n219) );
  NAND2X0 U19 ( .IN1(n90), .IN2(n89), .QN(n218) );
  NAND2X0 U20 ( .IN1(n131), .IN2(n130), .QN(n236) );
  NAND2X0 U21 ( .IN1(n142), .IN2(n141), .QN(n235) );
  NAND2X0 U22 ( .IN1(n159), .IN2(n158), .QN(n252) );
  NAND2X0 U23 ( .IN1(n169), .IN2(n168), .QN(n251) );
  NAND2X0 U24 ( .IN1(n716), .IN2(n273), .QN(n254) );
  NAND2X0 U25 ( .IN1(n273), .IN2(n834), .QN(n253) );
  NAND2X0 U26 ( .IN1(n188), .IN2(n187), .QN(n272) );
  NAND2X0 U27 ( .IN1(n198), .IN2(n197), .QN(n271) );
  NAND2X0 U28 ( .IN1(exp_diff_value[0]), .IN2(n6), .QN(n200) );
  NAND2X0 U29 ( .IN1(exp_diff_value[1]), .IN2(exp_diff_value[0]), .QN(n199) );
  NAND2X0 U30 ( .IN1(n84), .IN2(n83), .QN(n215) );
  NAND2X0 U31 ( .IN1(n135), .IN2(n134), .QN(n232) );
  NAND2X0 U32 ( .IN1(n163), .IN2(n162), .QN(n248) );
  NAND2X0 U33 ( .IN1(n202), .IN2(n201), .QN(n265) );
  NAND2X0 U34 ( .IN1(n192), .IN2(n191), .QN(n268) );
  NAND2X0 U35 ( .IN1(n68), .IN2(n69), .QN(n12) );
  NAND2X0 U36 ( .IN1(input_factor_02[16]), .IN2(n328), .QN(n68) );
  NAND2X0 U37 ( .IN1(input_factor_01[23]), .IN2(n559), .QN(n30) );
  NAND2X0 U38 ( .IN1(n549), .IN2(input_factor_02[25]), .QN(n31) );
  NAND2X0 U39 ( .IN1(input_factor_02[27]), .IN2(n589), .QN(n22) );
  NAND2X0 U40 ( .IN1(input_factor_02[26]), .IN2(n583), .QN(n20) );
  NAND2X0 U41 ( .IN1(n375), .IN2(n72), .QN(n220) );
  NAND2X0 U42 ( .IN1(n723), .IN2(pre_sig_res_01[9]), .QN(n645) );
  NAND2X0 U43 ( .IN1(n723), .IN2(pre_sig_res_01[10]), .QN(n651) );
  NAND2X0 U44 ( .IN1(n723), .IN2(pre_sig_res_01[11]), .QN(n657) );
  NAND2X0 U45 ( .IN1(n723), .IN2(pre_sig_res_01[12]), .QN(n663) );
  NAND2X0 U46 ( .IN1(n723), .IN2(pre_sig_res_01[13]), .QN(n669) );
  NAND2X0 U47 ( .IN1(n723), .IN2(pre_sig_res_01[15]), .QN(n678) );
  NAND2X0 U48 ( .IN1(n723), .IN2(pre_sig_res_01[16]), .QN(n682) );
  NAND2X0 U49 ( .IN1(n723), .IN2(pre_sig_res_01[17]), .QN(n688) );
  NAND2X0 U50 ( .IN1(n723), .IN2(pre_sig_res_01[18]), .QN(n694) );
  NAND2X0 U51 ( .IN1(n723), .IN2(pre_sig_res_01[19]), .QN(n700) );
  NAND2X0 U52 ( .IN1(n723), .IN2(pre_sig_res_01[20]), .QN(n706) );
  NAND2X0 U53 ( .IN1(n723), .IN2(pre_sig_res_01[21]), .QN(n712) );
  NAND2X0 U54 ( .IN1(n723), .IN2(pre_sig_res_01[22]), .QN(n724) );
  NAND2X0 U55 ( .IN1(n723), .IN2(add_output_exponent_w1[0]), .QN(n571) );
  NAND2X0 U56 ( .IN1(n723), .IN2(add_output_exponent_w1[1]), .QN(n575) );
  NAND2X0 U57 ( .IN1(n723), .IN2(add_output_exponent_w1[2]), .QN(n579) );
  NAND2X0 U58 ( .IN1(n723), .IN2(add_output_exponent_w1[3]), .QN(n585) );
  NAND2X0 U59 ( .IN1(n723), .IN2(add_output_exponent_w1[4]), .QN(n591) );
  NAND2X0 U60 ( .IN1(n723), .IN2(add_output_exponent_w1[5]), .QN(n597) );
  NAND2X0 U61 ( .IN1(n557), .IN2(n556), .QN(n718) );
  NAND2X0 U62 ( .IN1(n723), .IN2(add_output_exponent_w1[6]), .QN(n603) );
  NAND2X0 U63 ( .IN1(n518), .IN2(n828), .QN(n536) );
  NAND2X0 U64 ( .IN1(n515), .IN2(n524), .QN(n521) );
  NAND2X0 U65 ( .IN1(n220), .IN2(n361), .QN(n393) );
  NAND2X0 U66 ( .IN1(n516), .IN2(n801), .QN(n534) );
  NAND2X0 U67 ( .IN1(n517), .IN2(n768), .QN(n535) );
  NAND2X0 U68 ( .IN1(n773), .IN2(n757), .QN(n732) );
  NAND2X0 U69 ( .IN1(n731), .IN2(n744), .QN(n806) );
  NAND2X0 U70 ( .IN1(n514), .IN2(n502), .QN(n735) );
  NAND2X0 U71 ( .IN1(n514), .IN2(n506), .QN(n728) );
  NAND2X0 U72 ( .IN1(n397), .IN2(n396), .QN(n496) );
  NAND2X0 U73 ( .IN1(n414), .IN2(n830), .QN(n411) );
  NAND2X0 U74 ( .IN1(n401), .IN2(n398), .QN(n485) );
  NAND2X0 U75 ( .IN1(n404), .IN2(n399), .QN(n489) );
  NAND2X0 U76 ( .IN1(n400), .IN2(n570), .QN(n487) );
  NAND2X0 U77 ( .IN1(n77), .IN2(n76), .QN(n85) );
  NAND2X0 U78 ( .IN1(n88), .IN2(n87), .QN(n93) );
  NAND2X0 U79 ( .IN1(input_factor_02[0]), .IN2(n184), .QN(n119) );
  NAND2X0 U80 ( .IN1(n129), .IN2(n128), .QN(n136) );
  NAND2X0 U81 ( .IN1(n140), .IN2(n139), .QN(n145) );
  NAND2X0 U82 ( .IN1(input_factor_02[1]), .IN2(n184), .QN(n149) );
  NAND2X0 U83 ( .IN1(n157), .IN2(n156), .QN(n164) );
  NAND2X0 U84 ( .IN1(n167), .IN2(n166), .QN(n172) );
  NAND2X0 U85 ( .IN1(input_factor_02[2]), .IN2(n184), .QN(n176) );
  NAND2X0 U86 ( .IN1(n273), .IN2(n2), .QN(n182) );
  NAND2X0 U87 ( .IN1(n186), .IN2(n185), .QN(n193) );
  NAND2X0 U88 ( .IN1(n196), .IN2(n195), .QN(n203) );
  NAND2X0 U89 ( .IN1(input_factor_02[3]), .IN2(n184), .QN(n207) );
  NAND2X0 U90 ( .IN1(n92), .IN2(n91), .QN(n211) );
  NAND2X0 U91 ( .IN1(n82), .IN2(n81), .QN(n210) );
  NAND2X0 U92 ( .IN1(n133), .IN2(n132), .QN(n227) );
  NAND2X0 U93 ( .IN1(n144), .IN2(n143), .QN(n228) );
  NAND2X0 U94 ( .IN1(n161), .IN2(n160), .QN(n243) );
  NAND2X0 U95 ( .IN1(n171), .IN2(n170), .QN(n244) );
  NAND2X0 U96 ( .IN1(n190), .IN2(n189), .QN(n261) );
  NAND2X0 U97 ( .IN1(exp_diff_value[3]), .IN2(n353), .QN(n327) );
  NAND2X0 U98 ( .IN1(exp_diff_value[3]), .IN2(n351), .QN(n326) );
  NAND2X0 U99 ( .IN1(n327), .IN2(n326), .QN(n329) );
  NAND2X0 U100 ( .IN1(n2), .IN2(n353), .QN(n347) );
  NAND2X0 U101 ( .IN1(n2), .IN2(n351), .QN(n345) );
  NAND2X0 U102 ( .IN1(n364), .IN2(n74), .QN(n361) );
  NAND2X0 U103 ( .IN1(n353), .IN2(n352), .QN(n365) );
  NAND2X0 U104 ( .IN1(n352), .IN2(n351), .QN(n367) );
  NAND2X0 U105 ( .IN1(n612), .IN2(n611), .QN(N389) );
  NAND2X0 U106 ( .IN1(n616), .IN2(n615), .QN(N390) );
  NAND2X0 U107 ( .IN1(n620), .IN2(n619), .QN(N391) );
  NAND2X0 U108 ( .IN1(n624), .IN2(n623), .QN(N392) );
  NAND2X0 U109 ( .IN1(n628), .IN2(n627), .QN(N393) );
  NAND2X0 U110 ( .IN1(n632), .IN2(n631), .QN(N394) );
  NAND2X0 U111 ( .IN1(n636), .IN2(n635), .QN(N395) );
  NAND2X0 U112 ( .IN1(n640), .IN2(n639), .QN(N396) );
  NAND2X0 U113 ( .IN1(n721), .IN2(pre_sig_res_03[9]), .QN(n643) );
  NAND2X0 U114 ( .IN1(n720), .IN2(pre_sig_res_02[9]), .QN(n644) );
  NAND2X0 U115 ( .IN1(n721), .IN2(pre_sig_res_03[10]), .QN(n649) );
  NAND2X0 U116 ( .IN1(n720), .IN2(pre_sig_res_02[10]), .QN(n650) );
  NAND2X0 U117 ( .IN1(n721), .IN2(pre_sig_res_03[11]), .QN(n655) );
  NAND2X0 U118 ( .IN1(n720), .IN2(pre_sig_res_02[11]), .QN(n656) );
  NAND2X0 U119 ( .IN1(n721), .IN2(pre_sig_res_03[12]), .QN(n661) );
  NAND2X0 U120 ( .IN1(n720), .IN2(pre_sig_res_02[12]), .QN(n662) );
  NAND2X0 U121 ( .IN1(n721), .IN2(pre_sig_res_03[13]), .QN(n667) );
  NAND2X0 U122 ( .IN1(n720), .IN2(pre_sig_res_02[13]), .QN(n668) );
  NAND2X0 U123 ( .IN1(n7), .IN2(n8), .QN(N402) );
  NAND2X0 U124 ( .IN1(pre_sig_res_01[14]), .IN2(n723), .QN(n8) );
  NAND2X0 U125 ( .IN1(n721), .IN2(pre_sig_res_03[15]), .QN(n676) );
  NAND2X0 U126 ( .IN1(n720), .IN2(pre_sig_res_02[15]), .QN(n677) );
  NAND2X0 U127 ( .IN1(n722), .IN2(pre_sig_res_04[16]), .QN(n683) );
  NAND2X0 U128 ( .IN1(n722), .IN2(pre_sig_res_04[17]), .QN(n689) );
  NAND2X0 U129 ( .IN1(n722), .IN2(pre_sig_res_04[18]), .QN(n695) );
  NAND2X0 U130 ( .IN1(n722), .IN2(pre_sig_res_04[19]), .QN(n701) );
  NAND2X0 U131 ( .IN1(n722), .IN2(pre_sig_res_04[20]), .QN(n707) );
  NAND2X0 U132 ( .IN1(n722), .IN2(pre_sig_res_04[21]), .QN(n713) );
  NAND2X0 U133 ( .IN1(n722), .IN2(pre_sig_res_04[22]), .QN(n725) );
  NAND2X0 U134 ( .IN1(n722), .IN2(add_output_exponent_w4[0]), .QN(n572) );
  NAND2X0 U135 ( .IN1(n722), .IN2(add_output_exponent_w4[1]), .QN(n576) );
  NAND2X0 U136 ( .IN1(n722), .IN2(add_output_exponent_w4[2]), .QN(n580) );
  NAND2X0 U137 ( .IN1(n722), .IN2(add_output_exponent_w4[3]), .QN(n586) );
  NAND2X0 U138 ( .IN1(n722), .IN2(add_output_exponent_w4[4]), .QN(n592) );
  NAND2X0 U139 ( .IN1(n722), .IN2(add_output_exponent_w4[5]), .QN(n598) );
  NAND2X0 U140 ( .IN1(n722), .IN2(add_output_exponent_w4[6]), .QN(n604) );
  NAND2X0 U141 ( .IN1(n9), .IN2(n10), .QN(N387) );
  NAND2X0 U142 ( .IN1(n722), .IN2(add_output_exponent_w4[7]), .QN(n10) );
  NAND2X0 U143 ( .IN1(n521), .IN2(n520), .QN(N348) );
  NAND2X0 U144 ( .IN1(n538), .IN2(n808), .QN(n539) );
  NAND2X0 U145 ( .IN1(n538), .IN2(n828), .QN(n529) );
  NAND2X0 U146 ( .IN1(n538), .IN2(n830), .QN(n525) );
  NAND2X0 U147 ( .IN1(n523), .IN2(n522), .QN(N352) );
  NAND2X0 U148 ( .IN1(pre_sig_res_03[22]), .IN2(n832), .QN(n737) );
  NAND2X0 U149 ( .IN1(n821), .IN2(n736), .QN(n738) );
  NAND2X0 U150 ( .IN1(pre_sig_res_03[21]), .IN2(n832), .QN(n745) );
  NAND2X0 U151 ( .IN1(n821), .IN2(n744), .QN(n746) );
  NAND2X0 U152 ( .IN1(pre_sig_res_03[20]), .IN2(n832), .QN(n753) );
  NAND2X0 U153 ( .IN1(n821), .IN2(n752), .QN(n754) );
  NAND2X0 U154 ( .IN1(pre_sig_res_03[19]), .IN2(n832), .QN(n761) );
  NAND2X0 U155 ( .IN1(n821), .IN2(n760), .QN(n762) );
  NAND2X0 U156 ( .IN1(pre_sig_res_03[18]), .IN2(n832), .QN(n769) );
  NAND2X0 U157 ( .IN1(n821), .IN2(n768), .QN(n770) );
  NAND2X0 U158 ( .IN1(pre_sig_res_03[17]), .IN2(n832), .QN(n777) );
  NAND2X0 U159 ( .IN1(n821), .IN2(n776), .QN(n778) );
  NAND2X0 U160 ( .IN1(pre_sig_res_03[16]), .IN2(n832), .QN(n784) );
  NAND2X0 U161 ( .IN1(n821), .IN2(n801), .QN(n785) );
  NAND2X0 U162 ( .IN1(pre_sig_res_03[15]), .IN2(n832), .QN(n793) );
  NAND2X0 U163 ( .IN1(n821), .IN2(n809), .QN(n794) );
  NAND2X0 U164 ( .IN1(n728), .IN2(n735), .QN(n507) );
  NAND2X0 U165 ( .IN1(pre_sig_res_03[14]), .IN2(n861), .QN(n803) );
  NAND2X0 U166 ( .IN1(n831), .IN2(n801), .QN(n802) );
  NAND2X0 U167 ( .IN1(n821), .IN2(n800), .QN(n804) );
  NAND2X0 U168 ( .IN1(pre_sig_res_03[13]), .IN2(n832), .QN(n811) );
  NAND2X0 U169 ( .IN1(n831), .IN2(n809), .QN(n810) );
  NAND2X0 U170 ( .IN1(n821), .IN2(n808), .QN(n812) );
  NAND2X0 U171 ( .IN1(n816), .IN2(n815), .QN(n850) );
  NAND2X0 U172 ( .IN1(pre_sig_res_03[12]), .IN2(n832), .QN(n824) );
  NAND2X0 U173 ( .IN1(n821), .IN2(n828), .QN(n826) );
  NAND2X0 U174 ( .IN1(n414), .IN2(n828), .QN(n415) );
  NAND2X0 U175 ( .IN1(n419), .IN2(n809), .QN(n410) );
  NAND2X0 U176 ( .IN1(n420), .IN2(n808), .QN(n407) );
  NAND2X0 U177 ( .IN1(n406), .IN2(n405), .QN(N263) );
  NAND2X0 U178 ( .IN1(n351), .IN2(n116), .QN(n117) );
  NAND2X0 U179 ( .IN1(n353), .IN2(n86), .QN(n118) );
  NAND2X0 U180 ( .IN1(n351), .IN2(n146), .QN(n147) );
  NAND2X0 U181 ( .IN1(n353), .IN2(n137), .QN(n148) );
  NAND2X0 U182 ( .IN1(n351), .IN2(n173), .QN(n174) );
  NAND2X0 U183 ( .IN1(n353), .IN2(n165), .QN(n175) );
  NAND2X0 U184 ( .IN1(n351), .IN2(n204), .QN(n205) );
  NAND2X0 U185 ( .IN1(n353), .IN2(n194), .QN(n206) );
  NAND2X0 U186 ( .IN1(n280), .IN2(n298), .QN(n283) );
  NAND2X0 U187 ( .IN1(n281), .IN2(n300), .QN(n282) );
  NAND2X0 U188 ( .IN1(n286), .IN2(n298), .QN(n289) );
  NAND2X0 U189 ( .IN1(n287), .IN2(n300), .QN(n288) );
  NAND2X0 U190 ( .IN1(n292), .IN2(n298), .QN(n295) );
  NAND2X0 U191 ( .IN1(n293), .IN2(n300), .QN(n294) );
  NAND2X0 U192 ( .IN1(n299), .IN2(n298), .QN(n303) );
  NAND2X0 U193 ( .IN1(n301), .IN2(n300), .QN(n302) );
  NAND2X0 U194 ( .IN1(input_factor_01[14]), .IN2(n320), .QN(n321) );
  NAND2X0 U195 ( .IN1(n336), .IN2(n335), .QN(N168) );
  NAND2X0 U196 ( .IN1(n340), .IN2(n339), .QN(N169) );
  NAND2X0 U197 ( .IN1(n344), .IN2(n343), .QN(N170) );
  NAND2X0 U198 ( .IN1(n350), .IN2(n349), .QN(N171) );
  NAND2X0 U199 ( .IN1(n357), .IN2(n356), .QN(N172) );
  NAND2X0 U200 ( .IN1(n363), .IN2(n362), .QN(N173) );
  NAND2X0 U201 ( .IN1(n370), .IN2(n369), .QN(N174) );
  NAND2X0 U202 ( .IN1(n375), .IN2(n374), .QN(N175) );
  INVX0 U203 ( .INP(n393), .ZN(n392) );
  NOR2X0 U204 ( .IN1(n834), .IN2(n861), .QN(n835) );
  NOR2X0 U205 ( .IN1(n833), .IN2(n832), .QN(n836) );
  INVX0 U206 ( .INP(n563), .ZN(n838) );
  INVX0 U207 ( .INP(n419), .ZN(n491) );
  NOR2X0 U208 ( .IN1(n735), .IN2(n832), .QN(n821) );
  INVX0 U209 ( .INP(n829), .ZN(n819) );
  INVX0 U210 ( .INP(n808), .ZN(n820) );
  INVX0 U211 ( .INP(n809), .ZN(n798) );
  INVX0 U212 ( .INP(n776), .ZN(n789) );
  NOR2X0 U213 ( .IN1(n566), .IN2(n569), .QN(n720) );
  NOR2X0 U214 ( .IN1(n567), .IN2(n569), .QN(n721) );
  INVX0 U215 ( .INP(n752), .ZN(n765) );
  INVX0 U216 ( .INP(n456), .ZN(n565) );
  INVX0 U217 ( .INP(n564), .ZN(n514) );
  INVX0 U218 ( .INP(n760), .ZN(n773) );
  NOR2X0 U219 ( .IN1(n570), .IN2(n569), .QN(n723) );
  INVX0 U220 ( .INP(n4), .ZN(n18) );
  INVX0 U221 ( .INP(n220), .ZN(n716) );
  INVX0 U222 ( .INP(n320), .ZN(n360) );
  NOR2X0 U223 ( .IN1(n833), .IN2(n373), .QN(n353) );
  INVX0 U224 ( .INP(n834), .ZN(n833) );
  NOR2X0 U225 ( .IN1(n364), .IN2(n72), .QN(n834) );
  INVX0 U226 ( .INP(n328), .ZN(n372) );
  NOR2X0 U227 ( .IN1(exp_diff_value[1]), .IN2(exp_diff_value[0]), .QN(n328) );
  INVX0 U228 ( .INP(n398), .ZN(n494) );
  NOR2X0 U229 ( .IN1(add_sub_result_24_), .IN2(n395), .QN(n570) );
  MUX21X1 U230 ( .IN1(add_result[24]), .IN2(sub_result[24]), .S(n16), .Q(
        add_sub_result_24_) );
  INVX0 U231 ( .INP(n396), .ZN(n484) );
  INVX0 U232 ( .INP(n17), .ZN(n16) );
  INVX0 U233 ( .INP(n503), .ZN(n17) );
  INVX0 U234 ( .INP(n744), .ZN(n757) );
  INVX0 U235 ( .INP(n768), .ZN(n781) );
  INVX0 U236 ( .INP(n801), .ZN(n788) );
  INVX0 U237 ( .INP(n800), .ZN(n818) );
  INVX0 U238 ( .INP(n828), .ZN(n814) );
  INVX0 U239 ( .INP(n830), .ZN(n822) );
  MUX21X1 U240 ( .IN1(input_factor_01[31]), .IN2(n551), .S(input_factor_02[31]), .Q(n503) );
  INVX0 U241 ( .INP(input_factor_01[31]), .ZN(n551) );
  INVX0 U242 ( .INP(input_factor_02[22]), .ZN(n719) );
  INVX0 U243 ( .INP(n375), .ZN(n364) );
  NAND2X0 U244 ( .IN1(input_factor_02[29]), .IN2(n601), .QN(n44) );
  INVX0 U245 ( .INP(input_factor_02[23]), .ZN(n559) );
  INVX0 U246 ( .INP(input_factor_02[29]), .ZN(n602) );
  NAND4X0 U247 ( .IN1(n27), .IN2(n26), .IN3(n550), .IN4(n30), .QN(n375) );
  NAND3X0 U248 ( .IN1(n562), .IN2(n18), .IN3(n718), .QN(n569) );
  INVX0 U249 ( .INP(n447), .ZN(n730) );
  INVX0 U250 ( .INP(n442), .ZN(n741) );
  INVX0 U251 ( .INP(n736), .ZN(n749) );
  INVX0 U252 ( .INP(n831), .ZN(n817) );
  NOR2X0 U253 ( .IN1(n673), .IN2(n672), .QN(n7) );
  NOR2X0 U254 ( .IN1(n608), .IN2(n607), .QN(n9) );
  NAND3X0 U255 ( .IN1(n494), .IN2(n401), .IN3(n465), .QN(n483) );
  OR2X1 U256 ( .IN1(n561), .IN2(n765), .Q(n797) );
  NOR2X0 U257 ( .IN1(n11), .IN2(n12), .QN(n213) );
  NOR2X0 U258 ( .IN1(n699), .IN2(n199), .QN(n11) );
  NOR2X0 U259 ( .IN1(exp_diff_value[3]), .IN2(exp_diff_value[2]), .QN(n352) );
  NOR2X0 U260 ( .IN1(n220), .IN2(n373), .QN(n351) );
  NOR2X0 U261 ( .IN1(exp_diff_value[3]), .IN2(n1), .QN(n209) );
  MUX21X1 U262 ( .IN1(add_result[1]), .IN2(sub_result[1]), .S(n503), .Q(n828)
         );
  INVX0 U263 ( .INP(n200), .ZN(n15) );
  AND3X1 U264 ( .IN1(n391), .IN2(n390), .IN3(n389), .Q(n4) );
  INVX0 U265 ( .INP(n718), .ZN(n19) );
  AND2X1 U266 ( .IN1(exp_diff_value[1]), .IN2(n3), .Q(n5) );
  INVX0 U267 ( .INP(n199), .ZN(n14) );
  INVX0 U268 ( .INP(n5), .ZN(n13) );
  INVX0 U269 ( .INP(input_factor_01[29]), .ZN(n601) );
  OA222X1 U270 ( .IN1(input_factor_02[29]), .IN2(n601), .IN3(n602), .IN4(
        input_factor_01[29]), .IN5(input_factor_01[23]), .IN6(n559), .Q(n27)
         );
  INVX0 U271 ( .INP(input_factor_01[25]), .ZN(n549) );
  INVX0 U272 ( .INP(n31), .ZN(n25) );
  NOR2X0 U273 ( .IN1(input_factor_02[25]), .IN2(n549), .QN(n36) );
  INVX0 U274 ( .INP(input_factor_02[28]), .ZN(n596) );
  INVX0 U275 ( .INP(input_factor_02[26]), .ZN(n584) );
  INVX0 U276 ( .INP(input_factor_01[28]), .ZN(n595) );
  INVX0 U277 ( .INP(input_factor_01[26]), .ZN(n583) );
  NAND4X0 U278 ( .IN1(n39), .IN2(n29), .IN3(n43), .IN4(n20), .QN(n24) );
  INVX0 U279 ( .INP(input_factor_01[27]), .ZN(n589) );
  INVX0 U280 ( .INP(input_factor_02[27]), .ZN(n590) );
  INVX0 U281 ( .INP(input_factor_01[24]), .ZN(n548) );
  NOR2X0 U282 ( .IN1(n548), .IN2(input_factor_02[24]), .QN(n34) );
  INVX0 U283 ( .INP(n34), .ZN(n21) );
  NAND4X0 U284 ( .IN1(n22), .IN2(n28), .IN3(n32), .IN4(n21), .QN(n23) );
  NOR4X0 U285 ( .IN1(n25), .IN2(n36), .IN3(n24), .IN4(n23), .QN(n26) );
  INVX0 U286 ( .INP(input_factor_01[30]), .ZN(n550) );
  INVX0 U287 ( .INP(n28), .ZN(n42) );
  INVX0 U288 ( .INP(n29), .ZN(n38) );
  INVX0 U289 ( .INP(n30), .ZN(n33) );
  OA221X1 U290 ( .IN1(n34), .IN2(n33), .IN3(n34), .IN4(n32), .IN5(n31), .Q(n35) );
  OA22X1 U291 ( .IN1(n36), .IN2(n35), .IN3(input_factor_01[26]), .IN4(n584), 
        .Q(n37) );
  OA22X1 U292 ( .IN1(n38), .IN2(n37), .IN3(input_factor_01[27]), .IN4(n590), 
        .Q(n41) );
  INVX0 U293 ( .INP(n39), .ZN(n40) );
  AO221X1 U294 ( .IN1(n43), .IN2(n42), .IN3(n43), .IN4(n41), .IN5(n40), .Q(n45) );
  AO221X1 U295 ( .IN1(n45), .IN2(n44), .IN3(n602), .IN4(input_factor_01[29]), 
        .IN5(input_factor_01[30]), .Q(n72) );
  INVX0 U296 ( .INP(input_factor_02[21]), .ZN(n711) );
  INVX0 U297 ( .INP(input_factor_02[20]), .ZN(n705) );
  INVX0 U298 ( .INP(input_factor_02[19]), .ZN(n699) );
  INVX0 U299 ( .INP(input_factor_02[18]), .ZN(n693) );
  INVX0 U300 ( .INP(input_factor_02[17]), .ZN(n687) );
  INVX0 U301 ( .INP(input_factor_02[16]), .ZN(n681) );
  INVX0 U302 ( .INP(input_factor_02[15]), .ZN(n675) );
  INVX0 U303 ( .INP(input_factor_02[12]), .ZN(n660) );
  INVX0 U304 ( .INP(input_factor_02[11]), .ZN(n654) );
  INVX0 U305 ( .INP(input_factor_02[10]), .ZN(n648) );
  INVX0 U306 ( .INP(input_factor_02[9]), .ZN(n642) );
  INVX0 U307 ( .INP(input_factor_02[8]), .ZN(n638) );
  INVX0 U308 ( .INP(input_factor_02[7]), .ZN(n634) );
  INVX0 U309 ( .INP(input_factor_02[6]), .ZN(n630) );
  INVX0 U310 ( .INP(input_factor_02[5]), .ZN(n626) );
  INVX0 U311 ( .INP(input_factor_02[4]), .ZN(n622) );
  INVX0 U312 ( .INP(input_factor_02[3]), .ZN(n618) );
  INVX0 U313 ( .INP(input_factor_02[2]), .ZN(n614) );
  INVX0 U314 ( .INP(input_factor_01[0]), .ZN(n543) );
  NOR2X0 U315 ( .IN1(input_factor_02[0]), .IN2(n543), .QN(n46) );
  INVX0 U316 ( .INP(input_factor_02[1]), .ZN(n610) );
  AO222X1 U317 ( .IN1(input_factor_01[1]), .IN2(n46), .IN3(input_factor_01[1]), 
        .IN4(n610), .IN5(n46), .IN6(n610), .Q(n47) );
  AO222X1 U318 ( .IN1(input_factor_01[2]), .IN2(n614), .IN3(input_factor_01[2]), .IN4(n47), .IN5(n614), .IN6(n47), .Q(n48) );
  AO222X1 U319 ( .IN1(input_factor_01[3]), .IN2(n618), .IN3(input_factor_01[3]), .IN4(n48), .IN5(n618), .IN6(n48), .Q(n49) );
  AO222X1 U320 ( .IN1(input_factor_01[4]), .IN2(n622), .IN3(input_factor_01[4]), .IN4(n49), .IN5(n622), .IN6(n49), .Q(n50) );
  AO222X1 U321 ( .IN1(input_factor_01[5]), .IN2(n626), .IN3(input_factor_01[5]), .IN4(n50), .IN5(n626), .IN6(n50), .Q(n51) );
  AO222X1 U322 ( .IN1(input_factor_01[6]), .IN2(n630), .IN3(input_factor_01[6]), .IN4(n51), .IN5(n630), .IN6(n51), .Q(n52) );
  AO222X1 U323 ( .IN1(input_factor_01[7]), .IN2(n634), .IN3(input_factor_01[7]), .IN4(n52), .IN5(n634), .IN6(n52), .Q(n53) );
  AO222X1 U324 ( .IN1(input_factor_01[8]), .IN2(n638), .IN3(input_factor_01[8]), .IN4(n53), .IN5(n638), .IN6(n53), .Q(n54) );
  AO222X1 U325 ( .IN1(input_factor_01[9]), .IN2(n642), .IN3(input_factor_01[9]), .IN4(n54), .IN5(n642), .IN6(n54), .Q(n55) );
  AO222X1 U326 ( .IN1(input_factor_01[10]), .IN2(n648), .IN3(
        input_factor_01[10]), .IN4(n55), .IN5(n648), .IN6(n55), .Q(n56) );
  AO222X1 U327 ( .IN1(input_factor_01[11]), .IN2(n654), .IN3(
        input_factor_01[11]), .IN4(n56), .IN5(n654), .IN6(n56), .Q(n57) );
  AO222X1 U328 ( .IN1(input_factor_01[12]), .IN2(n660), .IN3(
        input_factor_01[12]), .IN4(n57), .IN5(n660), .IN6(n57), .Q(n59) );
  INVX0 U329 ( .INP(input_factor_01[13]), .ZN(n665) );
  INVX0 U330 ( .INP(input_factor_02[13]), .ZN(n666) );
  AO221X1 U331 ( .IN1(n59), .IN2(n58), .IN3(n666), .IN4(input_factor_01[13]), 
        .IN5(input_factor_01[14]), .Q(n60) );
  AO222X1 U332 ( .IN1(input_factor_01[15]), .IN2(n675), .IN3(
        input_factor_01[15]), .IN4(n60), .IN5(n675), .IN6(n60), .Q(n61) );
  AO222X1 U333 ( .IN1(input_factor_01[16]), .IN2(n681), .IN3(
        input_factor_01[16]), .IN4(n61), .IN5(n681), .IN6(n61), .Q(n62) );
  AO222X1 U334 ( .IN1(input_factor_01[17]), .IN2(n687), .IN3(
        input_factor_01[17]), .IN4(n62), .IN5(n687), .IN6(n62), .Q(n63) );
  AO222X1 U335 ( .IN1(input_factor_01[18]), .IN2(n693), .IN3(
        input_factor_01[18]), .IN4(n63), .IN5(n693), .IN6(n63), .Q(n64) );
  AO222X1 U336 ( .IN1(input_factor_01[19]), .IN2(n699), .IN3(
        input_factor_01[19]), .IN4(n64), .IN5(n699), .IN6(n64), .Q(n65) );
  AO222X1 U337 ( .IN1(input_factor_01[20]), .IN2(n705), .IN3(
        input_factor_01[20]), .IN4(n65), .IN5(n705), .IN6(n65), .Q(n66) );
  AO222X1 U338 ( .IN1(input_factor_01[21]), .IN2(n711), .IN3(
        input_factor_01[21]), .IN4(n66), .IN5(n711), .IN6(n66), .Q(n67) );
  AO222X1 U339 ( .IN1(input_factor_01[22]), .IN2(n719), .IN3(
        input_factor_01[22]), .IN4(n67), .IN5(n719), .IN6(n67), .Q(n74) );
  INVX0 U340 ( .INP(input_factor_01[14]), .ZN(n671) );
  NOR2X0 U341 ( .IN1(n392), .IN2(n671), .QN(N190) );
  AO22X1 U342 ( .IN1(input_factor_01[30]), .IN2(rst_n), .IN3(n861), .IN4(
        larger_exponent[7]), .Q(n839) );
  OA22X1 U344 ( .IN1(n687), .IN2(n200), .IN3(n693), .IN4(n13), .Q(n69) );
  AO222X1 U345 ( .IN1(n711), .IN2(n15), .IN3(n705), .IN4(n328), .IN5(n719), 
        .IN6(n5), .Q(n355) );
  MUX21X1 U346 ( .IN1(n213), .IN2(n355), .S(exp_diff_value[2]), .Q(n333) );
  AO22X1 U347 ( .IN1(input_factor_01[18]), .IN2(n5), .IN3(input_factor_01[16]), 
        .IN4(n328), .Q(n71) );
  AO22X1 U348 ( .IN1(input_factor_01[19]), .IN2(n14), .IN3(input_factor_01[17]), .IN4(n15), .Q(n70) );
  NOR2X0 U349 ( .IN1(n71), .IN2(n70), .QN(n216) );
  INVX0 U350 ( .INP(input_factor_01[22]), .ZN(n717) );
  INVX0 U351 ( .INP(input_factor_01[21]), .ZN(n710) );
  INVX0 U352 ( .INP(input_factor_01[20]), .ZN(n704) );
  AO222X1 U353 ( .IN1(n5), .IN2(n717), .IN3(n15), .IN4(n710), .IN5(n328), 
        .IN6(n704), .Q(n354) );
  MUX21X1 U354 ( .IN1(n216), .IN2(n354), .S(exp_diff_value[2]), .Q(n334) );
  OA22X1 U355 ( .IN1(n333), .IN2(n220), .IN3(n334), .IN4(n833), .Q(n75) );
  NOR3X0 U356 ( .IN1(exp_diff_value[5]), .IN2(exp_diff_value[6]), .IN3(
        exp_diff_value[7]), .QN(n73) );
  AND2X1 U357 ( .IN1(exp_diff_value[4]), .IN2(n73), .Q(n273) );
  NOR2X0 U358 ( .IN1(n375), .IN2(n74), .QN(n320) );
  OA22X1 U359 ( .IN1(n75), .IN2(n182), .IN3(n543), .IN4(n360), .Q(n120) );
  INVX0 U360 ( .INP(n361), .ZN(n184) );
  OR4X1 U361 ( .IN1(exp_diff_value[4]), .IN2(exp_diff_value[5]), .IN3(
        exp_diff_value[6]), .IN4(exp_diff_value[7]), .Q(n373) );
  INVX0 U362 ( .INP(input_factor_01[2]), .ZN(n613) );
  OA22X1 U363 ( .IN1(n613), .IN2(n13), .IN3(n543), .IN4(n372), .Q(n77) );
  INVX0 U364 ( .INP(input_factor_01[3]), .ZN(n617) );
  INVX0 U365 ( .INP(input_factor_01[1]), .ZN(n609) );
  OA22X1 U366 ( .IN1(n617), .IN2(n199), .IN3(n609), .IN4(n200), .Q(n76) );
  INVX0 U367 ( .INP(input_factor_01[6]), .ZN(n629) );
  INVX0 U368 ( .INP(input_factor_01[4]), .ZN(n621) );
  OA22X1 U369 ( .IN1(n629), .IN2(n13), .IN3(n621), .IN4(n372), .Q(n80) );
  INVX0 U370 ( .INP(input_factor_01[7]), .ZN(n633) );
  INVX0 U371 ( .INP(input_factor_01[5]), .ZN(n625) );
  OA22X1 U372 ( .IN1(n633), .IN2(n199), .IN3(n625), .IN4(n200), .Q(n79) );
  INVX0 U373 ( .INP(input_factor_01[10]), .ZN(n647) );
  INVX0 U374 ( .INP(input_factor_01[8]), .ZN(n637) );
  OA22X1 U375 ( .IN1(n647), .IN2(n13), .IN3(n637), .IN4(n372), .Q(n82) );
  INVX0 U376 ( .INP(input_factor_01[11]), .ZN(n653) );
  INVX0 U377 ( .INP(input_factor_01[9]), .ZN(n641) );
  OA22X1 U378 ( .IN1(n653), .IN2(n199), .IN3(n641), .IN4(n200), .Q(n81) );
  INVX0 U379 ( .INP(input_factor_01[12]), .ZN(n659) );
  OA22X1 U380 ( .IN1(n671), .IN2(n13), .IN3(n659), .IN4(n372), .Q(n84) );
  INVX0 U381 ( .INP(input_factor_01[15]), .ZN(n674) );
  OA22X1 U382 ( .IN1(n674), .IN2(n199), .IN3(n665), .IN4(n200), .Q(n83) );
  MUX21X1 U383 ( .IN1(n210), .IN2(n215), .S(exp_diff_value[2]), .Q(n281) );
  AO222X1 U384 ( .IN1(n85), .IN2(n352), .IN3(n219), .IN4(n209), .IN5(n281), 
        .IN6(exp_diff_value[3]), .Q(n86) );
  AOI22X1 U385 ( .IN1(input_factor_02[0]), .IN2(n328), .IN3(input_factor_02[2]), .IN4(n5), .QN(n88) );
  OA22X1 U386 ( .IN1(n610), .IN2(n200), .IN3(n618), .IN4(n199), .Q(n87) );
  OA22X1 U387 ( .IN1(n622), .IN2(n372), .IN3(n630), .IN4(n13), .Q(n90) );
  OA22X1 U388 ( .IN1(n626), .IN2(n200), .IN3(n634), .IN4(n199), .Q(n89) );
  OA22X1 U389 ( .IN1(n638), .IN2(n372), .IN3(n648), .IN4(n13), .Q(n92) );
  OA22X1 U390 ( .IN1(n654), .IN2(n199), .IN3(n642), .IN4(n200), .Q(n91) );
  AO222X1 U391 ( .IN1(input_factor_02[12]), .IN2(n328), .IN3(
        input_factor_02[13]), .IN4(n15), .IN5(input_factor_02[15]), .IN6(n14), 
        .Q(n212) );
  MUX21X1 U392 ( .IN1(n211), .IN2(n212), .S(exp_diff_value[2]), .Q(n280) );
  AO222X1 U393 ( .IN1(n93), .IN2(n352), .IN3(n218), .IN4(n209), .IN5(n280), 
        .IN6(exp_diff_value[3]), .Q(n116) );
  NAND4X0 U394 ( .IN1(n120), .IN2(n119), .IN3(n118), .IN4(n117), .QN(N152) );
  AO22X1 U395 ( .IN1(input_factor_02[17]), .IN2(n328), .IN3(
        input_factor_02[19]), .IN4(n5), .Q(n122) );
  AO22X1 U396 ( .IN1(input_factor_02[18]), .IN2(n15), .IN3(input_factor_02[20]), .IN4(n14), .Q(n121) );
  NOR2X0 U397 ( .IN1(n122), .IN2(n121), .QN(n230) );
  AO22X1 U398 ( .IN1(input_factor_02[21]), .IN2(n3), .IN3(input_factor_02[22]), 
        .IN4(n15), .Q(n123) );
  NOR2X0 U399 ( .IN1(n5), .IN2(n123), .QN(n358) );
  MUX21X1 U400 ( .IN1(n230), .IN2(n358), .S(exp_diff_value[2]), .Q(n338) );
  AO22X1 U401 ( .IN1(input_factor_01[19]), .IN2(n5), .IN3(input_factor_01[17]), 
        .IN4(n328), .Q(n125) );
  AO22X1 U402 ( .IN1(input_factor_01[20]), .IN2(n14), .IN3(input_factor_01[18]), .IN4(n15), .Q(n124) );
  NOR2X0 U403 ( .IN1(n125), .IN2(n124), .QN(n233) );
  AO22X1 U404 ( .IN1(input_factor_01[22]), .IN2(n15), .IN3(input_factor_01[21]), .IN4(n3), .Q(n126) );
  NOR2X0 U405 ( .IN1(n5), .IN2(n126), .QN(n359) );
  MUX21X1 U406 ( .IN1(n233), .IN2(n359), .S(exp_diff_value[2]), .Q(n337) );
  OA22X1 U407 ( .IN1(n220), .IN2(n338), .IN3(n833), .IN4(n337), .Q(n127) );
  OA22X1 U408 ( .IN1(n127), .IN2(n182), .IN3(n609), .IN4(n360), .Q(n150) );
  OA22X1 U409 ( .IN1(n617), .IN2(n13), .IN3(n609), .IN4(n372), .Q(n129) );
  OA22X1 U410 ( .IN1(n621), .IN2(n199), .IN3(n613), .IN4(n200), .Q(n128) );
  OA22X1 U411 ( .IN1(n633), .IN2(n13), .IN3(n625), .IN4(n372), .Q(n131) );
  OA22X1 U412 ( .IN1(n637), .IN2(n199), .IN3(n629), .IN4(n200), .Q(n130) );
  OA22X1 U413 ( .IN1(n653), .IN2(n13), .IN3(n641), .IN4(n372), .Q(n133) );
  OA22X1 U414 ( .IN1(n659), .IN2(n199), .IN3(n647), .IN4(n200), .Q(n132) );
  OA22X1 U415 ( .IN1(n674), .IN2(n13), .IN3(n665), .IN4(n372), .Q(n135) );
  INVX0 U416 ( .INP(input_factor_01[16]), .ZN(n680) );
  OA22X1 U417 ( .IN1(n680), .IN2(n199), .IN3(n671), .IN4(n200), .Q(n134) );
  MUX21X1 U418 ( .IN1(n227), .IN2(n232), .S(exp_diff_value[2]), .Q(n287) );
  AO222X1 U419 ( .IN1(n136), .IN2(n352), .IN3(n236), .IN4(n209), .IN5(n287), 
        .IN6(exp_diff_value[3]), .Q(n137) );
  OA22X1 U420 ( .IN1(n610), .IN2(n372), .IN3(n618), .IN4(n13), .Q(n140) );
  OA22X1 U421 ( .IN1(n614), .IN2(n200), .IN3(n622), .IN4(n199), .Q(n139) );
  OA22X1 U422 ( .IN1(n626), .IN2(n372), .IN3(n634), .IN4(n13), .Q(n142) );
  OA22X1 U423 ( .IN1(n630), .IN2(n200), .IN3(n638), .IN4(n199), .Q(n141) );
  OA22X1 U424 ( .IN1(n654), .IN2(n13), .IN3(n642), .IN4(n372), .Q(n144) );
  OA22X1 U425 ( .IN1(n660), .IN2(n199), .IN3(n648), .IN4(n200), .Q(n143) );
  AO222X1 U426 ( .IN1(input_factor_02[15]), .IN2(n5), .IN3(input_factor_02[13]), .IN4(n328), .IN5(input_factor_02[16]), .IN6(n14), .Q(n229) );
  MUX21X1 U427 ( .IN1(n228), .IN2(n229), .S(exp_diff_value[2]), .Q(n286) );
  AO222X1 U428 ( .IN1(n145), .IN2(n352), .IN3(n235), .IN4(n209), .IN5(n286), 
        .IN6(exp_diff_value[3]), .Q(n146) );
  NAND4X0 U429 ( .IN1(n150), .IN2(n149), .IN3(n148), .IN4(n147), .QN(N153) );
  AO22X1 U430 ( .IN1(input_factor_02[18]), .IN2(n328), .IN3(
        input_factor_02[20]), .IN4(n5), .Q(n152) );
  AO22X1 U431 ( .IN1(input_factor_02[21]), .IN2(n14), .IN3(input_factor_02[19]), .IN4(n15), .Q(n151) );
  NOR2X0 U432 ( .IN1(n152), .IN2(n151), .QN(n246) );
  AO21X1 U433 ( .IN1(n719), .IN2(n3), .IN3(exp_diff_value[1]), .Q(n368) );
  MUX21X1 U434 ( .IN1(n246), .IN2(n368), .S(exp_diff_value[2]), .Q(n341) );
  AO22X1 U435 ( .IN1(input_factor_01[20]), .IN2(n5), .IN3(input_factor_01[18]), 
        .IN4(n328), .Q(n154) );
  AO22X1 U436 ( .IN1(input_factor_01[21]), .IN2(n14), .IN3(input_factor_01[19]), .IN4(n15), .Q(n153) );
  NOR2X0 U437 ( .IN1(n154), .IN2(n153), .QN(n249) );
  AO21X1 U438 ( .IN1(n717), .IN2(n3), .IN3(exp_diff_value[1]), .Q(n366) );
  MUX21X1 U439 ( .IN1(n249), .IN2(n366), .S(exp_diff_value[2]), .Q(n342) );
  OA22X1 U440 ( .IN1(n341), .IN2(n220), .IN3(n342), .IN4(n833), .Q(n155) );
  OA22X1 U441 ( .IN1(n155), .IN2(n182), .IN3(n613), .IN4(n360), .Q(n177) );
  OA22X1 U442 ( .IN1(n621), .IN2(n13), .IN3(n613), .IN4(n372), .Q(n157) );
  OA22X1 U443 ( .IN1(n625), .IN2(n199), .IN3(n617), .IN4(n200), .Q(n156) );
  OA22X1 U444 ( .IN1(n637), .IN2(n13), .IN3(n629), .IN4(n372), .Q(n159) );
  OA22X1 U445 ( .IN1(n641), .IN2(n199), .IN3(n633), .IN4(n200), .Q(n158) );
  OA22X1 U446 ( .IN1(n659), .IN2(n13), .IN3(n647), .IN4(n372), .Q(n161) );
  OA22X1 U447 ( .IN1(n665), .IN2(n199), .IN3(n653), .IN4(n200), .Q(n160) );
  OA22X1 U448 ( .IN1(n680), .IN2(n13), .IN3(n671), .IN4(n372), .Q(n163) );
  INVX0 U449 ( .INP(input_factor_01[17]), .ZN(n686) );
  OA22X1 U450 ( .IN1(n686), .IN2(n199), .IN3(n674), .IN4(n200), .Q(n162) );
  MUX21X1 U451 ( .IN1(n243), .IN2(n248), .S(exp_diff_value[2]), .Q(n293) );
  AO222X1 U452 ( .IN1(n164), .IN2(n352), .IN3(n252), .IN4(n209), .IN5(n293), 
        .IN6(exp_diff_value[3]), .Q(n165) );
  OA22X1 U453 ( .IN1(n614), .IN2(n372), .IN3(n622), .IN4(n13), .Q(n167) );
  OA22X1 U454 ( .IN1(n618), .IN2(n200), .IN3(n626), .IN4(n199), .Q(n166) );
  OA22X1 U455 ( .IN1(n630), .IN2(n372), .IN3(n638), .IN4(n13), .Q(n169) );
  OA22X1 U456 ( .IN1(n634), .IN2(n200), .IN3(n642), .IN4(n199), .Q(n168) );
  OA22X1 U457 ( .IN1(n660), .IN2(n13), .IN3(n648), .IN4(n372), .Q(n171) );
  OA22X1 U458 ( .IN1(n654), .IN2(n200), .IN3(n666), .IN4(n199), .Q(n170) );
  AO222X1 U459 ( .IN1(input_factor_02[15]), .IN2(n15), .IN3(
        input_factor_02[17]), .IN4(n14), .IN5(input_factor_02[16]), .IN6(n5), 
        .Q(n245) );
  MUX21X1 U460 ( .IN1(n244), .IN2(n245), .S(exp_diff_value[2]), .Q(n292) );
  AO222X1 U461 ( .IN1(n172), .IN2(n352), .IN3(n251), .IN4(n209), .IN5(n292), 
        .IN6(exp_diff_value[3]), .Q(n173) );
  NAND4X0 U462 ( .IN1(n177), .IN2(n176), .IN3(n175), .IN4(n174), .QN(N154) );
  AO22X1 U463 ( .IN1(input_factor_02[21]), .IN2(n5), .IN3(input_factor_02[19]), 
        .IN4(n328), .Q(n179) );
  AO22X1 U464 ( .IN1(input_factor_02[20]), .IN2(n15), .IN3(input_factor_02[22]), .IN4(n14), .Q(n178) );
  NOR2X0 U465 ( .IN1(n179), .IN2(n178), .QN(n266) );
  MUX21X1 U466 ( .IN1(n266), .IN2(n372), .S(exp_diff_value[2]), .Q(n346) );
  AO22X1 U467 ( .IN1(input_factor_01[21]), .IN2(n5), .IN3(input_factor_01[19]), 
        .IN4(n328), .Q(n181) );
  AO22X1 U468 ( .IN1(input_factor_01[22]), .IN2(n14), .IN3(input_factor_01[20]), .IN4(n15), .Q(n180) );
  NOR2X0 U469 ( .IN1(n181), .IN2(n180), .QN(n269) );
  MUX21X1 U470 ( .IN1(n269), .IN2(n372), .S(exp_diff_value[2]), .Q(n348) );
  OA22X1 U471 ( .IN1(n346), .IN2(n220), .IN3(n348), .IN4(n833), .Q(n183) );
  OA22X1 U472 ( .IN1(n183), .IN2(n182), .IN3(n617), .IN4(n360), .Q(n208) );
  OA22X1 U473 ( .IN1(n625), .IN2(n13), .IN3(n617), .IN4(n372), .Q(n186) );
  OA22X1 U474 ( .IN1(n629), .IN2(n199), .IN3(n621), .IN4(n200), .Q(n185) );
  OA22X1 U475 ( .IN1(n641), .IN2(n13), .IN3(n633), .IN4(n372), .Q(n188) );
  OA22X1 U476 ( .IN1(n647), .IN2(n199), .IN3(n637), .IN4(n200), .Q(n187) );
  OA22X1 U477 ( .IN1(n665), .IN2(n13), .IN3(n653), .IN4(n372), .Q(n190) );
  OA22X1 U478 ( .IN1(n671), .IN2(n199), .IN3(n659), .IN4(n200), .Q(n189) );
  OA22X1 U479 ( .IN1(n686), .IN2(n13), .IN3(n674), .IN4(n372), .Q(n192) );
  INVX0 U480 ( .INP(input_factor_01[18]), .ZN(n692) );
  OA22X1 U481 ( .IN1(n692), .IN2(n199), .IN3(n680), .IN4(n200), .Q(n191) );
  MUX21X1 U482 ( .IN1(n261), .IN2(n268), .S(exp_diff_value[2]), .Q(n301) );
  AO222X1 U483 ( .IN1(n193), .IN2(n352), .IN3(n272), .IN4(n209), .IN5(n301), 
        .IN6(exp_diff_value[3]), .Q(n194) );
  OA22X1 U484 ( .IN1(n618), .IN2(n372), .IN3(n626), .IN4(n13), .Q(n196) );
  OA22X1 U485 ( .IN1(n622), .IN2(n200), .IN3(n630), .IN4(n199), .Q(n195) );
  OA22X1 U486 ( .IN1(n634), .IN2(n372), .IN3(n642), .IN4(n13), .Q(n198) );
  OA22X1 U487 ( .IN1(n638), .IN2(n200), .IN3(n648), .IN4(n199), .Q(n197) );
  AO222X1 U488 ( .IN1(input_factor_02[11]), .IN2(n328), .IN3(
        input_factor_02[13]), .IN4(n5), .IN5(n15), .IN6(input_factor_02[12]), 
        .Q(n263) );
  OA22X1 U489 ( .IN1(n675), .IN2(n372), .IN3(n687), .IN4(n13), .Q(n202) );
  OA22X1 U490 ( .IN1(n681), .IN2(n200), .IN3(n693), .IN4(n199), .Q(n201) );
  MUX21X1 U491 ( .IN1(n263), .IN2(n265), .S(exp_diff_value[2]), .Q(n299) );
  AO222X1 U492 ( .IN1(n203), .IN2(n352), .IN3(n271), .IN4(n209), .IN5(n299), 
        .IN6(exp_diff_value[3]), .Q(n204) );
  NAND4X0 U493 ( .IN1(n208), .IN2(n207), .IN3(n206), .IN4(n205), .QN(N155) );
  AND2X1 U494 ( .IN1(n209), .IN2(n351), .Q(n264) );
  AND2X1 U495 ( .IN1(n353), .IN2(n209), .Q(n262) );
  AOI22X1 U496 ( .IN1(n264), .IN2(n211), .IN3(n262), .IN4(n210), .QN(n226) );
  INVX0 U497 ( .INP(n212), .ZN(n214) );
  MUX21X1 U498 ( .IN1(n214), .IN2(n213), .S(exp_diff_value[2]), .Q(n307) );
  INVX0 U499 ( .INP(n215), .ZN(n217) );
  MUX21X1 U500 ( .IN1(n217), .IN2(n216), .S(exp_diff_value[2]), .Q(n306) );
  OA22X1 U501 ( .IN1(n326), .IN2(n307), .IN3(n327), .IN4(n306), .Q(n225) );
  OA22X1 U502 ( .IN1(n622), .IN2(n361), .IN3(n621), .IN4(n360), .Q(n224) );
  AOI22X1 U503 ( .IN1(n353), .IN2(n219), .IN3(n351), .IN4(n218), .QN(n222) );
  OA22X1 U504 ( .IN1(n355), .IN2(n254), .IN3(n354), .IN4(n253), .Q(n221) );
  INVX0 U505 ( .INP(n352), .ZN(n371) );
  AO21X1 U506 ( .IN1(n222), .IN2(n221), .IN3(n371), .Q(n223) );
  NAND4X0 U507 ( .IN1(n226), .IN2(n225), .IN3(n224), .IN4(n223), .QN(N156) );
  AOI22X1 U508 ( .IN1(n264), .IN2(n228), .IN3(n262), .IN4(n227), .QN(n242) );
  INVX0 U509 ( .INP(n229), .ZN(n231) );
  MUX21X1 U510 ( .IN1(n231), .IN2(n230), .S(exp_diff_value[2]), .Q(n312) );
  INVX0 U511 ( .INP(n232), .ZN(n234) );
  MUX21X1 U512 ( .IN1(n234), .IN2(n233), .S(exp_diff_value[2]), .Q(n311) );
  OA22X1 U513 ( .IN1(n326), .IN2(n312), .IN3(n327), .IN4(n311), .Q(n241) );
  OA22X1 U514 ( .IN1(n626), .IN2(n361), .IN3(n625), .IN4(n360), .Q(n240) );
  AOI22X1 U515 ( .IN1(n353), .IN2(n236), .IN3(n351), .IN4(n235), .QN(n238) );
  OA22X1 U516 ( .IN1(n359), .IN2(n253), .IN3(n358), .IN4(n254), .Q(n237) );
  AO21X1 U517 ( .IN1(n238), .IN2(n237), .IN3(n371), .Q(n239) );
  NAND4X0 U518 ( .IN1(n242), .IN2(n241), .IN3(n240), .IN4(n239), .QN(N157) );
  AOI22X1 U519 ( .IN1(n264), .IN2(n244), .IN3(n262), .IN4(n243), .QN(n260) );
  INVX0 U520 ( .INP(n245), .ZN(n247) );
  MUX21X1 U521 ( .IN1(n247), .IN2(n246), .S(exp_diff_value[2]), .Q(n317) );
  INVX0 U522 ( .INP(n248), .ZN(n250) );
  MUX21X1 U523 ( .IN1(n250), .IN2(n249), .S(exp_diff_value[2]), .Q(n316) );
  OA22X1 U524 ( .IN1(n326), .IN2(n317), .IN3(n327), .IN4(n316), .Q(n259) );
  OA22X1 U525 ( .IN1(n630), .IN2(n361), .IN3(n629), .IN4(n360), .Q(n258) );
  AOI22X1 U526 ( .IN1(n353), .IN2(n252), .IN3(n351), .IN4(n251), .QN(n256) );
  OA22X1 U527 ( .IN1(n368), .IN2(n254), .IN3(n366), .IN4(n253), .Q(n255) );
  AO21X1 U528 ( .IN1(n256), .IN2(n255), .IN3(n371), .Q(n257) );
  NAND4X0 U529 ( .IN1(n260), .IN2(n259), .IN3(n258), .IN4(n257), .QN(N158) );
  AOI22X1 U530 ( .IN1(n264), .IN2(n263), .IN3(n262), .IN4(n261), .QN(n279) );
  INVX0 U531 ( .INP(n265), .ZN(n267) );
  MUX21X1 U532 ( .IN1(n267), .IN2(n266), .S(exp_diff_value[2]), .Q(n325) );
  INVX0 U533 ( .INP(n268), .ZN(n270) );
  MUX21X1 U534 ( .IN1(n270), .IN2(n269), .S(exp_diff_value[2]), .Q(n324) );
  OA22X1 U535 ( .IN1(n326), .IN2(n325), .IN3(n327), .IN4(n324), .Q(n278) );
  OA22X1 U536 ( .IN1(n634), .IN2(n361), .IN3(n633), .IN4(n360), .Q(n277) );
  AOI22X1 U537 ( .IN1(n353), .IN2(n272), .IN3(n351), .IN4(n271), .QN(n275) );
  NAND3X0 U538 ( .IN1(n273), .IN2(n328), .IN3(n375), .QN(n274) );
  AO21X1 U539 ( .IN1(n275), .IN2(n274), .IN3(n371), .Q(n276) );
  NAND4X0 U540 ( .IN1(n279), .IN2(n278), .IN3(n277), .IN4(n276), .QN(N159) );
  OA22X1 U541 ( .IN1(n334), .IN2(n327), .IN3(n333), .IN4(n326), .Q(n285) );
  OA22X1 U542 ( .IN1(n638), .IN2(n361), .IN3(n637), .IN4(n360), .Q(n284) );
  INVX0 U543 ( .INP(n345), .ZN(n298) );
  INVX0 U544 ( .INP(n347), .ZN(n300) );
  NAND4X0 U545 ( .IN1(n285), .IN2(n284), .IN3(n283), .IN4(n282), .QN(N160) );
  OA22X1 U546 ( .IN1(n338), .IN2(n326), .IN3(n337), .IN4(n327), .Q(n291) );
  OA22X1 U547 ( .IN1(n642), .IN2(n361), .IN3(n641), .IN4(n360), .Q(n290) );
  NAND4X0 U548 ( .IN1(n291), .IN2(n290), .IN3(n289), .IN4(n288), .QN(N161) );
  OA22X1 U549 ( .IN1(n342), .IN2(n327), .IN3(n341), .IN4(n326), .Q(n297) );
  OA22X1 U550 ( .IN1(n648), .IN2(n361), .IN3(n647), .IN4(n360), .Q(n296) );
  NAND4X0 U551 ( .IN1(n297), .IN2(n296), .IN3(n295), .IN4(n294), .QN(N162) );
  OA22X1 U552 ( .IN1(n348), .IN2(n327), .IN3(n346), .IN4(n326), .Q(n305) );
  OA22X1 U553 ( .IN1(n654), .IN2(n361), .IN3(n653), .IN4(n360), .Q(n304) );
  NAND4X0 U554 ( .IN1(n305), .IN2(n304), .IN3(n303), .IN4(n302), .QN(N163) );
  OA22X1 U555 ( .IN1(n307), .IN2(n345), .IN3(n306), .IN4(n347), .Q(n310) );
  OR2X1 U556 ( .IN1(n326), .IN2(exp_diff_value[2]), .Q(n319) );
  OR2X1 U557 ( .IN1(n327), .IN2(exp_diff_value[2]), .Q(n318) );
  OA22X1 U558 ( .IN1(n355), .IN2(n319), .IN3(n354), .IN4(n318), .Q(n309) );
  OA22X1 U559 ( .IN1(n660), .IN2(n361), .IN3(n659), .IN4(n360), .Q(n308) );
  NAND3X0 U560 ( .IN1(n310), .IN2(n309), .IN3(n308), .QN(N164) );
  OA22X1 U561 ( .IN1(n312), .IN2(n345), .IN3(n311), .IN4(n347), .Q(n315) );
  OA22X1 U562 ( .IN1(n359), .IN2(n318), .IN3(n358), .IN4(n319), .Q(n314) );
  OA22X1 U563 ( .IN1(n666), .IN2(n361), .IN3(n665), .IN4(n360), .Q(n313) );
  NAND3X0 U564 ( .IN1(n315), .IN2(n314), .IN3(n313), .QN(N165) );
  OA22X1 U565 ( .IN1(n317), .IN2(n345), .IN3(n316), .IN4(n347), .Q(n323) );
  OA22X1 U566 ( .IN1(n368), .IN2(n319), .IN3(n366), .IN4(n318), .Q(n322) );
  NAND3X0 U567 ( .IN1(n323), .IN2(n322), .IN3(n321), .QN(N166) );
  OA22X1 U568 ( .IN1(n325), .IN2(n345), .IN3(n324), .IN4(n347), .Q(n332) );
  OA22X1 U569 ( .IN1(n675), .IN2(n361), .IN3(n674), .IN4(n360), .Q(n331) );
  NAND3X0 U570 ( .IN1(n329), .IN2(n1), .IN3(n328), .QN(n330) );
  NAND3X0 U571 ( .IN1(n332), .IN2(n331), .IN3(n330), .QN(N167) );
  OA22X1 U572 ( .IN1(n334), .IN2(n347), .IN3(n333), .IN4(n345), .Q(n336) );
  OA22X1 U573 ( .IN1(n681), .IN2(n361), .IN3(n680), .IN4(n360), .Q(n335) );
  OA22X1 U574 ( .IN1(n338), .IN2(n345), .IN3(n337), .IN4(n347), .Q(n340) );
  OA22X1 U575 ( .IN1(n687), .IN2(n361), .IN3(n686), .IN4(n360), .Q(n339) );
  OA22X1 U576 ( .IN1(n342), .IN2(n347), .IN3(n341), .IN4(n345), .Q(n344) );
  OA22X1 U577 ( .IN1(n693), .IN2(n361), .IN3(n692), .IN4(n360), .Q(n343) );
  OA22X1 U578 ( .IN1(n348), .IN2(n347), .IN3(n346), .IN4(n345), .Q(n350) );
  INVX0 U579 ( .INP(input_factor_01[19]), .ZN(n698) );
  OA22X1 U580 ( .IN1(n699), .IN2(n361), .IN3(n698), .IN4(n360), .Q(n349) );
  OA22X1 U581 ( .IN1(n355), .IN2(n367), .IN3(n354), .IN4(n365), .Q(n357) );
  OA22X1 U582 ( .IN1(n705), .IN2(n361), .IN3(n704), .IN4(n360), .Q(n356) );
  OA22X1 U583 ( .IN1(n359), .IN2(n365), .IN3(n358), .IN4(n367), .Q(n363) );
  OA22X1 U584 ( .IN1(n711), .IN2(n361), .IN3(n710), .IN4(n360), .Q(n362) );
  NAND3X0 U585 ( .IN1(input_factor_01[22]), .IN2(input_factor_02[22]), .IN3(
        n364), .QN(n370) );
  OA22X1 U586 ( .IN1(n368), .IN2(n367), .IN3(n366), .IN4(n365), .Q(n369) );
  OR3X1 U587 ( .IN1(n373), .IN2(n372), .IN3(n371), .Q(n374) );
  MUX21X1 U588 ( .IN1(input_factor_01[0]), .IN2(input_factor_02[0]), .S(n392), 
        .Q(N176) );
  MUX21X1 U589 ( .IN1(input_factor_01[1]), .IN2(input_factor_02[1]), .S(n392), 
        .Q(N177) );
  MUX21X1 U590 ( .IN1(input_factor_01[2]), .IN2(input_factor_02[2]), .S(n392), 
        .Q(N178) );
  MUX21X1 U591 ( .IN1(input_factor_01[3]), .IN2(input_factor_02[3]), .S(n392), 
        .Q(N179) );
  MUX21X1 U592 ( .IN1(input_factor_01[4]), .IN2(input_factor_02[4]), .S(n392), 
        .Q(N180) );
  MUX21X1 U593 ( .IN1(input_factor_01[5]), .IN2(input_factor_02[5]), .S(n392), 
        .Q(N181) );
  MUX21X1 U594 ( .IN1(input_factor_01[6]), .IN2(input_factor_02[6]), .S(n392), 
        .Q(N182) );
  MUX21X1 U595 ( .IN1(input_factor_01[7]), .IN2(input_factor_02[7]), .S(n392), 
        .Q(N183) );
  MUX21X1 U596 ( .IN1(input_factor_01[8]), .IN2(input_factor_02[8]), .S(n392), 
        .Q(N184) );
  MUX21X1 U597 ( .IN1(input_factor_01[9]), .IN2(input_factor_02[9]), .S(n392), 
        .Q(N185) );
  MUX21X1 U598 ( .IN1(input_factor_01[10]), .IN2(input_factor_02[10]), .S(n392), .Q(N186) );
  MUX21X1 U599 ( .IN1(input_factor_01[11]), .IN2(input_factor_02[11]), .S(n392), .Q(N187) );
  MUX21X1 U600 ( .IN1(input_factor_01[12]), .IN2(input_factor_02[12]), .S(n392), .Q(N188) );
  MUX21X1 U601 ( .IN1(input_factor_01[13]), .IN2(input_factor_02[13]), .S(n392), .Q(N189) );
  MUX21X1 U602 ( .IN1(input_factor_01[15]), .IN2(input_factor_02[15]), .S(n392), .Q(N191) );
  MUX21X1 U603 ( .IN1(input_factor_01[16]), .IN2(input_factor_02[16]), .S(n392), .Q(N192) );
  MUX21X1 U604 ( .IN1(input_factor_01[17]), .IN2(input_factor_02[17]), .S(n392), .Q(N193) );
  MUX21X1 U605 ( .IN1(input_factor_01[18]), .IN2(input_factor_02[18]), .S(n392), .Q(N194) );
  MUX21X1 U606 ( .IN1(input_factor_01[19]), .IN2(input_factor_02[19]), .S(n392), .Q(N195) );
  MUX21X1 U607 ( .IN1(input_factor_01[20]), .IN2(input_factor_02[20]), .S(n392), .Q(N196) );
  MUX21X1 U608 ( .IN1(input_factor_01[21]), .IN2(input_factor_02[21]), .S(n392), .Q(N197) );
  MUX21X1 U609 ( .IN1(input_factor_01[22]), .IN2(input_factor_02[22]), .S(n392), .Q(N198) );
  MUX21X1 U610 ( .IN1(add_result[0]), .IN2(sub_result[0]), .S(n503), .Q(n830)
         );
  MUX21X1 U611 ( .IN1(add_result[2]), .IN2(sub_result[2]), .S(n503), .Q(n808)
         );
  MUX21X1 U612 ( .IN1(add_result[3]), .IN2(sub_result[3]), .S(n503), .Q(n800)
         );
  MUX21X1 U613 ( .IN1(add_result[4]), .IN2(sub_result[4]), .S(n503), .Q(n809)
         );
  MUX21X1 U614 ( .IN1(add_result[5]), .IN2(sub_result[5]), .S(n503), .Q(n801)
         );
  MUX21X1 U615 ( .IN1(add_result[6]), .IN2(sub_result[6]), .S(n503), .Q(n776)
         );
  MUX21X1 U616 ( .IN1(add_result[7]), .IN2(sub_result[7]), .S(n503), .Q(n768)
         );
  MUX21X1 U617 ( .IN1(add_result[9]), .IN2(sub_result[9]), .S(n503), .Q(n752)
         );
  MUX21X1 U618 ( .IN1(add_result[10]), .IN2(sub_result[10]), .S(n503), .Q(n744) );
  NOR4X0 U619 ( .IN1(n503), .IN2(add_result[14]), .IN3(add_result[15]), .IN4(
        add_result[13]), .QN(n512) );
  NOR4X0 U620 ( .IN1(sub_result[15]), .IN2(sub_result[14]), .IN3(
        sub_result[13]), .IN4(n17), .QN(n510) );
  NOR2X0 U621 ( .IN1(n512), .IN2(n510), .QN(n379) );
  MUX21X1 U622 ( .IN1(add_result[11]), .IN2(sub_result[11]), .S(n503), .Q(n736) );
  MUX21X1 U623 ( .IN1(add_result[16]), .IN2(sub_result[16]), .S(n16), .Q(n396)
         );
  MUX21X1 U624 ( .IN1(add_result[17]), .IN2(sub_result[17]), .S(n16), .Q(n465)
         );
  MUX21X1 U625 ( .IN1(add_result[20]), .IN2(sub_result[20]), .S(n16), .Q(n399)
         );
  INVX0 U626 ( .INP(n399), .ZN(n492) );
  MUX21X1 U627 ( .IN1(add_result[22]), .IN2(sub_result[22]), .S(n16), .Q(n400)
         );
  INVX0 U628 ( .INP(n400), .ZN(n376) );
  MUX21X1 U629 ( .IN1(add_result[23]), .IN2(sub_result[23]), .S(n16), .Q(n395)
         );
  MUX21X1 U630 ( .IN1(add_result[21]), .IN2(sub_result[21]), .S(n16), .Q(n402)
         );
  NOR2X0 U631 ( .IN1(n403), .IN2(n402), .QN(n404) );
  MUX21X1 U632 ( .IN1(add_result[19]), .IN2(sub_result[19]), .S(n16), .Q(n474)
         );
  NOR2X0 U633 ( .IN1(n377), .IN2(n474), .QN(n401) );
  MUX21X1 U634 ( .IN1(add_result[18]), .IN2(sub_result[18]), .S(n16), .Q(n398)
         );
  NOR2X0 U635 ( .IN1(n465), .IN2(n378), .QN(n397) );
  MUX21X1 U636 ( .IN1(add_result[12]), .IN2(sub_result[12]), .S(n16), .Q(n442)
         );
  NOR4X0 U637 ( .IN1(n379), .IN2(n736), .IN3(n564), .IN4(n442), .QN(n731) );
  MUX21X1 U638 ( .IN1(add_result[8]), .IN2(sub_result[8]), .S(n16), .Q(n760)
         );
  NOR3X0 U639 ( .IN1(n752), .IN2(n561), .IN3(n760), .QN(n517) );
  NOR2X0 U640 ( .IN1(n776), .IN2(n380), .QN(n516) );
  NOR2X0 U641 ( .IN1(n809), .IN2(n381), .QN(n524) );
  NOR2X0 U642 ( .IN1(n808), .IN2(n382), .QN(n518) );
  NAND3X0 U643 ( .IN1(n822), .IN2(n814), .IN3(n518), .QN(n562) );
  NOR4X0 U644 ( .IN1(input_factor_02[15]), .IN2(input_factor_02[16]), .IN3(
        input_factor_02[17]), .IN4(input_factor_02[18]), .QN(n391) );
  NOR4X0 U645 ( .IN1(input_factor_02[31]), .IN2(input_factor_02[27]), .IN3(
        input_factor_02[24]), .IN4(input_factor_02[25]), .QN(n390) );
  NAND4X0 U646 ( .IN1(n602), .IN2(n559), .IN3(n596), .IN4(n584), .QN(n388) );
  NOR4X0 U647 ( .IN1(input_factor_02[0]), .IN2(input_factor_02[1]), .IN3(
        input_factor_02[2]), .IN4(input_factor_02[3]), .QN(n386) );
  NOR4X0 U648 ( .IN1(input_factor_02[21]), .IN2(input_factor_02[19]), .IN3(
        input_factor_02[20]), .IN4(input_factor_02[22]), .QN(n385) );
  NOR4X0 U649 ( .IN1(input_factor_02[8]), .IN2(input_factor_02[9]), .IN3(
        input_factor_02[10]), .IN4(input_factor_02[13]), .QN(n384) );
  NOR4X0 U650 ( .IN1(input_factor_02[4]), .IN2(input_factor_02[5]), .IN3(
        input_factor_02[6]), .IN4(input_factor_02[7]), .QN(n383) );
  NAND4X0 U651 ( .IN1(n386), .IN2(n385), .IN3(n384), .IN4(n383), .QN(n387) );
  NOR4X0 U652 ( .IN1(input_factor_02[11]), .IN2(input_factor_02[12]), .IN3(
        n388), .IN4(n387), .QN(n389) );
  AO222X1 U653 ( .IN1(input_factor_01[31]), .IN2(n4), .IN3(input_factor_01[31]), .IN4(n393), .IN5(n392), .IN6(input_factor_02[31]), .Q(n394) );
  AND2X1 U654 ( .IN1(n562), .IN2(n394), .Q(N211) );
  MUX21X1 U655 ( .IN1(n830), .IN2(n828), .S(add_sub_result_24_), .Q(N226) );
  MUX21X1 U656 ( .IN1(n828), .IN2(n808), .S(add_sub_result_24_), .Q(N227) );
  MUX21X1 U657 ( .IN1(n808), .IN2(n800), .S(add_sub_result_24_), .Q(N228) );
  MUX21X1 U658 ( .IN1(n800), .IN2(n809), .S(add_sub_result_24_), .Q(N229) );
  MUX21X1 U659 ( .IN1(n809), .IN2(n801), .S(add_sub_result_24_), .Q(N230) );
  MUX21X1 U660 ( .IN1(n801), .IN2(n776), .S(add_sub_result_24_), .Q(N231) );
  MUX21X1 U661 ( .IN1(n776), .IN2(n768), .S(add_sub_result_24_), .Q(N232) );
  MUX21X1 U662 ( .IN1(n768), .IN2(n760), .S(add_sub_result_24_), .Q(N233) );
  MUX21X1 U663 ( .IN1(n760), .IN2(n752), .S(add_sub_result_24_), .Q(N234) );
  MUX21X1 U664 ( .IN1(n752), .IN2(n744), .S(add_sub_result_24_), .Q(N235) );
  MUX21X1 U665 ( .IN1(n744), .IN2(n736), .S(add_sub_result_24_), .Q(N236) );
  MUX21X1 U666 ( .IN1(n736), .IN2(n442), .S(add_sub_result_24_), .Q(N237) );
  MUX21X1 U667 ( .IN1(add_result[13]), .IN2(sub_result[13]), .S(n16), .Q(n447)
         );
  MUX21X1 U668 ( .IN1(n442), .IN2(n447), .S(add_sub_result_24_), .Q(N238) );
  MUX21X1 U669 ( .IN1(add_result[14]), .IN2(sub_result[14]), .S(n16), .Q(n501)
         );
  MUX21X1 U670 ( .IN1(n447), .IN2(n501), .S(add_sub_result_24_), .Q(N239) );
  MUX21X1 U671 ( .IN1(add_result[15]), .IN2(sub_result[15]), .S(n16), .Q(n456)
         );
  MUX21X1 U672 ( .IN1(n501), .IN2(n456), .S(add_sub_result_24_), .Q(N240) );
  MUX21X1 U673 ( .IN1(n456), .IN2(n396), .S(add_sub_result_24_), .Q(N241) );
  MUX21X1 U674 ( .IN1(n396), .IN2(n465), .S(add_sub_result_24_), .Q(N242) );
  MUX21X1 U675 ( .IN1(n465), .IN2(n398), .S(add_sub_result_24_), .Q(N243) );
  MUX21X1 U676 ( .IN1(n398), .IN2(n474), .S(add_sub_result_24_), .Q(N244) );
  MUX21X1 U677 ( .IN1(n474), .IN2(n399), .S(add_sub_result_24_), .Q(N245) );
  MUX21X1 U678 ( .IN1(n399), .IN2(n402), .S(add_sub_result_24_), .Q(N246) );
  MUX21X1 U679 ( .IN1(n402), .IN2(n400), .S(add_sub_result_24_), .Q(N247) );
  MUX21X1 U680 ( .IN1(n400), .IN2(n395), .S(add_sub_result_24_), .Q(N248) );
  NAND4X0 U681 ( .IN1(n496), .IN2(n485), .IN3(n489), .IN4(n487), .QN(N256) );
  INVX0 U682 ( .INP(n402), .ZN(n488) );
  NOR2X0 U683 ( .IN1(n488), .IN2(n403), .QN(n419) );
  NAND4X0 U684 ( .IN1(n496), .IN2(n483), .IN3(n489), .IN4(n491), .QN(N257) );
  NAND3X0 U685 ( .IN1(n404), .IN2(n492), .IN3(n474), .QN(n493) );
  NAND4X0 U686 ( .IN1(n496), .IN2(n485), .IN3(n493), .IN4(n483), .QN(N258) );
  NOR2X0 U687 ( .IN1(n822), .IN2(n487), .QN(N260) );
  INVX0 U688 ( .INP(n487), .ZN(n421) );
  AO22X1 U689 ( .IN1(n421), .IN2(n828), .IN3(n419), .IN4(n830), .Q(N261) );
  INVX0 U690 ( .INP(n489), .ZN(n420) );
  AO222X1 U691 ( .IN1(n830), .IN2(n420), .IN3(n828), .IN4(n419), .IN5(n808), 
        .IN6(n421), .Q(N262) );
  OA22X1 U692 ( .IN1(n814), .IN2(n489), .IN3(n822), .IN4(n493), .Q(n406) );
  OA22X1 U693 ( .IN1(n820), .IN2(n491), .IN3(n818), .IN4(n487), .Q(n405) );
  OA22X1 U694 ( .IN1(n798), .IN2(n487), .IN3(n818), .IN4(n491), .Q(n409) );
  OA22X1 U695 ( .IN1(n814), .IN2(n493), .IN3(n822), .IN4(n485), .Q(n408) );
  NAND3X0 U696 ( .IN1(n409), .IN2(n408), .IN3(n407), .QN(N264) );
  OA22X1 U697 ( .IN1(n788), .IN2(n487), .IN3(n818), .IN4(n489), .Q(n413) );
  OA22X1 U698 ( .IN1(n820), .IN2(n493), .IN3(n814), .IN4(n485), .Q(n412) );
  INVX0 U699 ( .INP(n483), .ZN(n414) );
  NAND4X0 U700 ( .IN1(n413), .IN2(n412), .IN3(n411), .IN4(n410), .QN(N265) );
  OA22X1 U701 ( .IN1(n798), .IN2(n489), .IN3(n818), .IN4(n493), .Q(n418) );
  OA22X1 U702 ( .IN1(n789), .IN2(n487), .IN3(n788), .IN4(n491), .Q(n417) );
  OA22X1 U703 ( .IN1(n820), .IN2(n485), .IN3(n822), .IN4(n496), .Q(n416) );
  NAND4X0 U704 ( .IN1(n418), .IN2(n417), .IN3(n416), .IN4(n415), .QN(N266) );
  NOR4X0 U705 ( .IN1(n421), .IN2(n420), .IN3(n419), .IN4(N258), .QN(n563) );
  OA22X1 U706 ( .IN1(n820), .IN2(n483), .IN3(n818), .IN4(n485), .Q(n425) );
  OA22X1 U707 ( .IN1(n781), .IN2(n487), .IN3(n788), .IN4(n489), .Q(n424) );
  OA22X1 U708 ( .IN1(n789), .IN2(n491), .IN3(n798), .IN4(n493), .Q(n423) );
  OA22X1 U709 ( .IN1(n814), .IN2(n496), .IN3(n822), .IN4(n838), .Q(n422) );
  NAND4X0 U710 ( .IN1(n425), .IN2(n424), .IN3(n423), .IN4(n422), .QN(N267) );
  OA22X1 U711 ( .IN1(n798), .IN2(n485), .IN3(n818), .IN4(n483), .Q(n429) );
  OA22X1 U712 ( .IN1(n773), .IN2(n487), .IN3(n789), .IN4(n489), .Q(n428) );
  OA22X1 U713 ( .IN1(n781), .IN2(n491), .IN3(n788), .IN4(n493), .Q(n427) );
  OA22X1 U714 ( .IN1(n820), .IN2(n496), .IN3(n814), .IN4(n838), .Q(n426) );
  NAND4X0 U715 ( .IN1(n429), .IN2(n428), .IN3(n427), .IN4(n426), .QN(N268) );
  OA22X1 U716 ( .IN1(n788), .IN2(n485), .IN3(n798), .IN4(n483), .Q(n433) );
  OA22X1 U717 ( .IN1(n765), .IN2(n487), .IN3(n781), .IN4(n489), .Q(n432) );
  OA22X1 U718 ( .IN1(n773), .IN2(n491), .IN3(n789), .IN4(n493), .Q(n431) );
  OA22X1 U719 ( .IN1(n820), .IN2(n838), .IN3(n818), .IN4(n496), .Q(n430) );
  NAND4X0 U720 ( .IN1(n433), .IN2(n432), .IN3(n431), .IN4(n430), .QN(N269) );
  OA22X1 U721 ( .IN1(n789), .IN2(n485), .IN3(n788), .IN4(n483), .Q(n437) );
  OA22X1 U722 ( .IN1(n773), .IN2(n489), .IN3(n757), .IN4(n487), .Q(n436) );
  OA22X1 U723 ( .IN1(n765), .IN2(n491), .IN3(n781), .IN4(n493), .Q(n435) );
  OA22X1 U724 ( .IN1(n798), .IN2(n496), .IN3(n818), .IN4(n838), .Q(n434) );
  NAND4X0 U725 ( .IN1(n437), .IN2(n436), .IN3(n435), .IN4(n434), .QN(N270) );
  OA22X1 U726 ( .IN1(n781), .IN2(n485), .IN3(n789), .IN4(n483), .Q(n441) );
  OA22X1 U727 ( .IN1(n749), .IN2(n487), .IN3(n765), .IN4(n489), .Q(n440) );
  OA22X1 U728 ( .IN1(n773), .IN2(n493), .IN3(n757), .IN4(n491), .Q(n439) );
  OA22X1 U729 ( .IN1(n788), .IN2(n496), .IN3(n798), .IN4(n838), .Q(n438) );
  NAND4X0 U730 ( .IN1(n441), .IN2(n440), .IN3(n439), .IN4(n438), .QN(N271) );
  OA22X1 U731 ( .IN1(n773), .IN2(n485), .IN3(n781), .IN4(n483), .Q(n446) );
  OA22X1 U732 ( .IN1(n741), .IN2(n487), .IN3(n757), .IN4(n489), .Q(n445) );
  OA22X1 U733 ( .IN1(n749), .IN2(n491), .IN3(n765), .IN4(n493), .Q(n444) );
  OA22X1 U734 ( .IN1(n789), .IN2(n496), .IN3(n788), .IN4(n838), .Q(n443) );
  NAND4X0 U735 ( .IN1(n446), .IN2(n445), .IN3(n444), .IN4(n443), .QN(N272) );
  OA22X1 U736 ( .IN1(n773), .IN2(n483), .IN3(n765), .IN4(n485), .Q(n451) );
  OA22X1 U737 ( .IN1(n749), .IN2(n489), .IN3(n730), .IN4(n487), .Q(n450) );
  OA22X1 U738 ( .IN1(n741), .IN2(n491), .IN3(n757), .IN4(n493), .Q(n449) );
  OA22X1 U739 ( .IN1(n781), .IN2(n496), .IN3(n789), .IN4(n838), .Q(n448) );
  NAND4X0 U740 ( .IN1(n451), .IN2(n450), .IN3(n449), .IN4(n448), .QN(N273) );
  OA22X1 U741 ( .IN1(n757), .IN2(n485), .IN3(n765), .IN4(n483), .Q(n455) );
  INVX0 U742 ( .INP(n501), .ZN(n495) );
  OA22X1 U743 ( .IN1(n495), .IN2(n487), .IN3(n741), .IN4(n489), .Q(n454) );
  OA22X1 U744 ( .IN1(n749), .IN2(n493), .IN3(n730), .IN4(n491), .Q(n453) );
  OA22X1 U745 ( .IN1(n773), .IN2(n496), .IN3(n781), .IN4(n838), .Q(n452) );
  NAND4X0 U746 ( .IN1(n455), .IN2(n454), .IN3(n453), .IN4(n452), .QN(N274) );
  OA22X1 U747 ( .IN1(n749), .IN2(n485), .IN3(n757), .IN4(n483), .Q(n460) );
  OA22X1 U748 ( .IN1(n565), .IN2(n487), .IN3(n730), .IN4(n489), .Q(n459) );
  OA22X1 U749 ( .IN1(n495), .IN2(n491), .IN3(n741), .IN4(n493), .Q(n458) );
  OA22X1 U750 ( .IN1(n773), .IN2(n838), .IN3(n765), .IN4(n496), .Q(n457) );
  NAND4X0 U751 ( .IN1(n460), .IN2(n459), .IN3(n458), .IN4(n457), .QN(N275) );
  OA22X1 U752 ( .IN1(n741), .IN2(n485), .IN3(n749), .IN4(n483), .Q(n464) );
  OA22X1 U753 ( .IN1(n495), .IN2(n489), .IN3(n484), .IN4(n487), .Q(n463) );
  OA22X1 U754 ( .IN1(n565), .IN2(n491), .IN3(n730), .IN4(n493), .Q(n462) );
  OA22X1 U755 ( .IN1(n757), .IN2(n496), .IN3(n765), .IN4(n838), .Q(n461) );
  NAND4X0 U756 ( .IN1(n464), .IN2(n463), .IN3(n462), .IN4(n461), .QN(N276) );
  OA22X1 U757 ( .IN1(n741), .IN2(n483), .IN3(n730), .IN4(n485), .Q(n469) );
  INVX0 U758 ( .INP(n465), .ZN(n486) );
  OA22X1 U759 ( .IN1(n565), .IN2(n489), .IN3(n486), .IN4(n487), .Q(n468) );
  OA22X1 U760 ( .IN1(n495), .IN2(n493), .IN3(n484), .IN4(n491), .Q(n467) );
  OA22X1 U761 ( .IN1(n749), .IN2(n496), .IN3(n757), .IN4(n838), .Q(n466) );
  NAND4X0 U762 ( .IN1(n469), .IN2(n468), .IN3(n467), .IN4(n466), .QN(N277) );
  OA22X1 U763 ( .IN1(n495), .IN2(n485), .IN3(n730), .IN4(n483), .Q(n473) );
  OA22X1 U764 ( .IN1(n494), .IN2(n487), .IN3(n484), .IN4(n489), .Q(n472) );
  OA22X1 U765 ( .IN1(n565), .IN2(n493), .IN3(n486), .IN4(n491), .Q(n471) );
  OA22X1 U766 ( .IN1(n741), .IN2(n496), .IN3(n749), .IN4(n838), .Q(n470) );
  NAND4X0 U767 ( .IN1(n473), .IN2(n472), .IN3(n471), .IN4(n470), .QN(N278) );
  OA22X1 U768 ( .IN1(n565), .IN2(n485), .IN3(n495), .IN4(n483), .Q(n478) );
  INVX0 U769 ( .INP(n474), .ZN(n490) );
  OA22X1 U770 ( .IN1(n486), .IN2(n489), .IN3(n490), .IN4(n487), .Q(n477) );
  OA22X1 U771 ( .IN1(n494), .IN2(n491), .IN3(n484), .IN4(n493), .Q(n476) );
  OA22X1 U772 ( .IN1(n741), .IN2(n838), .IN3(n730), .IN4(n496), .Q(n475) );
  NAND4X0 U773 ( .IN1(n478), .IN2(n477), .IN3(n476), .IN4(n475), .QN(N279) );
  OA22X1 U774 ( .IN1(n565), .IN2(n483), .IN3(n484), .IN4(n485), .Q(n482) );
  OA22X1 U775 ( .IN1(n494), .IN2(n489), .IN3(n492), .IN4(n487), .Q(n481) );
  OA22X1 U776 ( .IN1(n486), .IN2(n493), .IN3(n490), .IN4(n491), .Q(n480) );
  OA22X1 U777 ( .IN1(n495), .IN2(n496), .IN3(n730), .IN4(n838), .Q(n479) );
  NAND4X0 U778 ( .IN1(n482), .IN2(n481), .IN3(n480), .IN4(n479), .QN(N280) );
  OA22X1 U779 ( .IN1(n486), .IN2(n485), .IN3(n484), .IN4(n483), .Q(n500) );
  OA22X1 U780 ( .IN1(n490), .IN2(n489), .IN3(n488), .IN4(n487), .Q(n499) );
  OA22X1 U781 ( .IN1(n494), .IN2(n493), .IN3(n492), .IN4(n491), .Q(n498) );
  OA22X1 U782 ( .IN1(n565), .IN2(n496), .IN3(n495), .IN4(n838), .Q(n497) );
  NAND4X0 U783 ( .IN1(n500), .IN2(n499), .IN3(n498), .IN4(n497), .QN(N281) );
  NAND3X0 U784 ( .IN1(n501), .IN2(n514), .IN3(n565), .QN(n729) );
  AO22X1 U785 ( .IN1(n512), .IN2(add_result[12]), .IN3(n510), .IN4(
        sub_result[12]), .Q(n502) );
  INVX0 U786 ( .INP(n729), .ZN(n508) );
  NOR3X0 U787 ( .IN1(n503), .IN2(add_result[14]), .IN3(add_result[15]), .QN(
        n505) );
  NOR3X0 U788 ( .IN1(sub_result[14]), .IN2(sub_result[15]), .IN3(n17), .QN(
        n504) );
  AO22X1 U789 ( .IN1(n505), .IN2(add_result[13]), .IN3(n504), .IN4(
        sub_result[13]), .Q(n506) );
  NOR2X0 U790 ( .IN1(n508), .IN2(n507), .QN(N308) );
  INVX0 U791 ( .INP(add_result[12]), .ZN(n511) );
  INVX0 U792 ( .INP(sub_result[12]), .ZN(n509) );
  AO22X1 U793 ( .IN1(n512), .IN2(n511), .IN3(n510), .IN4(n509), .Q(n513) );
  NAND3X0 U794 ( .IN1(n514), .IN2(n736), .IN3(n513), .QN(n823) );
  NAND4X0 U795 ( .IN1(N308), .IN2(n823), .IN3(n806), .IN4(n797), .QN(n790) );
  NAND4X0 U796 ( .IN1(n806), .IN2(n729), .IN3(n735), .IN4(n790), .QN(N306) );
  NAND4X0 U797 ( .IN1(n797), .IN2(n728), .IN3(n735), .IN4(n790), .QN(N307) );
  AO22X1 U798 ( .IN1(n716), .IN2(exponent_factor_12[0]), .IN3(n834), .IN4(
        exponent_factor_21[0]), .Q(N34) );
  NAND3X0 U799 ( .IN1(n818), .IN2(n524), .IN3(n808), .QN(n537) );
  NAND3X0 U800 ( .IN1(n788), .IN2(n516), .IN3(n809), .QN(n532) );
  NAND3X0 U801 ( .IN1(n781), .IN2(n517), .IN3(n776), .QN(n533) );
  NAND3X0 U802 ( .IN1(n820), .IN2(n814), .IN3(n818), .QN(n515) );
  AND2X1 U803 ( .IN1(n532), .IN2(n534), .Q(n519) );
  NAND4X0 U804 ( .IN1(n521), .IN2(n519), .IN3(n533), .IN4(n535), .QN(n520) );
  NAND4X0 U805 ( .IN1(n537), .IN2(n532), .IN3(n533), .IN4(n520), .QN(N346) );
  NAND3X0 U806 ( .IN1(n519), .IN2(n536), .IN3(n520), .QN(N347) );
  NOR2X0 U807 ( .IN1(n822), .IN2(n535), .QN(N349) );
  AO22X1 U808 ( .IN1(n716), .IN2(exponent_factor_12[1]), .IN3(n834), .IN4(
        exponent_factor_21[1]), .Q(N35) );
  OAI22X1 U809 ( .IN1(n814), .IN2(n535), .IN3(n822), .IN4(n533), .QN(N350) );
  OAI222X1 U810 ( .IN1(n534), .IN2(n822), .IN3(n533), .IN4(n814), .IN5(n535), 
        .IN6(n820), .QN(N351) );
  OA22X1 U811 ( .IN1(n820), .IN2(n533), .IN3(n818), .IN4(n535), .Q(n523) );
  OA22X1 U812 ( .IN1(n814), .IN2(n534), .IN3(n822), .IN4(n532), .Q(n522) );
  OA22X1 U813 ( .IN1(n798), .IN2(n535), .IN3(n818), .IN4(n533), .Q(n527) );
  OA22X1 U814 ( .IN1(n820), .IN2(n534), .IN3(n814), .IN4(n532), .Q(n526) );
  AND2X1 U815 ( .IN1(n524), .IN2(n800), .Q(n538) );
  NAND3X0 U816 ( .IN1(n527), .IN2(n526), .IN3(n525), .QN(N353) );
  OA22X1 U817 ( .IN1(n788), .IN2(n535), .IN3(n798), .IN4(n533), .Q(n531) );
  OA22X1 U818 ( .IN1(n820), .IN2(n532), .IN3(n822), .IN4(n537), .Q(n530) );
  OR2X1 U819 ( .IN1(n534), .IN2(n818), .Q(n528) );
  NAND4X0 U820 ( .IN1(n531), .IN2(n530), .IN3(n529), .IN4(n528), .QN(N354) );
  OA22X1 U821 ( .IN1(n788), .IN2(n533), .IN3(n818), .IN4(n532), .Q(n542) );
  OA22X1 U822 ( .IN1(n789), .IN2(n535), .IN3(n798), .IN4(n534), .Q(n541) );
  OA22X1 U823 ( .IN1(n814), .IN2(n537), .IN3(n822), .IN4(n536), .Q(n540) );
  NAND4X0 U824 ( .IN1(n542), .IN2(n541), .IN3(n540), .IN4(n539), .QN(N355) );
  AO22X1 U825 ( .IN1(n716), .IN2(exponent_factor_12[2]), .IN3(n834), .IN4(
        exponent_factor_21[2]), .Q(N36) );
  AO22X1 U826 ( .IN1(n716), .IN2(exponent_factor_12[3]), .IN3(n834), .IN4(
        exponent_factor_21[3]), .Q(N37) );
  AO22X1 U827 ( .IN1(n716), .IN2(exponent_factor_12[4]), .IN3(n834), .IN4(
        exponent_factor_21[4]), .Q(N38) );
  NAND4X0 U828 ( .IN1(n633), .IN2(n629), .IN3(n625), .IN4(n621), .QN(n547) );
  NAND4X0 U829 ( .IN1(n617), .IN2(n613), .IN3(n543), .IN4(n609), .QN(n546) );
  NAND4X0 U830 ( .IN1(n674), .IN2(n671), .IN3(n665), .IN4(n659), .QN(n545) );
  NAND4X0 U831 ( .IN1(n653), .IN2(n647), .IN3(n641), .IN4(n637), .QN(n544) );
  NOR4X0 U832 ( .IN1(n547), .IN2(n546), .IN3(n545), .IN4(n544), .QN(n557) );
  NAND4X0 U833 ( .IN1(n549), .IN2(n601), .IN3(n589), .IN4(n548), .QN(n555) );
  INVX0 U834 ( .INP(input_factor_01[23]), .ZN(n558) );
  NAND4X0 U835 ( .IN1(n550), .IN2(n558), .IN3(n595), .IN4(n583), .QN(n554) );
  NAND4X0 U836 ( .IN1(n717), .IN2(n710), .IN3(n704), .IN4(n698), .QN(n553) );
  NAND4X0 U837 ( .IN1(n551), .IN2(n692), .IN3(n686), .IN4(n680), .QN(n552) );
  NOR4X0 U838 ( .IN1(n555), .IN2(n554), .IN3(n553), .IN4(n552), .QN(n556) );
  OA22X1 U839 ( .IN1(n559), .IN2(n718), .IN3(n18), .IN4(n558), .Q(n574) );
  INVX0 U840 ( .INP(n790), .ZN(n560) );
  OA21X1 U841 ( .IN1(n773), .IN2(n561), .IN3(n560), .Q(n567) );
  OA21X1 U842 ( .IN1(n565), .IN2(n564), .IN3(n563), .Q(n566) );
  AOI22X1 U843 ( .IN1(n721), .IN2(add_output_exponent_w3[0]), .IN3(n720), 
        .IN4(add_output_exponent_w2[0]), .QN(n573) );
  INVX0 U844 ( .INP(n569), .ZN(n568) );
  AND4X1 U845 ( .IN1(n570), .IN2(n568), .IN3(n567), .IN4(n566), .Q(n722) );
  NAND4X0 U846 ( .IN1(n574), .IN2(n573), .IN3(n572), .IN4(n571), .QN(N380) );
  AOI22X1 U847 ( .IN1(input_factor_02[24]), .IN2(n19), .IN3(n4), .IN4(
        input_factor_01[24]), .QN(n578) );
  AOI22X1 U848 ( .IN1(n721), .IN2(add_output_exponent_w3[1]), .IN3(n720), 
        .IN4(add_output_exponent_w2[1]), .QN(n577) );
  NAND4X0 U849 ( .IN1(n578), .IN2(n577), .IN3(n576), .IN4(n575), .QN(N381) );
  AOI22X1 U850 ( .IN1(input_factor_02[25]), .IN2(n19), .IN3(n4), .IN4(
        input_factor_01[25]), .QN(n582) );
  AOI22X1 U851 ( .IN1(n721), .IN2(add_output_exponent_w3[2]), .IN3(n720), 
        .IN4(add_output_exponent_w2[2]), .QN(n581) );
  NAND4X0 U852 ( .IN1(n582), .IN2(n581), .IN3(n580), .IN4(n579), .QN(N382) );
  OA22X1 U853 ( .IN1(n584), .IN2(n718), .IN3(n18), .IN4(n583), .Q(n588) );
  AOI22X1 U854 ( .IN1(n721), .IN2(add_output_exponent_w3[3]), .IN3(n720), 
        .IN4(add_output_exponent_w2[3]), .QN(n587) );
  NAND4X0 U855 ( .IN1(n588), .IN2(n587), .IN3(n586), .IN4(n585), .QN(N383) );
  OA22X1 U856 ( .IN1(n590), .IN2(n718), .IN3(n18), .IN4(n589), .Q(n594) );
  AOI22X1 U857 ( .IN1(n721), .IN2(add_output_exponent_w3[4]), .IN3(n720), 
        .IN4(add_output_exponent_w2[4]), .QN(n593) );
  NAND4X0 U858 ( .IN1(n594), .IN2(n593), .IN3(n592), .IN4(n591), .QN(N384) );
  OA22X1 U859 ( .IN1(n596), .IN2(n718), .IN3(n18), .IN4(n595), .Q(n600) );
  AOI22X1 U860 ( .IN1(n721), .IN2(add_output_exponent_w3[5]), .IN3(n720), 
        .IN4(add_output_exponent_w2[5]), .QN(n599) );
  NAND4X0 U861 ( .IN1(n600), .IN2(n599), .IN3(n598), .IN4(n597), .QN(N385) );
  OA22X1 U862 ( .IN1(n602), .IN2(n718), .IN3(n18), .IN4(n601), .Q(n606) );
  AOI22X1 U863 ( .IN1(n721), .IN2(add_output_exponent_w3[6]), .IN3(n720), 
        .IN4(add_output_exponent_w2[6]), .QN(n605) );
  NAND4X0 U864 ( .IN1(n606), .IN2(n605), .IN3(n604), .IN4(n603), .QN(N386) );
  AO22X1 U866 ( .IN1(n4), .IN2(input_factor_01[30]), .IN3(n723), .IN4(
        add_output_exponent_w1[7]), .Q(n608) );
  AO22X1 U867 ( .IN1(n721), .IN2(add_output_exponent_w3[7]), .IN3(n720), .IN4(
        add_output_exponent_w2[7]), .Q(n607) );
  AO222X1 U868 ( .IN1(input_factor_02[0]), .IN2(n19), .IN3(input_factor_01[0]), 
        .IN4(n4), .IN5(n723), .IN6(pre_sig_res_01[0]), .Q(N388) );
  AOI22X1 U869 ( .IN1(n720), .IN2(pre_sig_res_02[1]), .IN3(n723), .IN4(
        pre_sig_res_01[1]), .QN(n612) );
  OA22X1 U870 ( .IN1(n610), .IN2(n718), .IN3(n18), .IN4(n609), .Q(n611) );
  AO22X1 U871 ( .IN1(n716), .IN2(exponent_factor_12[5]), .IN3(n834), .IN4(
        exponent_factor_21[5]), .Q(N39) );
  AOI22X1 U872 ( .IN1(n720), .IN2(pre_sig_res_02[2]), .IN3(n723), .IN4(
        pre_sig_res_01[2]), .QN(n616) );
  OA22X1 U873 ( .IN1(n614), .IN2(n718), .IN3(n18), .IN4(n613), .Q(n615) );
  AOI22X1 U874 ( .IN1(n720), .IN2(pre_sig_res_02[3]), .IN3(n723), .IN4(
        pre_sig_res_01[3]), .QN(n620) );
  OA22X1 U875 ( .IN1(n618), .IN2(n718), .IN3(n18), .IN4(n617), .Q(n619) );
  AOI22X1 U876 ( .IN1(n720), .IN2(pre_sig_res_02[4]), .IN3(n723), .IN4(
        pre_sig_res_01[4]), .QN(n624) );
  OA22X1 U877 ( .IN1(n622), .IN2(n718), .IN3(n18), .IN4(n621), .Q(n623) );
  AOI22X1 U878 ( .IN1(n720), .IN2(pre_sig_res_02[5]), .IN3(n723), .IN4(
        pre_sig_res_01[5]), .QN(n628) );
  OA22X1 U879 ( .IN1(n626), .IN2(n718), .IN3(n18), .IN4(n625), .Q(n627) );
  AOI22X1 U880 ( .IN1(n720), .IN2(pre_sig_res_02[6]), .IN3(n723), .IN4(
        pre_sig_res_01[6]), .QN(n632) );
  OA22X1 U881 ( .IN1(n630), .IN2(n718), .IN3(n18), .IN4(n629), .Q(n631) );
  AOI22X1 U882 ( .IN1(n720), .IN2(pre_sig_res_02[7]), .IN3(n723), .IN4(
        pre_sig_res_01[7]), .QN(n636) );
  OA22X1 U883 ( .IN1(n634), .IN2(n718), .IN3(n18), .IN4(n633), .Q(n635) );
  AOI22X1 U884 ( .IN1(n720), .IN2(pre_sig_res_02[8]), .IN3(n723), .IN4(
        pre_sig_res_01[8]), .QN(n640) );
  OA22X1 U885 ( .IN1(n638), .IN2(n718), .IN3(n18), .IN4(n637), .Q(n639) );
  OA22X1 U886 ( .IN1(n642), .IN2(n718), .IN3(n18), .IN4(n641), .Q(n646) );
  NAND4X0 U887 ( .IN1(n646), .IN2(n645), .IN3(n644), .IN4(n643), .QN(N397) );
  OA22X1 U888 ( .IN1(n648), .IN2(n718), .IN3(n18), .IN4(n647), .Q(n652) );
  NAND4X0 U889 ( .IN1(n652), .IN2(n651), .IN3(n650), .IN4(n649), .QN(N398) );
  OA22X1 U890 ( .IN1(n654), .IN2(n718), .IN3(n18), .IN4(n653), .Q(n658) );
  NAND4X0 U891 ( .IN1(n658), .IN2(n657), .IN3(n656), .IN4(n655), .QN(N399) );
  AO22X1 U892 ( .IN1(n716), .IN2(exponent_factor_12[6]), .IN3(n834), .IN4(
        exponent_factor_21[6]), .Q(N40) );
  OA22X1 U893 ( .IN1(n660), .IN2(n718), .IN3(n18), .IN4(n659), .Q(n664) );
  NAND4X0 U894 ( .IN1(n664), .IN2(n663), .IN3(n662), .IN4(n661), .QN(N400) );
  OA22X1 U895 ( .IN1(n666), .IN2(n718), .IN3(n18), .IN4(n665), .Q(n670) );
  NAND4X0 U896 ( .IN1(n670), .IN2(n669), .IN3(n668), .IN4(n667), .QN(N401) );
  NOR2X0 U897 ( .IN1(n18), .IN2(n671), .QN(n673) );
  AO22X1 U898 ( .IN1(n721), .IN2(pre_sig_res_03[14]), .IN3(n720), .IN4(
        pre_sig_res_02[14]), .Q(n672) );
  OA22X1 U899 ( .IN1(n675), .IN2(n718), .IN3(n18), .IN4(n674), .Q(n679) );
  NAND4X0 U900 ( .IN1(n679), .IN2(n678), .IN3(n677), .IN4(n676), .QN(N403) );
  OA22X1 U901 ( .IN1(n681), .IN2(n718), .IN3(n18), .IN4(n680), .Q(n685) );
  AOI22X1 U902 ( .IN1(n721), .IN2(pre_sig_res_03[16]), .IN3(n720), .IN4(
        pre_sig_res_02[16]), .QN(n684) );
  NAND4X0 U903 ( .IN1(n685), .IN2(n684), .IN3(n683), .IN4(n682), .QN(N404) );
  OA22X1 U904 ( .IN1(n687), .IN2(n718), .IN3(n18), .IN4(n686), .Q(n691) );
  AOI22X1 U905 ( .IN1(n721), .IN2(pre_sig_res_03[17]), .IN3(n720), .IN4(
        pre_sig_res_02[17]), .QN(n690) );
  NAND4X0 U906 ( .IN1(n691), .IN2(n690), .IN3(n689), .IN4(n688), .QN(N405) );
  OA22X1 U907 ( .IN1(n693), .IN2(n718), .IN3(n18), .IN4(n692), .Q(n697) );
  AOI22X1 U908 ( .IN1(n721), .IN2(pre_sig_res_03[18]), .IN3(n720), .IN4(
        pre_sig_res_02[18]), .QN(n696) );
  NAND4X0 U909 ( .IN1(n697), .IN2(n696), .IN3(n695), .IN4(n694), .QN(N406) );
  OA22X1 U910 ( .IN1(n699), .IN2(n718), .IN3(n18), .IN4(n698), .Q(n703) );
  AOI22X1 U911 ( .IN1(n721), .IN2(pre_sig_res_03[19]), .IN3(n720), .IN4(
        pre_sig_res_02[19]), .QN(n702) );
  NAND4X0 U912 ( .IN1(n703), .IN2(n702), .IN3(n701), .IN4(n700), .QN(N407) );
  OA22X1 U913 ( .IN1(n705), .IN2(n718), .IN3(n18), .IN4(n704), .Q(n709) );
  AOI22X1 U914 ( .IN1(n721), .IN2(pre_sig_res_03[20]), .IN3(n720), .IN4(
        pre_sig_res_02[20]), .QN(n708) );
  NAND4X0 U915 ( .IN1(n709), .IN2(n708), .IN3(n707), .IN4(n706), .QN(N408) );
  OA22X1 U916 ( .IN1(n711), .IN2(n718), .IN3(n18), .IN4(n710), .Q(n715) );
  AOI22X1 U917 ( .IN1(n721), .IN2(pre_sig_res_03[21]), .IN3(n720), .IN4(
        pre_sig_res_02[21]), .QN(n714) );
  NAND4X0 U918 ( .IN1(n715), .IN2(n714), .IN3(n713), .IN4(n712), .QN(N409) );
  AO22X1 U919 ( .IN1(n716), .IN2(exponent_factor_12[7]), .IN3(n834), .IN4(
        exponent_factor_21[7]), .Q(N41) );
  OA22X1 U920 ( .IN1(n719), .IN2(n718), .IN3(n18), .IN4(n717), .Q(n727) );
  AOI22X1 U921 ( .IN1(n721), .IN2(pre_sig_res_03[22]), .IN3(n720), .IN4(
        pre_sig_res_02[22]), .QN(n726) );
  NAND4X0 U922 ( .IN1(n727), .IN2(n726), .IN3(n725), .IN4(n724), .QN(N410) );
  NOR2X0 U923 ( .IN1(n861), .IN2(n728), .QN(n829) );
  NOR2X0 U924 ( .IN1(n729), .IN2(n861), .QN(n831) );
  OA22X1 U925 ( .IN1(n741), .IN2(n819), .IN3(n730), .IN4(n817), .Q(n740) );
  OA22X1 U926 ( .IN1(n757), .IN2(n823), .IN3(n781), .IN4(n790), .Q(n734) );
  INVX0 U927 ( .INP(rst_n), .ZN(n832) );
  NAND3X0 U928 ( .IN1(n732), .IN2(n752), .IN3(n731), .QN(n733) );
  OA22X1 U929 ( .IN1(n861), .IN2(n734), .IN3(n832), .IN4(n733), .Q(n739) );
  NAND4X0 U930 ( .IN1(n740), .IN2(n739), .IN3(n738), .IN4(n737), .QN(n860) );
  OA22X1 U931 ( .IN1(n741), .IN2(n817), .IN3(n749), .IN4(n819), .Q(n748) );
  OA22X1 U932 ( .IN1(n781), .IN2(n797), .IN3(n789), .IN4(n790), .Q(n743) );
  OA22X1 U933 ( .IN1(n773), .IN2(n806), .IN3(n765), .IN4(n823), .Q(n742) );
  AO21X1 U934 ( .IN1(n743), .IN2(n742), .IN3(n861), .Q(n747) );
  NAND4X0 U935 ( .IN1(n748), .IN2(n747), .IN3(n746), .IN4(n745), .QN(n859) );
  OA22X1 U936 ( .IN1(n749), .IN2(n817), .IN3(n757), .IN4(n819), .Q(n756) );
  OA22X1 U937 ( .IN1(n789), .IN2(n797), .IN3(n788), .IN4(n790), .Q(n751) );
  OA22X1 U938 ( .IN1(n773), .IN2(n823), .IN3(n781), .IN4(n806), .Q(n750) );
  AO21X1 U939 ( .IN1(n751), .IN2(n750), .IN3(n861), .Q(n755) );
  NAND4X0 U940 ( .IN1(n756), .IN2(n755), .IN3(n754), .IN4(n753), .QN(n858) );
  OA22X1 U941 ( .IN1(n757), .IN2(n817), .IN3(n765), .IN4(n819), .Q(n764) );
  OA22X1 U942 ( .IN1(n788), .IN2(n797), .IN3(n798), .IN4(n790), .Q(n759) );
  OA22X1 U943 ( .IN1(n781), .IN2(n823), .IN3(n789), .IN4(n806), .Q(n758) );
  AO21X1 U944 ( .IN1(n759), .IN2(n758), .IN3(n861), .Q(n763) );
  NAND4X0 U945 ( .IN1(n764), .IN2(n763), .IN3(n762), .IN4(n761), .QN(n857) );
  OA22X1 U946 ( .IN1(n773), .IN2(n819), .IN3(n765), .IN4(n817), .Q(n772) );
  OA22X1 U947 ( .IN1(n798), .IN2(n797), .IN3(n818), .IN4(n790), .Q(n767) );
  OA22X1 U948 ( .IN1(n789), .IN2(n823), .IN3(n788), .IN4(n806), .Q(n766) );
  AO21X1 U949 ( .IN1(n767), .IN2(n766), .IN3(n861), .Q(n771) );
  NAND4X0 U950 ( .IN1(n772), .IN2(n771), .IN3(n770), .IN4(n769), .QN(n856) );
  OA22X1 U951 ( .IN1(n773), .IN2(n817), .IN3(n781), .IN4(n819), .Q(n780) );
  OA22X1 U952 ( .IN1(n820), .IN2(n790), .IN3(n818), .IN4(n797), .Q(n775) );
  OA22X1 U953 ( .IN1(n788), .IN2(n823), .IN3(n798), .IN4(n806), .Q(n774) );
  AO21X1 U954 ( .IN1(n775), .IN2(n774), .IN3(n861), .Q(n779) );
  NAND4X0 U955 ( .IN1(n780), .IN2(n779), .IN3(n778), .IN4(n777), .QN(n855) );
  OA22X1 U956 ( .IN1(n781), .IN2(n817), .IN3(n789), .IN4(n819), .Q(n787) );
  OA22X1 U957 ( .IN1(n820), .IN2(n797), .IN3(n814), .IN4(n790), .Q(n783) );
  OA22X1 U958 ( .IN1(n798), .IN2(n823), .IN3(n818), .IN4(n806), .Q(n782) );
  AO21X1 U959 ( .IN1(n783), .IN2(n782), .IN3(n861), .Q(n786) );
  NAND4X0 U960 ( .IN1(n787), .IN2(n786), .IN3(n785), .IN4(n784), .QN(n854) );
  OA22X1 U961 ( .IN1(n789), .IN2(n817), .IN3(n788), .IN4(n819), .Q(n796) );
  OA22X1 U962 ( .IN1(n814), .IN2(n797), .IN3(n822), .IN4(n790), .Q(n792) );
  OA22X1 U963 ( .IN1(n820), .IN2(n806), .IN3(n818), .IN4(n823), .Q(n791) );
  AO21X1 U964 ( .IN1(n792), .IN2(n791), .IN3(n861), .Q(n795) );
  NAND4X0 U965 ( .IN1(n796), .IN2(n795), .IN3(n794), .IN4(n793), .QN(n853) );
  OA222X1 U966 ( .IN1(n823), .IN2(n820), .IN3(n797), .IN4(n822), .IN5(n806), 
        .IN6(n814), .Q(n799) );
  OA22X1 U967 ( .IN1(n861), .IN2(n799), .IN3(n798), .IN4(n819), .Q(n805) );
  NAND4X0 U968 ( .IN1(n805), .IN2(n804), .IN3(n803), .IN4(n802), .QN(n852) );
  OA22X1 U969 ( .IN1(n814), .IN2(n823), .IN3(n822), .IN4(n806), .Q(n807) );
  OA22X1 U970 ( .IN1(n818), .IN2(n819), .IN3(n807), .IN4(n832), .Q(n813) );
  NAND4X0 U971 ( .IN1(n813), .IN2(n812), .IN3(n811), .IN4(n810), .QN(n851) );
  AOI22X1 U972 ( .IN1(pre_sig_res_03[11]), .IN2(n832), .IN3(n821), .IN4(n830), 
        .QN(n816) );
  OA22X1 U973 ( .IN1(n820), .IN2(n817), .IN3(n814), .IN4(n819), .Q(n815) );
  OA22X1 U974 ( .IN1(n820), .IN2(n819), .IN3(n818), .IN4(n817), .Q(n827) );
  OR3X1 U975 ( .IN1(n823), .IN2(n832), .IN3(n822), .Q(n825) );
  NAND4X0 U976 ( .IN1(n827), .IN2(n826), .IN3(n825), .IN4(n824), .QN(n849) );
  AO222X1 U977 ( .IN1(n830), .IN2(n829), .IN3(n828), .IN4(n831), .IN5(n832), 
        .IN6(pre_sig_res_03[10]), .Q(n848) );
  AO22X1 U978 ( .IN1(pre_sig_res_03[9]), .IN2(n832), .IN3(n831), .IN4(n830), 
        .Q(n847) );
  AO222X1 U979 ( .IN1(input_factor_02[23]), .IN2(n836), .IN3(
        input_factor_01[23]), .IN4(n835), .IN5(larger_exponent[0]), .IN6(n861), 
        .Q(n846) );
  AO222X1 U980 ( .IN1(input_factor_02[24]), .IN2(n836), .IN3(
        input_factor_01[24]), .IN4(n835), .IN5(n861), .IN6(larger_exponent[1]), 
        .Q(n845) );
  AO222X1 U981 ( .IN1(input_factor_02[25]), .IN2(n836), .IN3(
        input_factor_01[25]), .IN4(n835), .IN5(n861), .IN6(larger_exponent[2]), 
        .Q(n844) );
  AO222X1 U982 ( .IN1(input_factor_02[26]), .IN2(n836), .IN3(
        input_factor_01[26]), .IN4(n835), .IN5(n861), .IN6(larger_exponent[3]), 
        .Q(n843) );
  AO222X1 U983 ( .IN1(input_factor_02[27]), .IN2(n836), .IN3(
        input_factor_01[27]), .IN4(n835), .IN5(n861), .IN6(larger_exponent[4]), 
        .Q(n842) );
  AO222X1 U984 ( .IN1(input_factor_02[28]), .IN2(n836), .IN3(
        input_factor_01[28]), .IN4(n835), .IN5(n861), .IN6(larger_exponent[5]), 
        .Q(n841) );
  AO222X1 U985 ( .IN1(input_factor_02[29]), .IN2(n836), .IN3(
        input_factor_01[29]), .IN4(n835), .IN5(n861), .IN6(larger_exponent[6]), 
        .Q(n840) );
endmodule


module add_481 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_482 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_483 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_484 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_485 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_486 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_487 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_488 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_489 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_490 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_491 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_492 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_493 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_494 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_495 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_496 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_497 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_498 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_499 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_500 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_501 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_502 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_503 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_504 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(b), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(b), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module adder24_9 ( clk, rst_n, a, b, cin, out );
  input [23:0] a;
  input [23:0] b;
  output [24:0] out;
  input clk, rst_n, cin;
  wire   c_tmp;
  wire   [24:0] s;
  wire   [22:0] c;

  add_504 add_01 ( .s(s[0]), .a(a[0]), .b(b[0]), .ci(1'b0), .co(c[0]) );
  add_503 add_02 ( .s(s[1]), .a(a[1]), .b(b[1]), .ci(c[0]), .co(c[1]) );
  add_502 add_03 ( .s(s[2]), .a(a[2]), .b(b[2]), .ci(c[1]), .co(c[2]) );
  add_501 add_04 ( .s(s[3]), .a(a[3]), .b(b[3]), .ci(c[2]), .co(c[3]) );
  add_500 add_05 ( .s(s[4]), .a(a[4]), .b(b[4]), .ci(c[3]), .co(c[4]) );
  add_499 add_06 ( .s(s[5]), .a(a[5]), .b(b[5]), .ci(c[4]), .co(c[5]) );
  add_498 add_07 ( .s(s[6]), .a(a[6]), .b(b[6]), .ci(c[5]), .co(c[6]) );
  add_497 add_08 ( .s(s[7]), .a(a[7]), .b(b[7]), .ci(c[6]), .co(c[7]) );
  add_496 add_09 ( .s(s[8]), .a(a[8]), .b(b[8]), .ci(c[7]), .co(c[8]) );
  add_495 add_10 ( .s(s[9]), .a(a[9]), .b(b[9]), .ci(c[8]), .co(c[9]) );
  add_494 add_11 ( .s(s[10]), .a(a[10]), .b(b[10]), .ci(c[9]), .co(c[10]) );
  add_493 add_12 ( .s(s[11]), .a(a[11]), .b(b[11]), .ci(c_tmp), .co(c[11]) );
  add_492 add_13 ( .s(s[12]), .a(a[12]), .b(b[12]), .ci(c[11]), .co(c[12]) );
  add_491 add_14 ( .s(s[13]), .a(a[13]), .b(b[13]), .ci(c[12]), .co(c[13]) );
  add_490 add_15 ( .s(s[14]), .a(a[14]), .b(b[14]), .ci(c[13]), .co(c[14]) );
  add_489 add_16 ( .s(s[15]), .a(a[15]), .b(b[15]), .ci(c[14]), .co(c[15]) );
  add_488 add_17 ( .s(s[16]), .a(a[16]), .b(b[16]), .ci(c[15]), .co(c[16]) );
  add_487 add_18 ( .s(s[17]), .a(a[17]), .b(b[17]), .ci(c[16]), .co(c[17]) );
  add_486 add_19 ( .s(s[18]), .a(a[18]), .b(b[18]), .ci(c[17]), .co(c[18]) );
  add_485 add_20 ( .s(s[19]), .a(a[19]), .b(b[19]), .ci(c[18]), .co(c[19]) );
  add_484 add_21 ( .s(s[20]), .a(a[20]), .b(b[20]), .ci(c[19]), .co(c[20]) );
  add_483 add_22 ( .s(s[21]), .a(a[21]), .b(b[21]), .ci(c[20]), .co(c[21]) );
  add_482 add_23 ( .s(s[22]), .a(a[22]), .b(b[22]), .ci(c[21]), .co(c[22]) );
  add_481 add_24 ( .s(s[23]), .a(a[23]), .b(b[23]), .ci(c[22]), .co(s[24]) );
  DFFARX1 out_reg_10_ ( .D(s[10]), .CLK(clk), .RSTB(rst_n), .Q(out[10]) );
  DFFARX1 out_reg_9_ ( .D(s[9]), .CLK(clk), .RSTB(rst_n), .Q(out[9]) );
  DFFARX1 out_reg_8_ ( .D(s[8]), .CLK(clk), .RSTB(rst_n), .Q(out[8]) );
  DFFARX1 out_reg_7_ ( .D(s[7]), .CLK(clk), .RSTB(rst_n), .Q(out[7]) );
  DFFARX1 out_reg_6_ ( .D(s[6]), .CLK(clk), .RSTB(rst_n), .Q(out[6]) );
  DFFARX1 out_reg_5_ ( .D(s[5]), .CLK(clk), .RSTB(rst_n), .Q(out[5]) );
  DFFARX1 out_reg_4_ ( .D(s[4]), .CLK(clk), .RSTB(rst_n), .Q(out[4]) );
  DFFARX1 out_reg_3_ ( .D(s[3]), .CLK(clk), .RSTB(rst_n), .Q(out[3]) );
  DFFARX1 out_reg_2_ ( .D(s[2]), .CLK(clk), .RSTB(rst_n), .Q(out[2]) );
  DFFARX1 out_reg_1_ ( .D(s[1]), .CLK(clk), .RSTB(rst_n), .Q(out[1]) );
  DFFARX1 out_reg_0_ ( .D(s[0]), .CLK(clk), .RSTB(rst_n), .Q(out[0]) );
  DFFARX1 c_tmp_reg ( .D(c[10]), .CLK(clk), .RSTB(rst_n), .Q(c_tmp) );
  DFFARX1 out_reg_24_ ( .D(s[24]), .CLK(clk), .RSTB(rst_n), .Q(out[24]) );
  DFFARX1 out_reg_23_ ( .D(s[23]), .CLK(clk), .RSTB(rst_n), .Q(out[23]) );
  DFFARX1 out_reg_22_ ( .D(s[22]), .CLK(clk), .RSTB(rst_n), .Q(out[22]) );
  DFFARX1 out_reg_21_ ( .D(s[21]), .CLK(clk), .RSTB(rst_n), .Q(out[21]) );
  DFFARX1 out_reg_20_ ( .D(s[20]), .CLK(clk), .RSTB(rst_n), .Q(out[20]) );
  DFFARX1 out_reg_19_ ( .D(s[19]), .CLK(clk), .RSTB(rst_n), .Q(out[19]) );
  DFFARX1 out_reg_18_ ( .D(s[18]), .CLK(clk), .RSTB(rst_n), .Q(out[18]) );
  DFFARX1 out_reg_17_ ( .D(s[17]), .CLK(clk), .RSTB(rst_n), .Q(out[17]) );
  DFFARX1 out_reg_16_ ( .D(s[16]), .CLK(clk), .RSTB(rst_n), .Q(out[16]) );
  DFFARX1 out_reg_15_ ( .D(s[15]), .CLK(clk), .RSTB(rst_n), .Q(out[15]) );
  DFFARX1 out_reg_14_ ( .D(s[14]), .CLK(clk), .RSTB(rst_n), .Q(out[14]) );
  DFFARX1 out_reg_13_ ( .D(s[13]), .CLK(clk), .RSTB(rst_n), .Q(out[13]) );
  DFFARX1 out_reg_12_ ( .D(s[12]), .CLK(clk), .RSTB(rst_n), .Q(out[12]) );
  DFFARX1 out_reg_11_ ( .D(s[11]), .CLK(clk), .RSTB(rst_n), .Q(out[11]) );
endmodule


module add_505 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_506 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_507 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_508 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_509 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_510 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_511 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_512 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_513 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_514 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_515 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_516 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_517 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_518 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_519 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_520 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_521 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_522 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_523 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_524 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_525 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_526 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_527 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_528 ( s, a, ci, co, b_BAR );
  input a, ci, b_BAR;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(b_BAR), .IN2(n1), .QN(co) );
  INVX0 U2 ( .INP(a), .ZN(n1) );
  MUX21X1 U3 ( .IN1(a), .IN2(n1), .S(b_BAR), .Q(s) );
endmodule


module adder24_10 ( clk, rst_n, a, b, cin, out );
  input [23:0] a;
  input [23:0] b;
  output [24:0] out;
  input clk, rst_n, cin;
  wire   c_tmp, n_1_net_, n_2_net_, n_3_net_, n_4_net_, n_5_net_, n_6_net_,
         n_7_net_, n_8_net_, n_9_net_, n_10_net_, n_11_net_, n_12_net_,
         n_13_net_, n_14_net_, n_15_net_, n_16_net_, n_17_net_, n_18_net_,
         n_19_net_, n_20_net_, n_21_net_, n_22_net_, n_23_net_;
  wire   [24:0] s;
  wire   [23:0] c;

  add_528 add_01 ( .s(s[0]), .a(a[0]), .ci(1'b1), .co(c[0]), .b_BAR(b[0]) );
  add_527 add_02 ( .s(s[1]), .a(a[1]), .b(n_1_net_), .ci(c[0]), .co(c[1]) );
  add_526 add_03 ( .s(s[2]), .a(a[2]), .b(n_2_net_), .ci(c[1]), .co(c[2]) );
  add_525 add_04 ( .s(s[3]), .a(a[3]), .b(n_3_net_), .ci(c[2]), .co(c[3]) );
  add_524 add_05 ( .s(s[4]), .a(a[4]), .b(n_4_net_), .ci(c[3]), .co(c[4]) );
  add_523 add_06 ( .s(s[5]), .a(a[5]), .b(n_5_net_), .ci(c[4]), .co(c[5]) );
  add_522 add_07 ( .s(s[6]), .a(a[6]), .b(n_6_net_), .ci(c[5]), .co(c[6]) );
  add_521 add_08 ( .s(s[7]), .a(a[7]), .b(n_7_net_), .ci(c[6]), .co(c[7]) );
  add_520 add_09 ( .s(s[8]), .a(a[8]), .b(n_8_net_), .ci(c[7]), .co(c[8]) );
  add_519 add_10 ( .s(s[9]), .a(a[9]), .b(n_9_net_), .ci(c[8]), .co(c[9]) );
  add_518 add_11 ( .s(s[10]), .a(a[10]), .b(n_10_net_), .ci(c[9]), .co(c[10])
         );
  add_517 add_12 ( .s(s[11]), .a(a[11]), .b(n_11_net_), .ci(c_tmp), .co(c[11])
         );
  add_516 add_13 ( .s(s[12]), .a(a[12]), .b(n_12_net_), .ci(c[11]), .co(c[12])
         );
  add_515 add_14 ( .s(s[13]), .a(a[13]), .b(n_13_net_), .ci(c[12]), .co(c[13])
         );
  add_514 add_15 ( .s(s[14]), .a(a[14]), .b(n_14_net_), .ci(c[13]), .co(c[14])
         );
  add_513 add_16 ( .s(s[15]), .a(a[15]), .b(n_15_net_), .ci(c[14]), .co(c[15])
         );
  add_512 add_17 ( .s(s[16]), .a(a[16]), .b(n_16_net_), .ci(c[15]), .co(c[16])
         );
  add_511 add_18 ( .s(s[17]), .a(a[17]), .b(n_17_net_), .ci(c[16]), .co(c[17])
         );
  add_510 add_19 ( .s(s[18]), .a(a[18]), .b(n_18_net_), .ci(c[17]), .co(c[18])
         );
  add_509 add_20 ( .s(s[19]), .a(a[19]), .b(n_19_net_), .ci(c[18]), .co(c[19])
         );
  add_508 add_21 ( .s(s[20]), .a(a[20]), .b(n_20_net_), .ci(c[19]), .co(c[20])
         );
  add_507 add_22 ( .s(s[21]), .a(a[21]), .b(n_21_net_), .ci(c[20]), .co(c[21])
         );
  add_506 add_23 ( .s(s[22]), .a(a[22]), .b(n_22_net_), .ci(c[21]), .co(c[22])
         );
  add_505 add_24 ( .s(s[23]), .a(a[23]), .b(n_23_net_), .ci(c[22]), .co(c[23])
         );
  DFFARX1 out_reg_10_ ( .D(s[10]), .CLK(clk), .RSTB(rst_n), .Q(out[10]) );
  DFFARX1 out_reg_9_ ( .D(s[9]), .CLK(clk), .RSTB(rst_n), .Q(out[9]) );
  DFFARX1 out_reg_8_ ( .D(s[8]), .CLK(clk), .RSTB(rst_n), .Q(out[8]) );
  DFFARX1 out_reg_7_ ( .D(s[7]), .CLK(clk), .RSTB(rst_n), .Q(out[7]) );
  DFFARX1 out_reg_6_ ( .D(s[6]), .CLK(clk), .RSTB(rst_n), .Q(out[6]) );
  DFFARX1 out_reg_5_ ( .D(s[5]), .CLK(clk), .RSTB(rst_n), .Q(out[5]) );
  DFFARX1 out_reg_4_ ( .D(s[4]), .CLK(clk), .RSTB(rst_n), .Q(out[4]) );
  DFFARX1 out_reg_3_ ( .D(s[3]), .CLK(clk), .RSTB(rst_n), .Q(out[3]) );
  DFFARX1 out_reg_2_ ( .D(s[2]), .CLK(clk), .RSTB(rst_n), .Q(out[2]) );
  DFFARX1 out_reg_1_ ( .D(s[1]), .CLK(clk), .RSTB(rst_n), .Q(out[1]) );
  DFFARX1 out_reg_0_ ( .D(s[0]), .CLK(clk), .RSTB(rst_n), .Q(out[0]) );
  DFFARX1 c_tmp_reg ( .D(c[10]), .CLK(clk), .RSTB(rst_n), .Q(c_tmp) );
  DFFARX1 out_reg_24_ ( .D(s[24]), .CLK(clk), .RSTB(rst_n), .Q(out[24]) );
  DFFARX1 out_reg_23_ ( .D(s[23]), .CLK(clk), .RSTB(rst_n), .Q(out[23]) );
  DFFARX1 out_reg_22_ ( .D(s[22]), .CLK(clk), .RSTB(rst_n), .Q(out[22]) );
  DFFARX1 out_reg_21_ ( .D(s[21]), .CLK(clk), .RSTB(rst_n), .Q(out[21]) );
  DFFARX1 out_reg_20_ ( .D(s[20]), .CLK(clk), .RSTB(rst_n), .Q(out[20]) );
  DFFARX1 out_reg_19_ ( .D(s[19]), .CLK(clk), .RSTB(rst_n), .Q(out[19]) );
  DFFARX1 out_reg_18_ ( .D(s[18]), .CLK(clk), .RSTB(rst_n), .Q(out[18]) );
  DFFARX1 out_reg_17_ ( .D(s[17]), .CLK(clk), .RSTB(rst_n), .Q(out[17]) );
  DFFARX1 out_reg_16_ ( .D(s[16]), .CLK(clk), .RSTB(rst_n), .Q(out[16]) );
  DFFARX1 out_reg_15_ ( .D(s[15]), .CLK(clk), .RSTB(rst_n), .Q(out[15]) );
  DFFARX1 out_reg_14_ ( .D(s[14]), .CLK(clk), .RSTB(rst_n), .Q(out[14]) );
  DFFARX1 out_reg_13_ ( .D(s[13]), .CLK(clk), .RSTB(rst_n), .Q(out[13]) );
  DFFARX1 out_reg_12_ ( .D(s[12]), .CLK(clk), .RSTB(rst_n), .Q(out[12]) );
  DFFARX1 out_reg_11_ ( .D(s[11]), .CLK(clk), .RSTB(rst_n), .Q(out[11]) );
  INVX0 U3 ( .INP(b[1]), .ZN(n_1_net_) );
  INVX0 U4 ( .INP(b[2]), .ZN(n_2_net_) );
  INVX0 U5 ( .INP(b[3]), .ZN(n_3_net_) );
  INVX0 U6 ( .INP(b[4]), .ZN(n_4_net_) );
  INVX0 U7 ( .INP(b[5]), .ZN(n_5_net_) );
  INVX0 U8 ( .INP(b[6]), .ZN(n_6_net_) );
  INVX0 U9 ( .INP(b[7]), .ZN(n_7_net_) );
  INVX0 U10 ( .INP(b[8]), .ZN(n_8_net_) );
  INVX0 U11 ( .INP(b[9]), .ZN(n_9_net_) );
  INVX0 U12 ( .INP(b[10]), .ZN(n_10_net_) );
  INVX0 U13 ( .INP(c[23]), .ZN(s[24]) );
  INVX0 U14 ( .INP(b[11]), .ZN(n_11_net_) );
  INVX0 U15 ( .INP(b[12]), .ZN(n_12_net_) );
  INVX0 U16 ( .INP(b[13]), .ZN(n_13_net_) );
  INVX0 U17 ( .INP(b[14]), .ZN(n_14_net_) );
  INVX0 U18 ( .INP(b[15]), .ZN(n_15_net_) );
  INVX0 U19 ( .INP(b[16]), .ZN(n_16_net_) );
  INVX0 U20 ( .INP(b[17]), .ZN(n_17_net_) );
  INVX0 U21 ( .INP(b[18]), .ZN(n_18_net_) );
  INVX0 U22 ( .INP(b[19]), .ZN(n_19_net_) );
  INVX0 U23 ( .INP(b[20]), .ZN(n_20_net_) );
  INVX0 U24 ( .INP(b[21]), .ZN(n_21_net_) );
  INVX0 U25 ( .INP(b[22]), .ZN(n_22_net_) );
  INVX0 U26 ( .INP(b[23]), .ZN(n_23_net_) );
endmodule


module add_449 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  XNOR2X1 U1 ( .IN1(ci), .IN2(a), .Q(s) );
endmodule


module add_450 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_451 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_452 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_453 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_454 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_455 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_456 ( s, a, ci, co, b_BAR );
  input a, ci, b_BAR;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(b_BAR), .IN2(n1), .QN(co) );
  INVX0 U2 ( .INP(a), .ZN(n1) );
  MUX21X1 U3 ( .IN1(a), .IN2(n1), .S(b_BAR), .Q(s) );
endmodule


module adder8_33 ( out, a, b, cin );
  output [7:0] out;
  input [7:0] a;
  input [7:0] b;
  input cin;
  wire   n_1_net_, n_2_net_, n_4_net_;
  wire   [6:0] c;

  add_456 add_01 ( .s(out[0]), .a(a[0]), .ci(1'b1), .co(c[0]), .b_BAR(b[0]) );
  add_455 add_02 ( .s(out[1]), .a(a[1]), .b(n_1_net_), .ci(c[0]), .co(c[1]) );
  add_454 add_03 ( .s(out[2]), .a(a[2]), .b(n_2_net_), .ci(c[1]), .co(c[2]) );
  add_453 add_04 ( .s(out[3]), .a(a[3]), .b(1'b1), .ci(c[2]), .co(c[3]) );
  add_452 add_05 ( .s(out[4]), .a(a[4]), .b(n_4_net_), .ci(c[3]), .co(c[4]) );
  add_451 add_06 ( .s(out[5]), .a(a[5]), .b(1'b1), .ci(c[4]), .co(c[5]) );
  add_450 add_07 ( .s(out[6]), .a(a[6]), .b(1'b1), .ci(c[5]), .co(c[6]) );
  add_449 add_08 ( .s(out[7]), .a(a[7]), .b(1'b1), .ci(c[6]) );
  INVX0 U1 ( .INP(b[1]), .ZN(n_1_net_) );
  INVX0 U2 ( .INP(b[2]), .ZN(n_2_net_) );
  INVX0 U3 ( .INP(b[4]), .ZN(n_4_net_) );
endmodule


module add_457 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  XNOR2X1 U1 ( .IN1(ci), .IN2(a), .Q(s) );
endmodule


module add_458 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_459 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_460 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_461 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_462 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_463 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_464 ( s, a, ci, co, b_BAR );
  input a, ci, b_BAR;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(b_BAR), .IN2(n1), .QN(co) );
  INVX0 U2 ( .INP(a), .ZN(n1) );
  MUX21X1 U3 ( .IN1(a), .IN2(n1), .S(b_BAR), .Q(s) );
endmodule


module adder8_34 ( out, a, b, cin );
  output [7:0] out;
  input [7:0] a;
  input [7:0] b;
  input cin;
  wire   n_1_net_, n_2_net_, n_3_net_;
  wire   [6:0] c;

  add_464 add_01 ( .s(out[0]), .a(a[0]), .ci(1'b1), .co(c[0]), .b_BAR(b[0]) );
  add_463 add_02 ( .s(out[1]), .a(a[1]), .b(n_1_net_), .ci(c[0]), .co(c[1]) );
  add_462 add_03 ( .s(out[2]), .a(a[2]), .b(n_2_net_), .ci(c[1]), .co(c[2]) );
  add_461 add_04 ( .s(out[3]), .a(a[3]), .b(n_3_net_), .ci(c[2]), .co(c[3]) );
  add_460 add_05 ( .s(out[4]), .a(a[4]), .b(1'b1), .ci(c[3]), .co(c[4]) );
  add_459 add_06 ( .s(out[5]), .a(a[5]), .b(1'b1), .ci(c[4]), .co(c[5]) );
  add_458 add_07 ( .s(out[6]), .a(a[6]), .b(1'b1), .ci(c[5]), .co(c[6]) );
  add_457 add_08 ( .s(out[7]), .a(a[7]), .b(1'b1), .ci(c[6]) );
  INVX0 U1 ( .INP(b[1]), .ZN(n_1_net_) );
  INVX0 U2 ( .INP(b[2]), .ZN(n_2_net_) );
  INVX0 U3 ( .INP(b[3]), .ZN(n_3_net_) );
endmodule


module add_465 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  XNOR2X1 U1 ( .IN1(ci), .IN2(a), .Q(s) );
endmodule


module add_466 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_467 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_468 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_469 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_470 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_471 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_472 ( s, a, ci, co, b_BAR );
  input a, ci, b_BAR;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(b_BAR), .IN2(n1), .QN(co) );
  INVX0 U2 ( .INP(a), .ZN(n1) );
  MUX21X1 U3 ( .IN1(a), .IN2(n1), .S(b_BAR), .Q(s) );
endmodule


module adder8_35 ( out, a, b, cin );
  output [7:0] out;
  input [7:0] a;
  input [7:0] b;
  input cin;
  wire   n_1_net_, n_2_net_, n_3_net_;
  wire   [6:0] c;

  add_472 add_01 ( .s(out[0]), .a(a[0]), .ci(1'b1), .co(c[0]), .b_BAR(b[0]) );
  add_471 add_02 ( .s(out[1]), .a(a[1]), .b(n_1_net_), .ci(c[0]), .co(c[1]) );
  add_470 add_03 ( .s(out[2]), .a(a[2]), .b(n_2_net_), .ci(c[1]), .co(c[2]) );
  add_469 add_04 ( .s(out[3]), .a(a[3]), .b(n_3_net_), .ci(c[2]), .co(c[3]) );
  add_468 add_05 ( .s(out[4]), .a(a[4]), .b(1'b1), .ci(c[3]), .co(c[4]) );
  add_467 add_06 ( .s(out[5]), .a(a[5]), .b(1'b1), .ci(c[4]), .co(c[5]) );
  add_466 add_07 ( .s(out[6]), .a(a[6]), .b(1'b1), .ci(c[5]), .co(c[6]) );
  add_465 add_08 ( .s(out[7]), .a(a[7]), .b(1'b1), .ci(c[6]) );
  INVX0 U1 ( .INP(b[1]), .ZN(n_1_net_) );
  INVX0 U2 ( .INP(b[2]), .ZN(n_2_net_) );
  INVX0 U3 ( .INP(b[3]), .ZN(n_3_net_) );
endmodule


module add_473 ( s, a, b, co, ci_BAR );
  input a, b, ci_BAR;
  output s, co;


  XNOR2X1 U1 ( .IN1(a), .IN2(ci_BAR), .Q(s) );
endmodule


module add_474 ( s, a, b, ci, co_BAR );
  input a, b, ci;
  output s, co_BAR;


  NAND2X0 U1 ( .IN1(ci), .IN2(a), .QN(co_BAR) );
  OA21X1 U2 ( .IN1(ci), .IN2(a), .IN3(co_BAR), .Q(s) );
endmodule


module add_475 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_476 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_477 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_478 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_479 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_480 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(b), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(b), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module adder8_36 ( out, a, b, cin );
  output [7:0] out;
  input [7:0] a;
  input [7:0] b;
  input cin;

  wire   [6:0] c;

  add_480 add_01 ( .s(out[0]), .a(a[0]), .b(b[0]), .ci(1'b0), .co(c[0]) );
  add_479 add_02 ( .s(out[1]), .a(a[1]), .b(1'b0), .ci(c[0]), .co(c[1]) );
  add_478 add_03 ( .s(out[2]), .a(a[2]), .b(1'b0), .ci(c[1]), .co(c[2]) );
  add_477 add_04 ( .s(out[3]), .a(a[3]), .b(1'b0), .ci(c[2]), .co(c[3]) );
  add_476 add_05 ( .s(out[4]), .a(a[4]), .b(1'b0), .ci(c[3]), .co(c[4]) );
  add_475 add_06 ( .s(out[5]), .a(a[5]), .b(1'b0), .ci(c[4]), .co(c[5]) );
  add_474 add_07 ( .s(out[6]), .a(a[6]), .b(1'b0), .ci(c[5]), .co_BAR(c[6]) );
  add_473 add_08 ( .s(out[7]), .a(a[7]), .b(1'b0), .ci_BAR(c[6]) );
endmodule


module add_529 ( s, a, ci, co, b_BAR );
  input a, ci, b_BAR;
  output s, co;


  XNOR2X1 U1 ( .IN1(ci), .IN2(a), .Q(s) );
endmodule


module add_530 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_531 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_532 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_533 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_534 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_535 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_536 ( s, a, ci, co, b_BAR );
  input a, ci, b_BAR;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(b_BAR), .IN2(n1), .QN(co) );
  INVX0 U2 ( .INP(a), .ZN(n1) );
  MUX21X1 U3 ( .IN1(a), .IN2(n1), .S(b_BAR), .Q(s) );
endmodule


module adder8_37 ( out, a, b, cin );
  output [7:0] out;
  input [7:0] a;
  input [7:0] b;
  input cin;
  wire   n_1_net_, n_2_net_, n_3_net_, n_4_net_, n_5_net_, n_6_net_;
  wire   [6:0] c;

  add_536 add_01 ( .s(out[0]), .a(a[0]), .ci(1'b1), .co(c[0]), .b_BAR(b[0]) );
  add_535 add_02 ( .s(out[1]), .a(a[1]), .b(n_1_net_), .ci(c[0]), .co(c[1]) );
  add_534 add_03 ( .s(out[2]), .a(a[2]), .b(n_2_net_), .ci(c[1]), .co(c[2]) );
  add_533 add_04 ( .s(out[3]), .a(a[3]), .b(n_3_net_), .ci(c[2]), .co(c[3]) );
  add_532 add_05 ( .s(out[4]), .a(a[4]), .b(n_4_net_), .ci(c[3]), .co(c[4]) );
  add_531 add_06 ( .s(out[5]), .a(a[5]), .b(n_5_net_), .ci(c[4]), .co(c[5]) );
  add_530 add_07 ( .s(out[6]), .a(a[6]), .b(n_6_net_), .ci(c[5]), .co(c[6]) );
  add_529 add_08 ( .s(out[7]), .a(a[7]), .ci(c[6]), .b_BAR(1'b0) );
  INVX0 U1 ( .INP(b[1]), .ZN(n_1_net_) );
  INVX0 U2 ( .INP(b[2]), .ZN(n_2_net_) );
  INVX0 U3 ( .INP(b[3]), .ZN(n_3_net_) );
  INVX0 U4 ( .INP(b[4]), .ZN(n_4_net_) );
  INVX0 U5 ( .INP(b[5]), .ZN(n_5_net_) );
  INVX0 U6 ( .INP(b[6]), .ZN(n_6_net_) );
endmodule


module add_537 ( s, a, ci, co, b_BAR );
  input a, ci, b_BAR;
  output s, co;


  XNOR2X1 U1 ( .IN1(b_BAR), .IN2(ci), .Q(s) );
endmodule


module add_538 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_539 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_540 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_541 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_542 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_543 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_544 ( s, a, ci, co, b_BAR );
  input a, ci, b_BAR;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(b_BAR), .IN2(n1), .QN(co) );
  INVX0 U2 ( .INP(a), .ZN(n1) );
  MUX21X1 U3 ( .IN1(a), .IN2(n1), .S(b_BAR), .Q(s) );
endmodule


module adder8_38 ( out, a, b, cin );
  output [7:0] out;
  input [7:0] a;
  input [7:0] b;
  input cin;
  wire   n_1_net_, n_2_net_, n_3_net_, n_4_net_, n_5_net_, n_6_net_;
  wire   [6:0] c;

  add_544 add_01 ( .s(out[0]), .a(a[0]), .ci(1'b1), .co(c[0]), .b_BAR(b[0]) );
  add_543 add_02 ( .s(out[1]), .a(a[1]), .b(n_1_net_), .ci(c[0]), .co(c[1]) );
  add_542 add_03 ( .s(out[2]), .a(a[2]), .b(n_2_net_), .ci(c[1]), .co(c[2]) );
  add_541 add_04 ( .s(out[3]), .a(a[3]), .b(n_3_net_), .ci(c[2]), .co(c[3]) );
  add_540 add_05 ( .s(out[4]), .a(a[4]), .b(n_4_net_), .ci(c[3]), .co(c[4]) );
  add_539 add_06 ( .s(out[5]), .a(a[5]), .b(n_5_net_), .ci(c[4]), .co(c[5]) );
  add_538 add_07 ( .s(out[6]), .a(a[6]), .b(n_6_net_), .ci(c[5]), .co(c[6]) );
  add_537 add_08 ( .s(out[7]), .a(1'b0), .ci(c[6]), .b_BAR(b[7]) );
  INVX0 U1 ( .INP(b[1]), .ZN(n_1_net_) );
  INVX0 U2 ( .INP(b[2]), .ZN(n_2_net_) );
  INVX0 U3 ( .INP(b[3]), .ZN(n_3_net_) );
  INVX0 U4 ( .INP(b[4]), .ZN(n_4_net_) );
  INVX0 U5 ( .INP(b[5]), .ZN(n_5_net_) );
  INVX0 U6 ( .INP(b[6]), .ZN(n_6_net_) );
endmodule


module floating_point_adder_5 ( clk, rst_n, input_factor_01, input_factor_02, 
        output_adder );
  input [31:0] input_factor_01;
  input [31:0] input_factor_02;
  output [31:0] output_adder;
  input clk, rst_n;
  wire   N34, N35, N36, N37, N38, N39, N40, N41, N152, N153, N154, N155, N156,
         N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, N167,
         N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178,
         N179, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189,
         N190, N191, N192, N193, N194, N195, N196, N197, N198,
         add_sub_result_24_, N211, shift_temp_01_0_, N226, N227, N228, N229,
         N230, N231, N232, N233, N234, N235, N236, N237, N238, N239, N240,
         N241, N242, N243, N244, N245, N246, N247, N248, N256, N257, N258,
         N260, N261, N262, N263, N264, N265, N266, N267, N268, N269, N270,
         N271, N272, N273, N274, N275, N276, N277, N278, N279, N280, N281,
         N306, N307, N308, N346, N347, N348, N349, N350, N351, N352, N353,
         N354, N355, N380, N381, N382, N383, N384, N385, N386, N387, N388,
         N389, N390, N391, N392, N393, N394, N395, N396, N397, N398, N399,
         N400, N401, N402, N403, N404, N405, N406, N407, N408, N409, N410, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844;
  wire   [7:0] exp_diff_value;
  wire   [7:0] exponent_factor_21;
  wire   [7:0] exponent_factor_12;
  wire   [23:0] shift_smaller_factor;
  wire   [22:0] larger_factor;
  wire   [7:0] larger_exponent;
  wire   [24:0] add_result;
  wire   [24:0] sub_result;
  wire   [22:0] pre_sig_res_01;
  wire   [3:0] shift_temp_02;
  wire   [22:1] pre_sig_res_02;
  wire   [2:0] shift_temp_03;
  wire   [22:9] pre_sig_res_03;
  wire   [4:0] shift_temp_04;
  wire   [22:16] pre_sig_res_04;
  wire   [7:0] add_output_exponent_w1;
  wire   [7:0] add_output_exponent_w2;
  wire   [7:0] add_output_exponent_w3;
  wire   [7:0] add_output_exponent_w4;

  adder8_38 adder8_01 ( .out(exponent_factor_21), .a({1'b0, 
        input_factor_02[29:23]}), .b(input_factor_01[30:23]), .cin(1'b1) );
  adder8_37 adder8_02 ( .out(exponent_factor_12), .a(input_factor_01[30:23]), 
        .b({1'b0, input_factor_02[29:23]}), .cin(1'b1) );
  adder24_10 adder24_01 ( .clk(clk), .rst_n(rst_n), .a({shift_temp_04[4], 
        larger_factor}), .b(shift_smaller_factor), .cin(1'b1), .out(sub_result) );
  adder24_9 adder24_02 ( .clk(clk), .rst_n(rst_n), .a({shift_temp_04[4], 
        larger_factor}), .b(shift_smaller_factor), .cin(1'b0), .out(add_result) );
  adder8_36 adder8_03 ( .out(add_output_exponent_w1), .a(larger_exponent), .b(
        {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, shift_temp_01_0_}), .cin(
        1'b0) );
  adder8_35 adder8_04 ( .out(add_output_exponent_w2), .a(larger_exponent), .b(
        {1'b0, 1'b0, 1'b0, 1'b0, shift_temp_02}), .cin(1'b1) );
  adder8_34 adder8_05 ( .out(add_output_exponent_w3), .a(larger_exponent), .b(
        {1'b0, 1'b0, 1'b0, 1'b0, shift_temp_04[4], shift_temp_03}), .cin(1'b1)
         );
  adder8_33 adder8_06 ( .out(add_output_exponent_w4), .a(larger_exponent), .b(
        {1'b0, 1'b0, 1'b0, shift_temp_04[4], 1'b0, shift_temp_04[2:0]}), .cin(
        1'b1) );
  DFFARX1 exp_diff_value_reg_7_ ( .D(N41), .CLK(clk), .RSTB(rst_n), .Q(
        exp_diff_value[7]) );
  DFFARX1 exp_diff_value_reg_6_ ( .D(N40), .CLK(clk), .RSTB(rst_n), .Q(
        exp_diff_value[6]) );
  DFFARX1 exp_diff_value_reg_5_ ( .D(N39), .CLK(clk), .RSTB(rst_n), .Q(
        exp_diff_value[5]) );
  DFFARX1 exp_diff_value_reg_4_ ( .D(N38), .CLK(clk), .RSTB(rst_n), .Q(
        exp_diff_value[4]) );
  DFFARX1 exp_diff_value_reg_3_ ( .D(N37), .CLK(clk), .RSTB(rst_n), .Q(
        exp_diff_value[3]), .QN(n4) );
  DFFARX1 exp_diff_value_reg_2_ ( .D(N36), .CLK(clk), .RSTB(rst_n), .Q(
        exp_diff_value[2]), .QN(n1) );
  DFFARX1 exp_diff_value_reg_1_ ( .D(N35), .CLK(clk), .RSTB(rst_n), .Q(
        exp_diff_value[1]), .QN(n2) );
  DFFARX1 exp_diff_value_reg_0_ ( .D(N34), .CLK(clk), .RSTB(rst_n), .Q(
        exp_diff_value[0]), .QN(n3) );
  DFFARX1 larger_factor_reg_22_ ( .D(N198), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[22]) );
  DFFARX1 larger_factor_reg_21_ ( .D(N197), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[21]) );
  DFFARX1 larger_factor_reg_20_ ( .D(N196), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[20]) );
  DFFARX1 larger_factor_reg_19_ ( .D(N195), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[19]) );
  DFFARX1 larger_factor_reg_18_ ( .D(N194), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[18]) );
  DFFARX1 larger_factor_reg_17_ ( .D(N193), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[17]) );
  DFFARX1 larger_factor_reg_16_ ( .D(N192), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[16]) );
  DFFARX1 larger_factor_reg_15_ ( .D(N191), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[15]) );
  DFFARX1 larger_factor_reg_14_ ( .D(N190), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[14]) );
  DFFARX1 larger_factor_reg_13_ ( .D(N189), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[13]) );
  DFFARX1 larger_factor_reg_12_ ( .D(N188), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[12]) );
  DFFARX1 larger_factor_reg_11_ ( .D(N187), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[11]) );
  DFFARX1 larger_factor_reg_10_ ( .D(N186), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[10]) );
  DFFARX1 larger_factor_reg_9_ ( .D(N185), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[9]) );
  DFFARX1 larger_factor_reg_8_ ( .D(N184), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[8]) );
  DFFARX1 larger_factor_reg_7_ ( .D(N183), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[7]) );
  DFFARX1 larger_factor_reg_6_ ( .D(N182), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[6]) );
  DFFARX1 larger_factor_reg_5_ ( .D(N181), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[5]) );
  DFFARX1 larger_factor_reg_4_ ( .D(N180), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[4]) );
  DFFARX1 larger_factor_reg_3_ ( .D(N179), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[3]) );
  DFFARX1 larger_factor_reg_2_ ( .D(N178), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[2]) );
  DFFARX1 larger_factor_reg_1_ ( .D(N177), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[1]) );
  DFFARX1 larger_factor_reg_0_ ( .D(N176), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[0]) );
  DFFARX1 shift_smaller_factor_reg_23_ ( .D(N175), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[23]) );
  DFFARX1 shift_smaller_factor_reg_22_ ( .D(N174), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[22]) );
  DFFARX1 shift_smaller_factor_reg_21_ ( .D(N173), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[21]) );
  DFFARX1 shift_smaller_factor_reg_20_ ( .D(N172), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[20]) );
  DFFARX1 shift_smaller_factor_reg_19_ ( .D(N171), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[19]) );
  DFFARX1 shift_smaller_factor_reg_18_ ( .D(N170), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[18]) );
  DFFARX1 shift_smaller_factor_reg_17_ ( .D(N169), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[17]) );
  DFFARX1 shift_smaller_factor_reg_16_ ( .D(N168), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[16]) );
  DFFARX1 shift_smaller_factor_reg_15_ ( .D(N167), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[15]) );
  DFFARX1 shift_smaller_factor_reg_14_ ( .D(N166), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[14]) );
  DFFARX1 shift_smaller_factor_reg_13_ ( .D(N165), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[13]) );
  DFFARX1 shift_smaller_factor_reg_12_ ( .D(N164), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[12]) );
  DFFARX1 shift_smaller_factor_reg_11_ ( .D(N163), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[11]) );
  DFFARX1 shift_smaller_factor_reg_10_ ( .D(N162), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[10]) );
  DFFARX1 shift_smaller_factor_reg_9_ ( .D(N161), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[9]) );
  DFFARX1 shift_smaller_factor_reg_8_ ( .D(N160), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[8]) );
  DFFARX1 shift_smaller_factor_reg_7_ ( .D(N159), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[7]) );
  DFFARX1 shift_smaller_factor_reg_6_ ( .D(N158), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[6]) );
  DFFARX1 shift_smaller_factor_reg_5_ ( .D(N157), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[5]) );
  DFFARX1 shift_smaller_factor_reg_4_ ( .D(N156), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[4]) );
  DFFARX1 shift_smaller_factor_reg_3_ ( .D(N155), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[3]) );
  DFFARX1 shift_smaller_factor_reg_2_ ( .D(N154), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[2]) );
  DFFARX1 shift_smaller_factor_reg_1_ ( .D(N153), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[1]) );
  DFFARX1 shift_smaller_factor_reg_0_ ( .D(N152), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[0]) );
  DFFX1 larger_exponent_reg_7_ ( .D(n822), .CLK(clk), .Q(larger_exponent[7])
         );
  DFFX1 larger_exponent_reg_6_ ( .D(n823), .CLK(clk), .Q(larger_exponent[6])
         );
  DFFX1 larger_exponent_reg_5_ ( .D(n824), .CLK(clk), .Q(larger_exponent[5])
         );
  DFFX1 larger_exponent_reg_4_ ( .D(n825), .CLK(clk), .Q(larger_exponent[4])
         );
  DFFX1 larger_exponent_reg_3_ ( .D(n826), .CLK(clk), .Q(larger_exponent[3])
         );
  DFFX1 larger_exponent_reg_2_ ( .D(n827), .CLK(clk), .Q(larger_exponent[2])
         );
  DFFX1 larger_exponent_reg_1_ ( .D(n828), .CLK(clk), .Q(larger_exponent[1])
         );
  DFFX1 larger_exponent_reg_0_ ( .D(n829), .CLK(clk), .Q(larger_exponent[0])
         );
  DFFARX1 shift_temp_04_reg_4_ ( .D(1'b1), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_04[4]) );
  DFFARX1 shift_temp_01_reg_0_ ( .D(add_sub_result_24_), .CLK(clk), .RSTB(
        rst_n), .Q(shift_temp_01_0_) );
  DFFARX1 pre_sig_res_02_reg_1_ ( .D(N260), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[1]) );
  DFFARX1 pre_sig_res_02_reg_2_ ( .D(N261), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[2]) );
  DFFARX1 pre_sig_res_02_reg_3_ ( .D(N262), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[3]) );
  DFFARX1 pre_sig_res_02_reg_4_ ( .D(N263), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[4]) );
  DFFARX1 pre_sig_res_02_reg_5_ ( .D(N264), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[5]) );
  DFFARX1 pre_sig_res_02_reg_6_ ( .D(N265), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[6]) );
  DFFARX1 pre_sig_res_02_reg_7_ ( .D(N266), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[7]) );
  DFFARX1 shift_temp_02_reg_2_ ( .D(N258), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_02[2]) );
  DFFASX1 shift_temp_02_reg_3_ ( .D(n821), .CLK(clk), .SETB(rst_n), .QN(
        shift_temp_02[3]) );
  DFFARX1 pre_sig_res_02_reg_8_ ( .D(N267), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[8]) );
  DFFARX1 pre_sig_res_02_reg_9_ ( .D(N268), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[9]) );
  DFFARX1 pre_sig_res_02_reg_10_ ( .D(N269), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[10]) );
  DFFARX1 pre_sig_res_02_reg_11_ ( .D(N270), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[11]) );
  DFFARX1 pre_sig_res_02_reg_12_ ( .D(N271), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[12]) );
  DFFARX1 pre_sig_res_02_reg_13_ ( .D(N272), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[13]) );
  DFFARX1 pre_sig_res_02_reg_14_ ( .D(N273), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[14]) );
  DFFARX1 pre_sig_res_02_reg_15_ ( .D(N274), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[15]) );
  DFFARX1 pre_sig_res_02_reg_16_ ( .D(N275), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[16]) );
  DFFARX1 pre_sig_res_02_reg_17_ ( .D(N276), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[17]) );
  DFFARX1 pre_sig_res_02_reg_18_ ( .D(N277), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[18]) );
  DFFARX1 pre_sig_res_02_reg_19_ ( .D(N278), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[19]) );
  DFFARX1 pre_sig_res_02_reg_20_ ( .D(N279), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[20]) );
  DFFARX1 pre_sig_res_02_reg_21_ ( .D(N280), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[21]) );
  DFFARX1 pre_sig_res_02_reg_22_ ( .D(N281), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[22]) );
  DFFARX1 shift_temp_02_reg_1_ ( .D(N257), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_02[1]) );
  DFFARX1 shift_temp_02_reg_0_ ( .D(N256), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_02[0]) );
  DFFX1 pre_sig_res_03_reg_9_ ( .D(n830), .CLK(clk), .Q(pre_sig_res_03[9]) );
  DFFX1 pre_sig_res_03_reg_10_ ( .D(n831), .CLK(clk), .Q(pre_sig_res_03[10])
         );
  DFFX1 pre_sig_res_03_reg_12_ ( .D(n832), .CLK(clk), .Q(pre_sig_res_03[12])
         );
  DFFX1 pre_sig_res_03_reg_11_ ( .D(n833), .CLK(clk), .Q(pre_sig_res_03[11])
         );
  DFFX1 pre_sig_res_03_reg_13_ ( .D(n834), .CLK(clk), .Q(pre_sig_res_03[13])
         );
  DFFX1 pre_sig_res_03_reg_14_ ( .D(n835), .CLK(clk), .Q(pre_sig_res_03[14])
         );
  DFFARX1 shift_temp_03_reg_2_ ( .D(N308), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_03[2]) );
  DFFARX1 shift_temp_03_reg_0_ ( .D(N306), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_03[0]) );
  DFFARX1 shift_temp_03_reg_1_ ( .D(N307), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_03[1]) );
  DFFX1 pre_sig_res_03_reg_15_ ( .D(n836), .CLK(clk), .Q(pre_sig_res_03[15])
         );
  DFFX1 pre_sig_res_03_reg_16_ ( .D(n837), .CLK(clk), .Q(pre_sig_res_03[16])
         );
  DFFX1 pre_sig_res_03_reg_17_ ( .D(n838), .CLK(clk), .Q(pre_sig_res_03[17])
         );
  DFFX1 pre_sig_res_03_reg_18_ ( .D(n839), .CLK(clk), .Q(pre_sig_res_03[18])
         );
  DFFX1 pre_sig_res_03_reg_19_ ( .D(n840), .CLK(clk), .Q(pre_sig_res_03[19])
         );
  DFFX1 pre_sig_res_03_reg_20_ ( .D(n841), .CLK(clk), .Q(pre_sig_res_03[20])
         );
  DFFX1 pre_sig_res_03_reg_21_ ( .D(n842), .CLK(clk), .Q(pre_sig_res_03[21])
         );
  DFFX1 pre_sig_res_03_reg_22_ ( .D(n843), .CLK(clk), .Q(pre_sig_res_03[22])
         );
  DFFARX1 pre_sig_res_04_reg_16_ ( .D(N349), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_04[16]) );
  DFFARX1 pre_sig_res_04_reg_17_ ( .D(N350), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_04[17]) );
  DFFARX1 pre_sig_res_04_reg_18_ ( .D(N351), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_04[18]) );
  DFFARX1 pre_sig_res_04_reg_19_ ( .D(N352), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_04[19]) );
  DFFARX1 pre_sig_res_04_reg_20_ ( .D(N353), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_04[20]) );
  DFFARX1 pre_sig_res_04_reg_21_ ( .D(N354), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_04[21]) );
  DFFARX1 pre_sig_res_04_reg_22_ ( .D(N355), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_04[22]) );
  DFFARX1 add_output_sign_reg ( .D(N211), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[31]) );
  DFFARX1 pre_sig_res_01_reg_0_ ( .D(N226), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[0]) );
  DFFARX1 pre_sig_res_01_reg_1_ ( .D(N227), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[1]) );
  DFFARX1 pre_sig_res_01_reg_2_ ( .D(N228), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[2]) );
  DFFARX1 pre_sig_res_01_reg_3_ ( .D(N229), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[3]) );
  DFFARX1 pre_sig_res_01_reg_4_ ( .D(N230), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[4]) );
  DFFARX1 pre_sig_res_01_reg_5_ ( .D(N231), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[5]) );
  DFFARX1 pre_sig_res_01_reg_6_ ( .D(N232), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[6]) );
  DFFARX1 pre_sig_res_01_reg_7_ ( .D(N233), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[7]) );
  DFFARX1 pre_sig_res_01_reg_8_ ( .D(N234), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[8]) );
  DFFARX1 pre_sig_res_01_reg_9_ ( .D(N235), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[9]) );
  DFFARX1 pre_sig_res_01_reg_10_ ( .D(N236), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[10]) );
  DFFARX1 pre_sig_res_01_reg_11_ ( .D(N237), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[11]) );
  DFFARX1 pre_sig_res_01_reg_12_ ( .D(N238), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[12]) );
  DFFARX1 pre_sig_res_01_reg_13_ ( .D(N239), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[13]) );
  DFFARX1 pre_sig_res_01_reg_14_ ( .D(N240), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[14]) );
  DFFARX1 pre_sig_res_01_reg_15_ ( .D(N241), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[15]) );
  DFFARX1 pre_sig_res_01_reg_16_ ( .D(N242), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[16]) );
  DFFARX1 pre_sig_res_01_reg_17_ ( .D(N243), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[17]) );
  DFFARX1 pre_sig_res_01_reg_18_ ( .D(N244), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[18]) );
  DFFARX1 pre_sig_res_01_reg_19_ ( .D(N245), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[19]) );
  DFFARX1 pre_sig_res_01_reg_20_ ( .D(N246), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[20]) );
  DFFARX1 pre_sig_res_01_reg_21_ ( .D(N247), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[21]) );
  DFFARX1 pre_sig_res_01_reg_22_ ( .D(N248), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[22]) );
  DFFARX1 shift_temp_04_reg_2_ ( .D(N348), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_04[2]) );
  DFFARX1 shift_temp_04_reg_1_ ( .D(N347), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_04[1]) );
  DFFARX1 shift_temp_04_reg_0_ ( .D(N346), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_04[0]) );
  DFFARX1 add_output_exponent_reg_7_ ( .D(N387), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[30]) );
  DFFARX1 add_output_exponent_reg_6_ ( .D(N386), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[29]) );
  DFFARX1 add_output_exponent_reg_5_ ( .D(N385), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[28]) );
  DFFARX1 add_output_exponent_reg_4_ ( .D(N384), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[27]) );
  DFFARX1 add_output_exponent_reg_3_ ( .D(N383), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[26]) );
  DFFARX1 add_output_exponent_reg_2_ ( .D(N382), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[25]) );
  DFFARX1 add_output_exponent_reg_1_ ( .D(N381), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[24]) );
  DFFARX1 add_output_exponent_reg_0_ ( .D(N380), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[23]) );
  DFFARX1 add_output_significands_reg_22_ ( .D(N410), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[22]) );
  DFFARX1 add_output_significands_reg_21_ ( .D(N409), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[21]) );
  DFFARX1 add_output_significands_reg_20_ ( .D(N408), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[20]) );
  DFFARX1 add_output_significands_reg_19_ ( .D(N407), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[19]) );
  DFFARX1 add_output_significands_reg_18_ ( .D(N406), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[18]) );
  DFFARX1 add_output_significands_reg_17_ ( .D(N405), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[17]) );
  DFFARX1 add_output_significands_reg_16_ ( .D(N404), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[16]) );
  DFFARX1 add_output_significands_reg_15_ ( .D(N403), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[15]) );
  DFFARX1 add_output_significands_reg_14_ ( .D(N402), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[14]) );
  DFFARX1 add_output_significands_reg_13_ ( .D(N401), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[13]) );
  DFFARX1 add_output_significands_reg_12_ ( .D(N400), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[12]) );
  DFFARX1 add_output_significands_reg_11_ ( .D(N399), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[11]) );
  DFFARX1 add_output_significands_reg_10_ ( .D(N398), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[10]) );
  DFFARX1 add_output_significands_reg_9_ ( .D(N397), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[9]) );
  DFFARX1 add_output_significands_reg_8_ ( .D(N396), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[8]) );
  DFFARX1 add_output_significands_reg_7_ ( .D(N395), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[7]) );
  DFFARX1 add_output_significands_reg_6_ ( .D(N394), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[6]) );
  DFFARX1 add_output_significands_reg_5_ ( .D(N393), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[5]) );
  DFFARX1 add_output_significands_reg_4_ ( .D(N392), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[4]) );
  DFFARX1 add_output_significands_reg_3_ ( .D(N391), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[3]) );
  DFFARX1 add_output_significands_reg_2_ ( .D(N390), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[2]) );
  DFFARX1 add_output_significands_reg_1_ ( .D(N389), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[1]) );
  DFFARX1 add_output_significands_reg_0_ ( .D(N388), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[0]) );
  INVX1 U5 ( .INP(rst_n), .ZN(n844) );
  NAND2X0 U3 ( .IN1(input_factor_02[11]), .IN2(n638), .QN(n57) );
  NAND2X0 U4 ( .IN1(n482), .IN2(n395), .QN(n562) );
  NAND2X0 U6 ( .IN1(input_factor_02[16]), .IN2(n370), .QN(n70) );
  NAND2X0 U7 ( .IN1(input_factor_02[24]), .IN2(n541), .QN(n34) );
  NAND2X0 U8 ( .IN1(input_factor_01[27]), .IN2(n588), .QN(n30) );
  NAND2X0 U9 ( .IN1(input_factor_01[26]), .IN2(n582), .QN(n31) );
  NAND2X0 U10 ( .IN1(input_factor_01[28]), .IN2(n594), .QN(n41) );
  NAND2X0 U11 ( .IN1(input_factor_02[28]), .IN2(n593), .QN(n45) );
  NAND2X0 U12 ( .IN1(n801), .IN2(n522), .QN(n381) );
  NAND2X0 U13 ( .IN1(n771), .IN2(n514), .QN(n380) );
  NAND2X0 U14 ( .IN1(n764), .IN2(n515), .QN(n379) );
  NAND2X0 U15 ( .IN1(n740), .IN2(n714), .QN(n559) );
  NAND2X0 U16 ( .IN1(n399), .IN2(n492), .QN(n377) );
  NAND2X0 U17 ( .IN1(n490), .IN2(n402), .QN(n376) );
  NAND2X0 U18 ( .IN1(n375), .IN2(n568), .QN(n401) );
  NAND2X0 U19 ( .IN1(n91), .IN2(n90), .QN(n217) );
  NAND2X0 U20 ( .IN1(n166), .IN2(n165), .QN(n250) );
  NAND2X0 U21 ( .IN1(n200), .IN2(n199), .QN(n269) );
  NAND2X0 U22 ( .IN1(exp_diff_value[1]), .IN2(exp_diff_value[0]), .QN(n198) );
  NAND2X0 U23 ( .IN1(exp_diff_value[1]), .IN2(n3), .QN(n196) );
  NAND2X0 U24 ( .IN1(exp_diff_value[0]), .IN2(n2), .QN(n197) );
  NAND2X0 U25 ( .IN1(n353), .IN2(n217), .QN(n218) );
  NAND2X0 U26 ( .IN1(n698), .IN2(n268), .QN(n248) );
  NAND2X0 U27 ( .IN1(n164), .IN2(n163), .QN(n246) );
  NAND2X0 U28 ( .IN1(n353), .IN2(n250), .QN(n251) );
  NAND2X0 U29 ( .IN1(n268), .IN2(n817), .QN(n252) );
  NAND2X0 U30 ( .IN1(n195), .IN2(n194), .QN(n265) );
  NAND2X0 U31 ( .IN1(n353), .IN2(n269), .QN(n270) );
  NAND2X0 U32 ( .IN1(n126), .IN2(n125), .QN(n230) );
  NAND2X0 U33 ( .IN1(n70), .IN2(n71), .QN(n18) );
  NAND2X0 U34 ( .IN1(n693), .IN2(n2), .QN(n120) );
  NAND2X0 U35 ( .IN1(input_factor_02[19]), .IN2(n683), .QN(n65) );
  NAND2X0 U36 ( .IN1(n702), .IN2(n3), .QN(n147) );
  NAND2X0 U37 ( .IN1(input_factor_01[23]), .IN2(n557), .QN(n32) );
  NAND2X0 U38 ( .IN1(n542), .IN2(input_factor_02[25]), .QN(n33) );
  NAND2X0 U39 ( .IN1(input_factor_02[27]), .IN2(n587), .QN(n24) );
  NAND2X0 U40 ( .IN1(input_factor_02[26]), .IN2(n581), .QN(n22) );
  NAND2X0 U41 ( .IN1(n373), .IN2(n74), .QN(n176) );
  NAND2X0 U42 ( .IN1(n706), .IN2(pre_sig_res_01[9]), .QN(n630) );
  NAND2X0 U43 ( .IN1(n706), .IN2(pre_sig_res_01[10]), .QN(n636) );
  NAND2X0 U44 ( .IN1(n706), .IN2(pre_sig_res_01[11]), .QN(n642) );
  NAND2X0 U45 ( .IN1(n706), .IN2(pre_sig_res_01[13]), .QN(n651) );
  NAND2X0 U46 ( .IN1(n706), .IN2(pre_sig_res_01[14]), .QN(n657) );
  NAND2X0 U47 ( .IN1(n706), .IN2(pre_sig_res_01[15]), .QN(n663) );
  NAND2X0 U48 ( .IN1(n706), .IN2(pre_sig_res_01[16]), .QN(n667) );
  NAND2X0 U49 ( .IN1(n706), .IN2(pre_sig_res_01[17]), .QN(n673) );
  NAND2X0 U50 ( .IN1(n706), .IN2(pre_sig_res_01[18]), .QN(n679) );
  NAND2X0 U51 ( .IN1(n706), .IN2(pre_sig_res_01[19]), .QN(n685) );
  NAND2X0 U52 ( .IN1(n706), .IN2(pre_sig_res_01[21]), .QN(n694) );
  NAND2X0 U53 ( .IN1(n706), .IN2(pre_sig_res_01[22]), .QN(n707) );
  NAND2X0 U54 ( .IN1(n706), .IN2(add_output_exponent_w1[0]), .QN(n569) );
  NAND2X0 U55 ( .IN1(n706), .IN2(add_output_exponent_w1[1]), .QN(n573) );
  NAND2X0 U56 ( .IN1(n706), .IN2(add_output_exponent_w1[2]), .QN(n577) );
  NAND2X0 U57 ( .IN1(n706), .IN2(add_output_exponent_w1[3]), .QN(n583) );
  NAND2X0 U58 ( .IN1(n706), .IN2(add_output_exponent_w1[4]), .QN(n589) );
  NAND2X0 U59 ( .IN1(n706), .IN2(add_output_exponent_w1[5]), .QN(n595) );
  NAND2X0 U60 ( .IN1(n706), .IN2(add_output_exponent_w1[6]), .QN(n601) );
  NAND2X0 U61 ( .IN1(n516), .IN2(n811), .QN(n534) );
  NAND2X0 U62 ( .IN1(n513), .IN2(n522), .QN(n519) );
  NAND2X0 U63 ( .IN1(n176), .IN2(n360), .QN(n391) );
  NAND2X0 U64 ( .IN1(n514), .IN2(n784), .QN(n532) );
  NAND2X0 U65 ( .IN1(n515), .IN2(n751), .QN(n533) );
  NAND2X0 U66 ( .IN1(n756), .IN2(n740), .QN(n715) );
  NAND2X0 U67 ( .IN1(n714), .IN2(n727), .QN(n789) );
  NAND2X0 U68 ( .IN1(n512), .IN2(n500), .QN(n718) );
  NAND2X0 U69 ( .IN1(n512), .IN2(n504), .QN(n711) );
  NAND2X0 U70 ( .IN1(n395), .IN2(n394), .QN(n494) );
  NAND2X0 U71 ( .IN1(n412), .IN2(n813), .QN(n409) );
  NAND2X0 U72 ( .IN1(n399), .IN2(n396), .QN(n483) );
  NAND2X0 U73 ( .IN1(n402), .IN2(n397), .QN(n487) );
  NAND2X0 U74 ( .IN1(n398), .IN2(n568), .QN(n485) );
  NAND2X0 U75 ( .IN1(n162), .IN2(n161), .QN(n167) );
  NAND2X0 U76 ( .IN1(n268), .IN2(n4), .QN(n177) );
  NAND2X0 U77 ( .IN1(n817), .IN2(n372), .QN(n271) );
  NAND2X0 U78 ( .IN1(n698), .IN2(n372), .QN(n232) );
  NAND2X0 U79 ( .IN1(n191), .IN2(n190), .QN(n201) );
  NAND2X0 U80 ( .IN1(n89), .IN2(n88), .QN(n215) );
  NAND2X0 U81 ( .IN1(n218), .IN2(n219), .QN(n16) );
  NAND2X0 U82 ( .IN1(n4), .IN2(n1), .QN(n275) );
  NAND2X0 U83 ( .IN1(n251), .IN2(n253), .QN(n14) );
  NAND2X0 U84 ( .IN1(n354), .IN2(n207), .QN(n262) );
  NAND2X0 U85 ( .IN1(n270), .IN2(n273), .QN(n12) );
  NAND2X0 U86 ( .IN1(exp_diff_value[3]), .IN2(n354), .QN(n330) );
  NAND2X0 U87 ( .IN1(n307), .IN2(n1), .QN(n322) );
  NAND2X0 U88 ( .IN1(n330), .IN2(n329), .QN(n331) );
  NAND2X0 U89 ( .IN1(n353), .IN2(n4), .QN(n347) );
  NAND2X0 U90 ( .IN1(n354), .IN2(n4), .QN(n349) );
  NAND2X0 U91 ( .IN1(n363), .IN2(n69), .QN(n360) );
  NAND2X0 U92 ( .IN1(n2), .IN2(n147), .QN(n367) );
  NAND2X0 U93 ( .IN1(n371), .IN2(n353), .QN(n366) );
  NAND2X0 U94 ( .IN1(n354), .IN2(n371), .QN(n364) );
  NAND2X0 U95 ( .IN1(n608), .IN2(n607), .QN(N390) );
  NAND2X0 U96 ( .IN1(n610), .IN2(n609), .QN(N391) );
  NAND2X0 U97 ( .IN1(n612), .IN2(n611), .QN(N392) );
  NAND2X0 U98 ( .IN1(n616), .IN2(n615), .QN(N393) );
  NAND2X0 U99 ( .IN1(n618), .IN2(n617), .QN(N394) );
  NAND2X0 U100 ( .IN1(n621), .IN2(n620), .QN(N395) );
  NAND2X0 U101 ( .IN1(n625), .IN2(n624), .QN(N396) );
  NAND2X0 U102 ( .IN1(n704), .IN2(pre_sig_res_03[9]), .QN(n628) );
  NAND2X0 U103 ( .IN1(n703), .IN2(pre_sig_res_02[9]), .QN(n629) );
  NAND2X0 U104 ( .IN1(n704), .IN2(pre_sig_res_03[10]), .QN(n634) );
  NAND2X0 U105 ( .IN1(n703), .IN2(pre_sig_res_02[10]), .QN(n635) );
  NAND2X0 U106 ( .IN1(n704), .IN2(pre_sig_res_03[11]), .QN(n640) );
  NAND2X0 U107 ( .IN1(n703), .IN2(pre_sig_res_02[11]), .QN(n641) );
  NAND2X0 U108 ( .IN1(n7), .IN2(n8), .QN(N400) );
  NAND2X0 U109 ( .IN1(pre_sig_res_01[12]), .IN2(n706), .QN(n8) );
  NAND2X0 U110 ( .IN1(n704), .IN2(pre_sig_res_03[13]), .QN(n649) );
  NAND2X0 U111 ( .IN1(n703), .IN2(pre_sig_res_02[13]), .QN(n650) );
  NAND2X0 U112 ( .IN1(n704), .IN2(pre_sig_res_03[14]), .QN(n655) );
  NAND2X0 U113 ( .IN1(n703), .IN2(pre_sig_res_02[14]), .QN(n656) );
  NAND2X0 U114 ( .IN1(n704), .IN2(pre_sig_res_03[15]), .QN(n661) );
  NAND2X0 U115 ( .IN1(n703), .IN2(pre_sig_res_02[15]), .QN(n662) );
  NAND2X0 U116 ( .IN1(n705), .IN2(pre_sig_res_04[16]), .QN(n668) );
  NAND2X0 U117 ( .IN1(n705), .IN2(pre_sig_res_04[17]), .QN(n674) );
  NAND2X0 U118 ( .IN1(n705), .IN2(pre_sig_res_04[18]), .QN(n680) );
  NAND2X0 U119 ( .IN1(n705), .IN2(pre_sig_res_04[19]), .QN(n686) );
  NAND2X0 U120 ( .IN1(n5), .IN2(n6), .QN(N408) );
  NAND2X0 U121 ( .IN1(n705), .IN2(pre_sig_res_04[20]), .QN(n6) );
  NAND2X0 U122 ( .IN1(n705), .IN2(pre_sig_res_04[21]), .QN(n695) );
  NAND2X0 U123 ( .IN1(n705), .IN2(pre_sig_res_04[22]), .QN(n708) );
  NAND2X0 U124 ( .IN1(n705), .IN2(add_output_exponent_w4[0]), .QN(n570) );
  NAND2X0 U125 ( .IN1(n705), .IN2(add_output_exponent_w4[1]), .QN(n574) );
  NAND2X0 U126 ( .IN1(n705), .IN2(add_output_exponent_w4[2]), .QN(n578) );
  NAND2X0 U127 ( .IN1(n705), .IN2(add_output_exponent_w4[3]), .QN(n584) );
  NAND2X0 U128 ( .IN1(n705), .IN2(add_output_exponent_w4[4]), .QN(n590) );
  NAND2X0 U129 ( .IN1(n705), .IN2(add_output_exponent_w4[5]), .QN(n596) );
  NAND2X0 U130 ( .IN1(n705), .IN2(add_output_exponent_w4[6]), .QN(n602) );
  NAND2X0 U131 ( .IN1(n9), .IN2(n10), .QN(N387) );
  NAND2X0 U132 ( .IN1(n705), .IN2(add_output_exponent_w4[7]), .QN(n10) );
  NAND2X0 U133 ( .IN1(n519), .IN2(n518), .QN(N348) );
  NAND2X0 U134 ( .IN1(n536), .IN2(n791), .QN(n537) );
  NAND2X0 U135 ( .IN1(n536), .IN2(n811), .QN(n527) );
  NAND2X0 U136 ( .IN1(n536), .IN2(n813), .QN(n523) );
  NAND2X0 U137 ( .IN1(n521), .IN2(n520), .QN(N352) );
  NAND2X0 U138 ( .IN1(pre_sig_res_03[22]), .IN2(n815), .QN(n720) );
  NAND2X0 U139 ( .IN1(n804), .IN2(n719), .QN(n721) );
  NAND2X0 U140 ( .IN1(pre_sig_res_03[21]), .IN2(n815), .QN(n728) );
  NAND2X0 U141 ( .IN1(n804), .IN2(n727), .QN(n729) );
  NAND2X0 U142 ( .IN1(pre_sig_res_03[20]), .IN2(n815), .QN(n736) );
  NAND2X0 U143 ( .IN1(n804), .IN2(n735), .QN(n737) );
  NAND2X0 U144 ( .IN1(pre_sig_res_03[19]), .IN2(n815), .QN(n744) );
  NAND2X0 U145 ( .IN1(n804), .IN2(n743), .QN(n745) );
  NAND2X0 U146 ( .IN1(pre_sig_res_03[18]), .IN2(n815), .QN(n752) );
  NAND2X0 U147 ( .IN1(n804), .IN2(n751), .QN(n753) );
  NAND2X0 U148 ( .IN1(pre_sig_res_03[17]), .IN2(n815), .QN(n760) );
  NAND2X0 U149 ( .IN1(n804), .IN2(n759), .QN(n761) );
  NAND2X0 U150 ( .IN1(pre_sig_res_03[16]), .IN2(n815), .QN(n767) );
  NAND2X0 U151 ( .IN1(n804), .IN2(n784), .QN(n768) );
  NAND2X0 U152 ( .IN1(pre_sig_res_03[15]), .IN2(n815), .QN(n776) );
  NAND2X0 U153 ( .IN1(n804), .IN2(n792), .QN(n777) );
  NAND2X0 U154 ( .IN1(n711), .IN2(n718), .QN(n505) );
  NAND2X0 U155 ( .IN1(pre_sig_res_03[14]), .IN2(n844), .QN(n786) );
  NAND2X0 U156 ( .IN1(n814), .IN2(n784), .QN(n785) );
  NAND2X0 U157 ( .IN1(n804), .IN2(n783), .QN(n787) );
  NAND2X0 U158 ( .IN1(pre_sig_res_03[13]), .IN2(n815), .QN(n794) );
  NAND2X0 U159 ( .IN1(n814), .IN2(n792), .QN(n793) );
  NAND2X0 U160 ( .IN1(n804), .IN2(n791), .QN(n795) );
  NAND2X0 U161 ( .IN1(n799), .IN2(n798), .QN(n833) );
  NAND2X0 U162 ( .IN1(pre_sig_res_03[12]), .IN2(n815), .QN(n807) );
  NAND2X0 U163 ( .IN1(n804), .IN2(n811), .QN(n809) );
  NAND2X0 U164 ( .IN1(n412), .IN2(n811), .QN(n413) );
  NAND2X0 U165 ( .IN1(n417), .IN2(n792), .QN(n408) );
  NAND2X0 U166 ( .IN1(n418), .IN2(n791), .QN(n405) );
  NAND2X0 U167 ( .IN1(n404), .IN2(n403), .QN(N263) );
  NAND2X0 U168 ( .IN1(n308), .IN2(input_factor_01[0]), .QN(n119) );
  NAND2X0 U169 ( .IN1(n146), .IN2(n145), .QN(N153) );
  NAND2X0 U170 ( .IN1(n308), .IN2(input_factor_01[2]), .QN(n172) );
  NAND2X0 U171 ( .IN1(n308), .IN2(input_factor_01[3]), .QN(n206) );
  NAND2X0 U172 ( .IN1(input_factor_01[4]), .IN2(n308), .QN(n222) );
  NAND2X0 U173 ( .IN1(input_factor_01[6]), .IN2(n308), .QN(n256) );
  NAND2X0 U174 ( .IN1(input_factor_01[7]), .IN2(n308), .QN(n277) );
  NAND2X0 U175 ( .IN1(input_factor_01[12]), .IN2(n308), .QN(n309) );
  NAND2X0 U176 ( .IN1(n338), .IN2(n337), .QN(N168) );
  NAND2X0 U177 ( .IN1(n342), .IN2(n341), .QN(N169) );
  NAND2X0 U178 ( .IN1(n346), .IN2(n345), .QN(N170) );
  NAND2X0 U179 ( .IN1(n352), .IN2(n351), .QN(N171) );
  NAND2X0 U180 ( .IN1(n362), .IN2(n361), .QN(N173) );
  NAND2X0 U181 ( .IN1(n369), .IN2(n368), .QN(N174) );
  NAND2X0 U182 ( .IN1(n374), .IN2(n373), .QN(N175) );
  INVX0 U183 ( .INP(n391), .ZN(n390) );
  NOR2X0 U184 ( .IN1(n817), .IN2(n844), .QN(n818) );
  NOR2X0 U185 ( .IN1(n816), .IN2(n815), .QN(n819) );
  INVX0 U186 ( .INP(n561), .ZN(n821) );
  INVX0 U187 ( .INP(n417), .ZN(n489) );
  NOR2X0 U188 ( .IN1(n718), .IN2(n815), .QN(n804) );
  INVX0 U189 ( .INP(n812), .ZN(n802) );
  INVX0 U190 ( .INP(n791), .ZN(n803) );
  INVX0 U191 ( .INP(n792), .ZN(n781) );
  INVX0 U192 ( .INP(n759), .ZN(n772) );
  NOR2X0 U193 ( .IN1(n564), .IN2(n567), .QN(n703) );
  NOR2X0 U194 ( .IN1(n565), .IN2(n567), .QN(n704) );
  INVX0 U195 ( .INP(n735), .ZN(n748) );
  INVX0 U196 ( .INP(n454), .ZN(n563) );
  INVX0 U197 ( .INP(n562), .ZN(n512) );
  INVX0 U198 ( .INP(n743), .ZN(n756) );
  NOR2X0 U199 ( .IN1(n568), .IN2(n567), .QN(n706) );
  INVX0 U200 ( .INP(n689), .ZN(n700) );
  NAND2X0 U201 ( .IN1(exp_diff_value[2]), .IN2(n4), .QN(n214) );
  INVX0 U202 ( .INP(n197), .ZN(n185) );
  INVX0 U203 ( .INP(n196), .ZN(n193) );
  NOR2X0 U204 ( .IN1(n363), .IN2(n74), .QN(n817) );
  INVX0 U205 ( .INP(n308), .ZN(n359) );
  NOR2X0 U206 ( .IN1(exp_diff_value[1]), .IN2(exp_diff_value[0]), .QN(n370) );
  INVX0 U207 ( .INP(n176), .ZN(n698) );
  INVX0 U208 ( .INP(n396), .ZN(n492) );
  NOR2X0 U209 ( .IN1(add_sub_result_24_), .IN2(n393), .QN(n568) );
  MUX21X1 U210 ( .IN1(add_result[24]), .IN2(sub_result[24]), .S(n20), .Q(
        add_sub_result_24_) );
  INVX0 U211 ( .INP(n394), .ZN(n482) );
  INVX0 U212 ( .INP(n21), .ZN(n20) );
  INVX0 U213 ( .INP(n501), .ZN(n21) );
  INVX0 U214 ( .INP(n727), .ZN(n740) );
  INVX0 U215 ( .INP(n751), .ZN(n764) );
  INVX0 U216 ( .INP(n784), .ZN(n771) );
  INVX0 U217 ( .INP(n783), .ZN(n801) );
  INVX0 U218 ( .INP(n811), .ZN(n797) );
  INVX0 U219 ( .INP(n813), .ZN(n805) );
  MUX21X1 U220 ( .IN1(input_factor_01[31]), .IN2(n547), .S(input_factor_02[31]), .Q(n501) );
  INVX0 U221 ( .INP(input_factor_01[31]), .ZN(n547) );
  INVX0 U222 ( .INP(n373), .ZN(n363) );
  NAND2X0 U223 ( .IN1(input_factor_02[29]), .IN2(n599), .QN(n46) );
  INVX0 U224 ( .INP(input_factor_02[23]), .ZN(n557) );
  INVX0 U225 ( .INP(input_factor_02[29]), .ZN(n600) );
  NAND4X0 U226 ( .IN1(n29), .IN2(n28), .IN3(n543), .IN4(n32), .QN(n373) );
  INVX0 U227 ( .INP(n445), .ZN(n713) );
  INVX0 U228 ( .INP(n719), .ZN(n732) );
  INVX0 U229 ( .INP(n440), .ZN(n724) );
  INVX0 U230 ( .INP(n814), .ZN(n800) );
  NOR2X0 U231 ( .IN1(n15), .IN2(n16), .QN(n221) );
  NOR2X0 U232 ( .IN1(n355), .IN2(n252), .QN(n15) );
  NOR2X0 U233 ( .IN1(n11), .IN2(n12), .QN(n276) );
  NOR2X0 U234 ( .IN1(n271), .IN2(n272), .QN(n11) );
  NOR2X0 U235 ( .IN1(n13), .IN2(n14), .QN(n255) );
  NOR2X0 U236 ( .IN1(n365), .IN2(n252), .QN(n13) );
  NOR2X0 U237 ( .IN1(n646), .IN2(n645), .QN(n7) );
  NOR2X0 U238 ( .IN1(n691), .IN2(n690), .QN(n5) );
  NOR2X0 U239 ( .IN1(n606), .IN2(n605), .QN(n9) );
  NAND3X0 U240 ( .IN1(n492), .IN2(n399), .IN3(n463), .QN(n481) );
  OR2X1 U241 ( .IN1(n559), .IN2(n748), .Q(n780) );
  NOR2X0 U242 ( .IN1(n17), .IN2(n18), .QN(n211) );
  NOR2X0 U243 ( .IN1(n684), .IN2(n198), .QN(n17) );
  INVX0 U244 ( .INP(n370), .ZN(n19) );
  NOR4X0 U245 ( .IN1(n389), .IN2(n388), .IN3(n387), .IN4(n386), .QN(n689) );
  MUX21X1 U246 ( .IN1(add_result[1]), .IN2(sub_result[1]), .S(n501), .Q(n811)
         );
  INVX0 U247 ( .INP(input_factor_01[29]), .ZN(n599) );
  OA222X1 U248 ( .IN1(input_factor_02[29]), .IN2(n599), .IN3(n600), .IN4(
        input_factor_01[29]), .IN5(input_factor_01[23]), .IN6(n557), .Q(n29)
         );
  INVX0 U249 ( .INP(input_factor_01[25]), .ZN(n542) );
  INVX0 U250 ( .INP(n33), .ZN(n27) );
  NOR2X0 U251 ( .IN1(input_factor_02[25]), .IN2(n542), .QN(n38) );
  INVX0 U252 ( .INP(input_factor_02[28]), .ZN(n594) );
  INVX0 U253 ( .INP(input_factor_02[26]), .ZN(n582) );
  INVX0 U254 ( .INP(input_factor_01[28]), .ZN(n593) );
  INVX0 U255 ( .INP(input_factor_01[26]), .ZN(n581) );
  NAND4X0 U256 ( .IN1(n41), .IN2(n31), .IN3(n45), .IN4(n22), .QN(n26) );
  INVX0 U257 ( .INP(input_factor_01[27]), .ZN(n587) );
  INVX0 U258 ( .INP(input_factor_02[27]), .ZN(n588) );
  INVX0 U259 ( .INP(input_factor_01[24]), .ZN(n541) );
  NOR2X0 U260 ( .IN1(n541), .IN2(input_factor_02[24]), .QN(n36) );
  INVX0 U261 ( .INP(n36), .ZN(n23) );
  NAND4X0 U262 ( .IN1(n24), .IN2(n30), .IN3(n34), .IN4(n23), .QN(n25) );
  NOR4X0 U263 ( .IN1(n27), .IN2(n38), .IN3(n26), .IN4(n25), .QN(n28) );
  INVX0 U264 ( .INP(input_factor_01[30]), .ZN(n543) );
  INVX0 U265 ( .INP(n30), .ZN(n44) );
  INVX0 U266 ( .INP(n31), .ZN(n40) );
  INVX0 U267 ( .INP(n32), .ZN(n35) );
  OA221X1 U268 ( .IN1(n36), .IN2(n35), .IN3(n36), .IN4(n34), .IN5(n33), .Q(n37) );
  OA22X1 U269 ( .IN1(n38), .IN2(n37), .IN3(input_factor_01[26]), .IN4(n582), 
        .Q(n39) );
  OA22X1 U270 ( .IN1(n40), .IN2(n39), .IN3(input_factor_01[27]), .IN4(n588), 
        .Q(n43) );
  INVX0 U271 ( .INP(n41), .ZN(n42) );
  AO221X1 U272 ( .IN1(n45), .IN2(n44), .IN3(n45), .IN4(n43), .IN5(n42), .Q(n47) );
  AO221X1 U273 ( .IN1(n47), .IN2(n46), .IN3(n600), .IN4(input_factor_01[29]), 
        .IN5(input_factor_01[30]), .Q(n74) );
  INVX0 U274 ( .INP(input_factor_02[22]), .ZN(n702) );
  INVX0 U275 ( .INP(input_factor_02[21]), .ZN(n693) );
  INVX0 U276 ( .INP(input_factor_02[18]), .ZN(n678) );
  INVX0 U277 ( .INP(input_factor_02[17]), .ZN(n672) );
  INVX0 U278 ( .INP(input_factor_02[16]), .ZN(n666) );
  INVX0 U279 ( .INP(input_factor_02[15]), .ZN(n660) );
  INVX0 U280 ( .INP(input_factor_02[14]), .ZN(n654) );
  INVX0 U281 ( .INP(input_factor_02[13]), .ZN(n648) );
  INVX0 U282 ( .INP(input_factor_02[10]), .ZN(n633) );
  INVX0 U283 ( .INP(input_factor_02[9]), .ZN(n627) );
  INVX0 U284 ( .INP(input_factor_02[8]), .ZN(n623) );
  INVX0 U285 ( .INP(input_factor_02[7]), .ZN(n274) );
  INVX0 U286 ( .INP(input_factor_02[6]), .ZN(n254) );
  INVX0 U287 ( .INP(input_factor_02[5]), .ZN(n614) );
  INVX0 U288 ( .INP(input_factor_02[4]), .ZN(n220) );
  INVX0 U289 ( .INP(input_factor_02[3]), .ZN(n189) );
  INVX0 U290 ( .INP(input_factor_02[2]), .ZN(n160) );
  INVX0 U291 ( .INP(input_factor_02[0]), .ZN(n76) );
  AO21X1 U292 ( .IN1(input_factor_01[0]), .IN2(n76), .IN3(input_factor_01[1]), 
        .Q(n48) );
  AO222X1 U293 ( .IN1(input_factor_01[2]), .IN2(n160), .IN3(input_factor_01[2]), .IN4(n48), .IN5(n160), .IN6(n48), .Q(n49) );
  AO222X1 U294 ( .IN1(input_factor_01[3]), .IN2(n189), .IN3(input_factor_01[3]), .IN4(n49), .IN5(n189), .IN6(n49), .Q(n50) );
  AO222X1 U295 ( .IN1(input_factor_01[4]), .IN2(n220), .IN3(input_factor_01[4]), .IN4(n50), .IN5(n220), .IN6(n50), .Q(n51) );
  AO222X1 U296 ( .IN1(input_factor_01[5]), .IN2(n614), .IN3(input_factor_01[5]), .IN4(n51), .IN5(n614), .IN6(n51), .Q(n52) );
  AO222X1 U297 ( .IN1(input_factor_01[6]), .IN2(n254), .IN3(input_factor_01[6]), .IN4(n52), .IN5(n254), .IN6(n52), .Q(n53) );
  AO222X1 U298 ( .IN1(input_factor_01[7]), .IN2(n274), .IN3(input_factor_01[7]), .IN4(n53), .IN5(n274), .IN6(n53), .Q(n54) );
  AO222X1 U299 ( .IN1(input_factor_01[8]), .IN2(n623), .IN3(input_factor_01[8]), .IN4(n54), .IN5(n623), .IN6(n54), .Q(n55) );
  AO222X1 U300 ( .IN1(input_factor_01[9]), .IN2(n627), .IN3(input_factor_01[9]), .IN4(n55), .IN5(n627), .IN6(n55), .Q(n56) );
  AO222X1 U301 ( .IN1(input_factor_01[10]), .IN2(n633), .IN3(
        input_factor_01[10]), .IN4(n56), .IN5(n633), .IN6(n56), .Q(n58) );
  INVX0 U302 ( .INP(input_factor_01[11]), .ZN(n638) );
  INVX0 U303 ( .INP(input_factor_02[11]), .ZN(n639) );
  AO221X1 U304 ( .IN1(n58), .IN2(n57), .IN3(n639), .IN4(input_factor_01[11]), 
        .IN5(input_factor_01[12]), .Q(n59) );
  AO222X1 U305 ( .IN1(input_factor_01[13]), .IN2(n648), .IN3(
        input_factor_01[13]), .IN4(n59), .IN5(n648), .IN6(n59), .Q(n60) );
  AO222X1 U306 ( .IN1(input_factor_01[14]), .IN2(n654), .IN3(
        input_factor_01[14]), .IN4(n60), .IN5(n654), .IN6(n60), .Q(n61) );
  AO222X1 U307 ( .IN1(input_factor_01[15]), .IN2(n660), .IN3(
        input_factor_01[15]), .IN4(n61), .IN5(n660), .IN6(n61), .Q(n62) );
  AO222X1 U308 ( .IN1(input_factor_01[16]), .IN2(n666), .IN3(
        input_factor_01[16]), .IN4(n62), .IN5(n666), .IN6(n62), .Q(n63) );
  AO222X1 U309 ( .IN1(input_factor_01[17]), .IN2(n672), .IN3(
        input_factor_01[17]), .IN4(n63), .IN5(n672), .IN6(n63), .Q(n64) );
  AO222X1 U310 ( .IN1(input_factor_01[18]), .IN2(n678), .IN3(
        input_factor_01[18]), .IN4(n64), .IN5(n678), .IN6(n64), .Q(n66) );
  INVX0 U311 ( .INP(input_factor_01[19]), .ZN(n683) );
  INVX0 U312 ( .INP(input_factor_02[19]), .ZN(n684) );
  AO221X1 U313 ( .IN1(n66), .IN2(n65), .IN3(n684), .IN4(input_factor_01[19]), 
        .IN5(input_factor_01[20]), .Q(n67) );
  AO222X1 U314 ( .IN1(input_factor_01[21]), .IN2(n693), .IN3(
        input_factor_01[21]), .IN4(n67), .IN5(n693), .IN6(n67), .Q(n68) );
  AO222X1 U315 ( .IN1(input_factor_01[22]), .IN2(n702), .IN3(
        input_factor_01[22]), .IN4(n68), .IN5(n702), .IN6(n68), .Q(n69) );
  INVX0 U316 ( .INP(input_factor_01[1]), .ZN(n143) );
  NOR2X0 U317 ( .IN1(n390), .IN2(n143), .QN(N177) );
  INVX0 U318 ( .INP(input_factor_01[12]), .ZN(n644) );
  NOR2X0 U319 ( .IN1(n390), .IN2(n644), .QN(N188) );
  INVX0 U320 ( .INP(input_factor_01[20]), .ZN(n546) );
  NOR2X0 U321 ( .IN1(n390), .IN2(n546), .QN(N196) );
  AO22X1 U322 ( .IN1(input_factor_01[30]), .IN2(rst_n), .IN3(n844), .IN4(
        larger_exponent[7]), .Q(n822) );
  NOR2X0 U324 ( .IN1(n373), .IN2(n69), .QN(n308) );
  OA22X1 U325 ( .IN1(n678), .IN2(n196), .IN3(n672), .IN4(n197), .Q(n71) );
  NAND3X0 U326 ( .IN1(n19), .IN2(n147), .IN3(n120), .QN(n356) );
  MUX21X1 U327 ( .IN1(n211), .IN2(n356), .S(exp_diff_value[2]), .Q(n335) );
  AO22X1 U328 ( .IN1(input_factor_01[18]), .IN2(n193), .IN3(
        input_factor_01[16]), .IN4(n370), .Q(n73) );
  INVX0 U329 ( .INP(n198), .ZN(n192) );
  AO22X1 U330 ( .IN1(input_factor_01[19]), .IN2(n192), .IN3(
        input_factor_01[17]), .IN4(n185), .Q(n72) );
  NOR2X0 U331 ( .IN1(n73), .IN2(n72), .QN(n208) );
  INVX0 U332 ( .INP(input_factor_01[22]), .ZN(n699) );
  INVX0 U333 ( .INP(input_factor_01[21]), .ZN(n692) );
  AO222X1 U334 ( .IN1(n193), .IN2(n699), .IN3(n185), .IN4(n692), .IN5(n370), 
        .IN6(n546), .Q(n355) );
  MUX21X1 U335 ( .IN1(n208), .IN2(n355), .S(exp_diff_value[2]), .Q(n336) );
  INVX0 U336 ( .INP(n817), .ZN(n816) );
  OA22X1 U337 ( .IN1(n335), .IN2(n176), .IN3(n336), .IN4(n816), .Q(n77) );
  NOR3X0 U338 ( .IN1(exp_diff_value[5]), .IN2(exp_diff_value[6]), .IN3(
        exp_diff_value[7]), .QN(n75) );
  AND2X1 U339 ( .IN1(exp_diff_value[4]), .IN2(n75), .Q(n268) );
  OA22X1 U340 ( .IN1(n77), .IN2(n177), .IN3(n76), .IN4(n360), .Q(n118) );
  AO22X1 U341 ( .IN1(input_factor_01[10]), .IN2(n193), .IN3(input_factor_01[8]), .IN4(n370), .Q(n80) );
  AO22X1 U342 ( .IN1(input_factor_01[11]), .IN2(n192), .IN3(input_factor_01[9]), .IN4(n185), .Q(n79) );
  NOR2X0 U343 ( .IN1(n80), .IN2(n79), .QN(n210) );
  AO22X1 U344 ( .IN1(input_factor_01[14]), .IN2(n193), .IN3(
        input_factor_01[12]), .IN4(n370), .Q(n82) );
  AO22X1 U345 ( .IN1(input_factor_01[15]), .IN2(n192), .IN3(
        input_factor_01[13]), .IN4(n185), .Q(n81) );
  NOR2X0 U346 ( .IN1(n82), .IN2(n81), .QN(n209) );
  MUX21X1 U347 ( .IN1(n210), .IN2(n209), .S(exp_diff_value[2]), .Q(n283) );
  AO22X1 U348 ( .IN1(input_factor_01[2]), .IN2(n193), .IN3(input_factor_01[0]), 
        .IN4(n370), .Q(n84) );
  AO22X1 U349 ( .IN1(input_factor_01[3]), .IN2(n192), .IN3(input_factor_01[1]), 
        .IN4(n185), .Q(n83) );
  NOR2X0 U350 ( .IN1(n84), .IN2(n83), .QN(n87) );
  AO22X1 U351 ( .IN1(input_factor_01[6]), .IN2(n193), .IN3(input_factor_01[4]), 
        .IN4(n370), .Q(n86) );
  AO22X1 U352 ( .IN1(input_factor_01[7]), .IN2(n192), .IN3(input_factor_01[5]), 
        .IN4(n185), .Q(n85) );
  NOR2X0 U353 ( .IN1(n86), .IN2(n85), .QN(n216) );
  OA222X1 U354 ( .IN1(n4), .IN2(n283), .IN3(n275), .IN4(n87), .IN5(n214), 
        .IN6(n216), .Q(n116) );
  NOR4X0 U355 ( .IN1(exp_diff_value[4]), .IN2(exp_diff_value[5]), .IN3(
        exp_diff_value[6]), .IN4(exp_diff_value[7]), .QN(n372) );
  AO222X1 U356 ( .IN1(input_factor_02[0]), .IN2(n370), .IN3(input_factor_02[3]), .IN4(n192), .IN5(input_factor_02[2]), .IN6(n193), .Q(n92) );
  INVX0 U357 ( .INP(n275), .ZN(n371) );
  OA22X1 U358 ( .IN1(n633), .IN2(n196), .IN3(n623), .IN4(n19), .Q(n89) );
  OA22X1 U359 ( .IN1(n639), .IN2(n198), .IN3(n627), .IN4(n197), .Q(n88) );
  AO222X1 U360 ( .IN1(input_factor_02[15]), .IN2(n192), .IN3(
        input_factor_02[13]), .IN4(n185), .IN5(input_factor_02[14]), .IN6(n193), .Q(n213) );
  MUX21X1 U361 ( .IN1(n215), .IN2(n213), .S(exp_diff_value[2]), .Q(n281) );
  OA22X1 U362 ( .IN1(n254), .IN2(n196), .IN3(n220), .IN4(n19), .Q(n91) );
  OA22X1 U363 ( .IN1(n614), .IN2(n197), .IN3(n274), .IN4(n198), .Q(n90) );
  INVX0 U364 ( .INP(n214), .ZN(n207) );
  AOI222X1 U365 ( .IN1(n92), .IN2(n371), .IN3(exp_diff_value[3]), .IN4(n281), 
        .IN5(n217), .IN6(n207), .QN(n93) );
  OA22X1 U366 ( .IN1(n116), .IN2(n271), .IN3(n93), .IN4(n232), .Q(n117) );
  NAND3X0 U367 ( .IN1(n119), .IN2(n118), .IN3(n117), .QN(N152) );
  AO222X1 U368 ( .IN1(input_factor_02[18]), .IN2(n185), .IN3(
        input_factor_02[19]), .IN4(n193), .IN5(input_factor_02[17]), .IN6(n370), .Q(n229) );
  INVX0 U369 ( .INP(n229), .ZN(n121) );
  AOI22X1 U370 ( .IN1(input_factor_02[22]), .IN2(n185), .IN3(n3), .IN4(n120), 
        .QN(n358) );
  MUX21X1 U371 ( .IN1(n121), .IN2(n358), .S(exp_diff_value[2]), .Q(n339) );
  AO22X1 U372 ( .IN1(input_factor_01[19]), .IN2(n193), .IN3(
        input_factor_01[17]), .IN4(n370), .Q(n123) );
  AO22X1 U373 ( .IN1(input_factor_01[20]), .IN2(n192), .IN3(
        input_factor_01[18]), .IN4(n185), .Q(n122) );
  NOR2X0 U374 ( .IN1(n123), .IN2(n122), .QN(n226) );
  AO22X1 U375 ( .IN1(input_factor_01[22]), .IN2(n185), .IN3(
        input_factor_01[21]), .IN4(n3), .Q(n124) );
  NOR2X0 U376 ( .IN1(n193), .IN2(n124), .QN(n357) );
  MUX21X1 U377 ( .IN1(n226), .IN2(n357), .S(exp_diff_value[2]), .Q(n340) );
  OA22X1 U378 ( .IN1(n176), .IN2(n339), .IN3(n816), .IN4(n340), .Q(n132) );
  AO222X1 U379 ( .IN1(input_factor_02[10]), .IN2(n185), .IN3(
        input_factor_02[9]), .IN4(n370), .IN5(input_factor_02[11]), .IN6(n193), 
        .Q(n231) );
  OA22X1 U380 ( .IN1(n660), .IN2(n196), .IN3(n648), .IN4(n19), .Q(n126) );
  OA22X1 U381 ( .IN1(n654), .IN2(n197), .IN3(n666), .IN4(n198), .Q(n125) );
  MUX21X1 U382 ( .IN1(n231), .IN2(n230), .S(exp_diff_value[2]), .Q(n127) );
  INVX0 U383 ( .INP(n127), .ZN(n287) );
  OA222X1 U384 ( .IN1(n160), .IN2(n197), .IN3(n189), .IN4(n196), .IN5(n220), 
        .IN6(n198), .Q(n130) );
  AO22X1 U385 ( .IN1(input_factor_02[5]), .IN2(n370), .IN3(input_factor_02[7]), 
        .IN4(n193), .Q(n129) );
  AO22X1 U386 ( .IN1(input_factor_02[6]), .IN2(n185), .IN3(input_factor_02[8]), 
        .IN4(n192), .Q(n128) );
  NOR2X0 U387 ( .IN1(n129), .IN2(n128), .QN(n233) );
  OA222X1 U388 ( .IN1(n4), .IN2(n287), .IN3(n275), .IN4(n130), .IN5(n214), 
        .IN6(n233), .Q(n131) );
  OA22X1 U389 ( .IN1(n132), .IN2(n177), .IN3(n131), .IN4(n232), .Q(n146) );
  AO22X1 U390 ( .IN1(input_factor_01[11]), .IN2(n193), .IN3(input_factor_01[9]), .IN4(n370), .Q(n134) );
  AO22X1 U391 ( .IN1(input_factor_01[12]), .IN2(n192), .IN3(
        input_factor_01[10]), .IN4(n185), .Q(n133) );
  NOR2X0 U392 ( .IN1(n134), .IN2(n133), .QN(n228) );
  AO22X1 U393 ( .IN1(input_factor_01[15]), .IN2(n193), .IN3(
        input_factor_01[13]), .IN4(n370), .Q(n136) );
  AO22X1 U394 ( .IN1(input_factor_01[16]), .IN2(n192), .IN3(
        input_factor_01[14]), .IN4(n185), .Q(n135) );
  NOR2X0 U395 ( .IN1(n136), .IN2(n135), .QN(n227) );
  MUX21X1 U396 ( .IN1(n228), .IN2(n227), .S(exp_diff_value[2]), .Q(n288) );
  AO22X1 U397 ( .IN1(input_factor_01[3]), .IN2(n193), .IN3(input_factor_01[1]), 
        .IN4(n370), .Q(n139) );
  AO22X1 U398 ( .IN1(input_factor_01[4]), .IN2(n192), .IN3(input_factor_01[2]), 
        .IN4(n185), .Q(n137) );
  NOR2X0 U399 ( .IN1(n139), .IN2(n137), .QN(n142) );
  AO22X1 U400 ( .IN1(input_factor_01[7]), .IN2(n193), .IN3(input_factor_01[5]), 
        .IN4(n370), .Q(n141) );
  AO22X1 U401 ( .IN1(input_factor_01[8]), .IN2(n192), .IN3(input_factor_01[6]), 
        .IN4(n185), .Q(n140) );
  NOR2X0 U402 ( .IN1(n141), .IN2(n140), .QN(n234) );
  OA222X1 U403 ( .IN1(n4), .IN2(n288), .IN3(n275), .IN4(n142), .IN5(n214), 
        .IN6(n234), .Q(n144) );
  OA22X1 U404 ( .IN1(n144), .IN2(n271), .IN3(n143), .IN4(n359), .Q(n145) );
  OA222X1 U405 ( .IN1(n693), .IN2(n198), .IN3(n678), .IN4(n19), .IN5(n684), 
        .IN6(n197), .Q(n244) );
  MUX21X1 U406 ( .IN1(n244), .IN2(n367), .S(exp_diff_value[2]), .Q(n343) );
  AO22X1 U407 ( .IN1(input_factor_01[20]), .IN2(n193), .IN3(
        input_factor_01[18]), .IN4(n370), .Q(n149) );
  AO22X1 U408 ( .IN1(input_factor_01[21]), .IN2(n192), .IN3(
        input_factor_01[19]), .IN4(n185), .Q(n148) );
  NOR2X0 U409 ( .IN1(n149), .IN2(n148), .QN(n241) );
  AO21X1 U410 ( .IN1(n699), .IN2(n3), .IN3(exp_diff_value[1]), .Q(n365) );
  MUX21X1 U411 ( .IN1(n241), .IN2(n365), .S(exp_diff_value[2]), .Q(n344) );
  OA22X1 U412 ( .IN1(n343), .IN2(n176), .IN3(n344), .IN4(n816), .Q(n150) );
  OA22X1 U413 ( .IN1(n150), .IN2(n177), .IN3(n160), .IN4(n360), .Q(n171) );
  AO22X1 U414 ( .IN1(input_factor_01[12]), .IN2(n193), .IN3(
        input_factor_01[10]), .IN4(n370), .Q(n152) );
  AO22X1 U415 ( .IN1(input_factor_01[13]), .IN2(n192), .IN3(
        input_factor_01[11]), .IN4(n185), .Q(n151) );
  NOR2X0 U416 ( .IN1(n152), .IN2(n151), .QN(n243) );
  AO22X1 U417 ( .IN1(input_factor_01[16]), .IN2(n193), .IN3(
        input_factor_01[14]), .IN4(n370), .Q(n154) );
  AO22X1 U418 ( .IN1(input_factor_01[17]), .IN2(n192), .IN3(
        input_factor_01[15]), .IN4(n185), .Q(n153) );
  NOR2X0 U419 ( .IN1(n154), .IN2(n153), .QN(n242) );
  MUX21X1 U420 ( .IN1(n243), .IN2(n242), .S(exp_diff_value[2]), .Q(n294) );
  AO22X1 U421 ( .IN1(input_factor_01[4]), .IN2(n193), .IN3(input_factor_01[2]), 
        .IN4(n370), .Q(n156) );
  AO22X1 U422 ( .IN1(input_factor_01[5]), .IN2(n192), .IN3(input_factor_01[3]), 
        .IN4(n185), .Q(n155) );
  NOR2X0 U423 ( .IN1(n156), .IN2(n155), .QN(n159) );
  AO22X1 U424 ( .IN1(input_factor_01[8]), .IN2(n193), .IN3(input_factor_01[6]), 
        .IN4(n370), .Q(n158) );
  AO22X1 U425 ( .IN1(input_factor_01[9]), .IN2(n192), .IN3(input_factor_01[7]), 
        .IN4(n185), .Q(n157) );
  NOR2X0 U426 ( .IN1(n158), .IN2(n157), .QN(n249) );
  OA222X1 U427 ( .IN1(n4), .IN2(n294), .IN3(n275), .IN4(n159), .IN5(n214), 
        .IN6(n249), .Q(n169) );
  OA22X1 U428 ( .IN1(n160), .IN2(n19), .IN3(n220), .IN4(n196), .Q(n162) );
  OA22X1 U429 ( .IN1(n189), .IN2(n197), .IN3(n614), .IN4(n198), .Q(n161) );
  AO222X1 U430 ( .IN1(input_factor_02[10]), .IN2(n370), .IN3(
        input_factor_02[13]), .IN4(n192), .IN5(input_factor_02[11]), .IN6(n185), .Q(n247) );
  OA22X1 U431 ( .IN1(n654), .IN2(n19), .IN3(n666), .IN4(n196), .Q(n164) );
  OA22X1 U432 ( .IN1(n660), .IN2(n197), .IN3(n672), .IN4(n198), .Q(n163) );
  MUX21X1 U433 ( .IN1(n247), .IN2(n246), .S(exp_diff_value[2]), .Q(n292) );
  OA22X1 U434 ( .IN1(n254), .IN2(n19), .IN3(n623), .IN4(n196), .Q(n166) );
  OA22X1 U435 ( .IN1(n274), .IN2(n197), .IN3(n627), .IN4(n198), .Q(n165) );
  AOI222X1 U436 ( .IN1(n167), .IN2(n371), .IN3(exp_diff_value[3]), .IN4(n292), 
        .IN5(n250), .IN6(n207), .QN(n168) );
  OA22X1 U437 ( .IN1(n169), .IN2(n271), .IN3(n168), .IN4(n232), .Q(n170) );
  NAND3X0 U438 ( .IN1(n172), .IN2(n171), .IN3(n170), .QN(N154) );
  AO222X1 U439 ( .IN1(input_factor_02[21]), .IN2(n193), .IN3(
        input_factor_02[19]), .IN4(n370), .IN5(input_factor_02[22]), .IN6(n192), .Q(n264) );
  MUX21X1 U440 ( .IN1(n264), .IN2(n370), .S(exp_diff_value[2]), .Q(n173) );
  INVX0 U441 ( .INP(n173), .ZN(n348) );
  AO22X1 U442 ( .IN1(input_factor_01[21]), .IN2(n193), .IN3(
        input_factor_01[19]), .IN4(n370), .Q(n175) );
  AO22X1 U443 ( .IN1(input_factor_01[22]), .IN2(n192), .IN3(
        input_factor_01[20]), .IN4(n185), .Q(n174) );
  NOR2X0 U444 ( .IN1(n175), .IN2(n174), .QN(n260) );
  MUX21X1 U445 ( .IN1(n260), .IN2(n19), .S(exp_diff_value[2]), .Q(n350) );
  OA22X1 U446 ( .IN1(n348), .IN2(n176), .IN3(n350), .IN4(n816), .Q(n178) );
  OA22X1 U447 ( .IN1(n178), .IN2(n177), .IN3(n189), .IN4(n360), .Q(n205) );
  AO22X1 U448 ( .IN1(input_factor_01[13]), .IN2(n193), .IN3(
        input_factor_01[11]), .IN4(n370), .Q(n180) );
  AO22X1 U449 ( .IN1(input_factor_01[14]), .IN2(n192), .IN3(
        input_factor_01[12]), .IN4(n185), .Q(n179) );
  NOR2X0 U450 ( .IN1(n180), .IN2(n179), .QN(n263) );
  AO22X1 U451 ( .IN1(input_factor_01[17]), .IN2(n193), .IN3(
        input_factor_01[15]), .IN4(n370), .Q(n182) );
  AO22X1 U452 ( .IN1(input_factor_01[18]), .IN2(n192), .IN3(
        input_factor_01[16]), .IN4(n185), .Q(n181) );
  NOR2X0 U453 ( .IN1(n182), .IN2(n181), .QN(n261) );
  MUX21X1 U454 ( .IN1(n263), .IN2(n261), .S(exp_diff_value[2]), .Q(n300) );
  AO22X1 U455 ( .IN1(input_factor_01[5]), .IN2(n193), .IN3(input_factor_01[3]), 
        .IN4(n370), .Q(n184) );
  AO22X1 U456 ( .IN1(input_factor_01[6]), .IN2(n192), .IN3(input_factor_01[4]), 
        .IN4(n185), .Q(n183) );
  NOR2X0 U457 ( .IN1(n184), .IN2(n183), .QN(n188) );
  AO22X1 U458 ( .IN1(input_factor_01[9]), .IN2(n193), .IN3(input_factor_01[7]), 
        .IN4(n370), .Q(n187) );
  AO22X1 U459 ( .IN1(input_factor_01[10]), .IN2(n192), .IN3(input_factor_01[8]), .IN4(n185), .Q(n186) );
  NOR2X0 U460 ( .IN1(n187), .IN2(n186), .QN(n272) );
  OA222X1 U461 ( .IN1(n4), .IN2(n300), .IN3(n275), .IN4(n188), .IN5(n214), 
        .IN6(n272), .Q(n203) );
  OA22X1 U462 ( .IN1(n189), .IN2(n19), .IN3(n614), .IN4(n196), .Q(n191) );
  OA22X1 U463 ( .IN1(n254), .IN2(n198), .IN3(n220), .IN4(n197), .Q(n190) );
  AO222X1 U464 ( .IN1(input_factor_02[11]), .IN2(n370), .IN3(
        input_factor_02[13]), .IN4(n193), .IN5(n192), .IN6(input_factor_02[14]), .Q(n266) );
  OA22X1 U465 ( .IN1(n660), .IN2(n19), .IN3(n672), .IN4(n196), .Q(n195) );
  OA22X1 U466 ( .IN1(n678), .IN2(n198), .IN3(n666), .IN4(n197), .Q(n194) );
  MUX21X1 U467 ( .IN1(n266), .IN2(n265), .S(exp_diff_value[2]), .Q(n298) );
  OA22X1 U468 ( .IN1(n274), .IN2(n19), .IN3(n627), .IN4(n196), .Q(n200) );
  OA22X1 U469 ( .IN1(n633), .IN2(n198), .IN3(n623), .IN4(n197), .Q(n199) );
  AOI222X1 U470 ( .IN1(n201), .IN2(n371), .IN3(exp_diff_value[3]), .IN4(n298), 
        .IN5(n269), .IN6(n207), .QN(n202) );
  OA22X1 U471 ( .IN1(n203), .IN2(n271), .IN3(n202), .IN4(n232), .Q(n204) );
  NAND3X0 U472 ( .IN1(n206), .IN2(n205), .IN3(n204), .QN(N155) );
  INVX0 U473 ( .INP(n271), .ZN(n354) );
  MUX21X1 U474 ( .IN1(n209), .IN2(n208), .S(exp_diff_value[2]), .Q(n305) );
  OA22X1 U475 ( .IN1(n210), .IN2(n262), .IN3(n305), .IN4(n330), .Q(n225) );
  INVX0 U476 ( .INP(n211), .ZN(n212) );
  MUX21X1 U477 ( .IN1(n213), .IN2(n212), .S(exp_diff_value[2]), .Q(n304) );
  NOR2X0 U478 ( .IN1(n4), .IN2(n232), .QN(n307) );
  NOR2X0 U479 ( .IN1(n214), .IN2(n232), .QN(n267) );
  AOI22X1 U480 ( .IN1(n304), .IN2(n307), .IN3(n267), .IN4(n215), .QN(n224) );
  OA22X1 U481 ( .IN1(n216), .IN2(n271), .IN3(n356), .IN4(n248), .Q(n219) );
  INVX0 U482 ( .INP(n232), .ZN(n353) );
  OA22X1 U483 ( .IN1(n221), .IN2(n275), .IN3(n220), .IN4(n360), .Q(n223) );
  NAND4X0 U484 ( .IN1(n225), .IN2(n224), .IN3(n223), .IN4(n222), .QN(N156) );
  MUX21X1 U485 ( .IN1(n227), .IN2(n226), .S(exp_diff_value[2]), .Q(n313) );
  OA22X1 U486 ( .IN1(n228), .IN2(n262), .IN3(n330), .IN4(n313), .Q(n240) );
  MUX21X1 U487 ( .IN1(n230), .IN2(n229), .S(exp_diff_value[2]), .Q(n312) );
  AOI22X1 U488 ( .IN1(n307), .IN2(n312), .IN3(n267), .IN4(n231), .QN(n239) );
  INVX0 U489 ( .INP(input_factor_01[5]), .ZN(n613) );
  OA22X1 U490 ( .IN1(n614), .IN2(n360), .IN3(n613), .IN4(n359), .Q(n238) );
  OA22X1 U491 ( .IN1(n234), .IN2(n271), .IN3(n233), .IN4(n232), .Q(n236) );
  OA22X1 U492 ( .IN1(n357), .IN2(n252), .IN3(n358), .IN4(n248), .Q(n235) );
  AO21X1 U493 ( .IN1(n236), .IN2(n235), .IN3(n275), .Q(n237) );
  NAND4X0 U494 ( .IN1(n240), .IN2(n239), .IN3(n238), .IN4(n237), .QN(N157) );
  MUX21X1 U495 ( .IN1(n242), .IN2(n241), .S(exp_diff_value[2]), .Q(n319) );
  OA22X1 U496 ( .IN1(n243), .IN2(n262), .IN3(n319), .IN4(n330), .Q(n259) );
  INVX0 U497 ( .INP(n244), .ZN(n245) );
  MUX21X1 U498 ( .IN1(n246), .IN2(n245), .S(exp_diff_value[2]), .Q(n318) );
  AOI22X1 U499 ( .IN1(n318), .IN2(n307), .IN3(n267), .IN4(n247), .QN(n258) );
  OA22X1 U500 ( .IN1(n249), .IN2(n271), .IN3(n367), .IN4(n248), .Q(n253) );
  OA22X1 U501 ( .IN1(n255), .IN2(n275), .IN3(n254), .IN4(n360), .Q(n257) );
  NAND4X0 U502 ( .IN1(n259), .IN2(n258), .IN3(n257), .IN4(n256), .QN(N158) );
  MUX21X1 U503 ( .IN1(n261), .IN2(n260), .S(exp_diff_value[2]), .Q(n327) );
  OA22X1 U504 ( .IN1(n263), .IN2(n262), .IN3(n327), .IN4(n330), .Q(n280) );
  MUX21X1 U505 ( .IN1(n265), .IN2(n264), .S(exp_diff_value[2]), .Q(n326) );
  AOI22X1 U506 ( .IN1(n326), .IN2(n307), .IN3(n267), .IN4(n266), .QN(n279) );
  NAND3X0 U507 ( .IN1(n268), .IN2(n370), .IN3(n373), .QN(n273) );
  OA22X1 U508 ( .IN1(n276), .IN2(n275), .IN3(n274), .IN4(n360), .Q(n278) );
  NAND4X0 U509 ( .IN1(n280), .IN2(n279), .IN3(n278), .IN4(n277), .QN(N159) );
  INVX0 U510 ( .INP(n307), .ZN(n329) );
  OA22X1 U511 ( .IN1(n336), .IN2(n330), .IN3(n335), .IN4(n329), .Q(n286) );
  INVX0 U512 ( .INP(n281), .ZN(n282) );
  OA22X1 U513 ( .IN1(n283), .IN2(n349), .IN3(n282), .IN4(n347), .Q(n285) );
  INVX0 U514 ( .INP(input_factor_01[8]), .ZN(n622) );
  OA22X1 U515 ( .IN1(n623), .IN2(n360), .IN3(n622), .IN4(n359), .Q(n284) );
  NAND3X0 U516 ( .IN1(n286), .IN2(n285), .IN3(n284), .QN(N160) );
  OA22X1 U517 ( .IN1(n329), .IN2(n339), .IN3(n330), .IN4(n340), .Q(n291) );
  OA22X1 U518 ( .IN1(n349), .IN2(n288), .IN3(n347), .IN4(n287), .Q(n290) );
  INVX0 U519 ( .INP(input_factor_01[9]), .ZN(n626) );
  OA22X1 U520 ( .IN1(n627), .IN2(n360), .IN3(n626), .IN4(n359), .Q(n289) );
  NAND3X0 U521 ( .IN1(n291), .IN2(n290), .IN3(n289), .QN(N161) );
  OA22X1 U522 ( .IN1(n344), .IN2(n330), .IN3(n343), .IN4(n329), .Q(n297) );
  INVX0 U523 ( .INP(n292), .ZN(n293) );
  OA22X1 U524 ( .IN1(n294), .IN2(n349), .IN3(n293), .IN4(n347), .Q(n296) );
  INVX0 U525 ( .INP(input_factor_01[10]), .ZN(n632) );
  OA22X1 U526 ( .IN1(n633), .IN2(n360), .IN3(n632), .IN4(n359), .Q(n295) );
  NAND3X0 U527 ( .IN1(n297), .IN2(n296), .IN3(n295), .QN(N162) );
  OA22X1 U528 ( .IN1(n350), .IN2(n330), .IN3(n348), .IN4(n329), .Q(n303) );
  INVX0 U529 ( .INP(n298), .ZN(n299) );
  OA22X1 U530 ( .IN1(n300), .IN2(n349), .IN3(n299), .IN4(n347), .Q(n302) );
  OA22X1 U531 ( .IN1(n639), .IN2(n360), .IN3(n638), .IN4(n359), .Q(n301) );
  NAND3X0 U532 ( .IN1(n303), .IN2(n302), .IN3(n301), .QN(N163) );
  INVX0 U533 ( .INP(n304), .ZN(n306) );
  OA22X1 U534 ( .IN1(n306), .IN2(n347), .IN3(n305), .IN4(n349), .Q(n311) );
  OR2X1 U535 ( .IN1(n330), .IN2(exp_diff_value[2]), .Q(n321) );
  OA22X1 U536 ( .IN1(n356), .IN2(n322), .IN3(n355), .IN4(n321), .Q(n310) );
  NAND3X0 U537 ( .IN1(n311), .IN2(n310), .IN3(n309), .QN(N164) );
  INVX0 U538 ( .INP(n312), .ZN(n314) );
  OA22X1 U539 ( .IN1(n314), .IN2(n347), .IN3(n313), .IN4(n349), .Q(n317) );
  OA22X1 U540 ( .IN1(n358), .IN2(n322), .IN3(n357), .IN4(n321), .Q(n316) );
  INVX0 U541 ( .INP(input_factor_01[13]), .ZN(n647) );
  OA22X1 U542 ( .IN1(n648), .IN2(n360), .IN3(n647), .IN4(n359), .Q(n315) );
  NAND3X0 U543 ( .IN1(n317), .IN2(n316), .IN3(n315), .QN(N165) );
  INVX0 U544 ( .INP(n318), .ZN(n320) );
  OA22X1 U545 ( .IN1(n320), .IN2(n347), .IN3(n319), .IN4(n349), .Q(n325) );
  OA22X1 U546 ( .IN1(n367), .IN2(n322), .IN3(n365), .IN4(n321), .Q(n324) );
  INVX0 U547 ( .INP(input_factor_01[14]), .ZN(n653) );
  OA22X1 U548 ( .IN1(n654), .IN2(n360), .IN3(n653), .IN4(n359), .Q(n323) );
  NAND3X0 U549 ( .IN1(n325), .IN2(n324), .IN3(n323), .QN(N166) );
  INVX0 U550 ( .INP(n326), .ZN(n328) );
  OA22X1 U551 ( .IN1(n328), .IN2(n347), .IN3(n327), .IN4(n349), .Q(n334) );
  INVX0 U552 ( .INP(input_factor_01[15]), .ZN(n659) );
  OA22X1 U553 ( .IN1(n660), .IN2(n360), .IN3(n659), .IN4(n359), .Q(n333) );
  NAND3X0 U554 ( .IN1(n331), .IN2(n1), .IN3(n370), .QN(n332) );
  NAND3X0 U555 ( .IN1(n334), .IN2(n333), .IN3(n332), .QN(N167) );
  OA22X1 U556 ( .IN1(n336), .IN2(n349), .IN3(n335), .IN4(n347), .Q(n338) );
  INVX0 U557 ( .INP(input_factor_01[16]), .ZN(n665) );
  OA22X1 U558 ( .IN1(n666), .IN2(n360), .IN3(n665), .IN4(n359), .Q(n337) );
  OA22X1 U559 ( .IN1(n349), .IN2(n340), .IN3(n347), .IN4(n339), .Q(n342) );
  INVX0 U560 ( .INP(input_factor_01[17]), .ZN(n671) );
  OA22X1 U561 ( .IN1(n672), .IN2(n360), .IN3(n671), .IN4(n359), .Q(n341) );
  OA22X1 U562 ( .IN1(n344), .IN2(n349), .IN3(n343), .IN4(n347), .Q(n346) );
  INVX0 U563 ( .INP(input_factor_01[18]), .ZN(n677) );
  OA22X1 U564 ( .IN1(n678), .IN2(n360), .IN3(n677), .IN4(n359), .Q(n345) );
  OA22X1 U565 ( .IN1(n350), .IN2(n349), .IN3(n348), .IN4(n347), .Q(n352) );
  OA22X1 U566 ( .IN1(n684), .IN2(n360), .IN3(n683), .IN4(n359), .Q(n351) );
  OAI222X1 U567 ( .IN1(n366), .IN2(n356), .IN3(n359), .IN4(n546), .IN5(n364), 
        .IN6(n355), .QN(N172) );
  OA22X1 U568 ( .IN1(n358), .IN2(n366), .IN3(n357), .IN4(n364), .Q(n362) );
  OA22X1 U569 ( .IN1(n693), .IN2(n360), .IN3(n692), .IN4(n359), .Q(n361) );
  NAND3X0 U570 ( .IN1(input_factor_01[22]), .IN2(input_factor_02[22]), .IN3(
        n363), .QN(n369) );
  OA22X1 U571 ( .IN1(n367), .IN2(n366), .IN3(n365), .IN4(n364), .Q(n368) );
  NAND3X0 U572 ( .IN1(n372), .IN2(n371), .IN3(n370), .QN(n374) );
  MUX21X1 U573 ( .IN1(input_factor_01[0]), .IN2(input_factor_02[0]), .S(n390), 
        .Q(N176) );
  MUX21X1 U574 ( .IN1(input_factor_01[2]), .IN2(input_factor_02[2]), .S(n390), 
        .Q(N178) );
  MUX21X1 U575 ( .IN1(input_factor_01[3]), .IN2(input_factor_02[3]), .S(n390), 
        .Q(N179) );
  MUX21X1 U576 ( .IN1(input_factor_01[4]), .IN2(input_factor_02[4]), .S(n390), 
        .Q(N180) );
  MUX21X1 U577 ( .IN1(input_factor_01[5]), .IN2(input_factor_02[5]), .S(n390), 
        .Q(N181) );
  MUX21X1 U578 ( .IN1(input_factor_01[6]), .IN2(input_factor_02[6]), .S(n390), 
        .Q(N182) );
  MUX21X1 U579 ( .IN1(input_factor_01[7]), .IN2(input_factor_02[7]), .S(n390), 
        .Q(N183) );
  MUX21X1 U580 ( .IN1(input_factor_01[8]), .IN2(input_factor_02[8]), .S(n390), 
        .Q(N184) );
  MUX21X1 U581 ( .IN1(input_factor_01[9]), .IN2(input_factor_02[9]), .S(n390), 
        .Q(N185) );
  MUX21X1 U582 ( .IN1(input_factor_01[10]), .IN2(input_factor_02[10]), .S(n390), .Q(N186) );
  MUX21X1 U583 ( .IN1(input_factor_01[11]), .IN2(input_factor_02[11]), .S(n390), .Q(N187) );
  MUX21X1 U584 ( .IN1(input_factor_01[13]), .IN2(input_factor_02[13]), .S(n390), .Q(N189) );
  MUX21X1 U585 ( .IN1(input_factor_01[14]), .IN2(input_factor_02[14]), .S(n390), .Q(N190) );
  MUX21X1 U586 ( .IN1(input_factor_01[15]), .IN2(input_factor_02[15]), .S(n390), .Q(N191) );
  MUX21X1 U587 ( .IN1(input_factor_01[16]), .IN2(input_factor_02[16]), .S(n390), .Q(N192) );
  MUX21X1 U588 ( .IN1(input_factor_01[17]), .IN2(input_factor_02[17]), .S(n390), .Q(N193) );
  MUX21X1 U589 ( .IN1(input_factor_01[18]), .IN2(input_factor_02[18]), .S(n390), .Q(N194) );
  MUX21X1 U590 ( .IN1(input_factor_01[19]), .IN2(input_factor_02[19]), .S(n390), .Q(N195) );
  MUX21X1 U591 ( .IN1(input_factor_01[21]), .IN2(input_factor_02[21]), .S(n390), .Q(N197) );
  MUX21X1 U592 ( .IN1(input_factor_01[22]), .IN2(input_factor_02[22]), .S(n390), .Q(N198) );
  MUX21X1 U593 ( .IN1(add_result[0]), .IN2(sub_result[0]), .S(n501), .Q(n813)
         );
  MUX21X1 U594 ( .IN1(add_result[2]), .IN2(sub_result[2]), .S(n501), .Q(n791)
         );
  MUX21X1 U595 ( .IN1(add_result[3]), .IN2(sub_result[3]), .S(n501), .Q(n783)
         );
  MUX21X1 U596 ( .IN1(add_result[4]), .IN2(sub_result[4]), .S(n501), .Q(n792)
         );
  MUX21X1 U597 ( .IN1(add_result[5]), .IN2(sub_result[5]), .S(n501), .Q(n784)
         );
  MUX21X1 U598 ( .IN1(add_result[6]), .IN2(sub_result[6]), .S(n501), .Q(n759)
         );
  MUX21X1 U599 ( .IN1(add_result[7]), .IN2(sub_result[7]), .S(n501), .Q(n751)
         );
  MUX21X1 U600 ( .IN1(add_result[9]), .IN2(sub_result[9]), .S(n501), .Q(n735)
         );
  MUX21X1 U601 ( .IN1(add_result[10]), .IN2(sub_result[10]), .S(n501), .Q(n727) );
  NOR4X0 U602 ( .IN1(n501), .IN2(add_result[14]), .IN3(add_result[15]), .IN4(
        add_result[13]), .QN(n510) );
  NOR4X0 U603 ( .IN1(sub_result[15]), .IN2(sub_result[14]), .IN3(
        sub_result[13]), .IN4(n21), .QN(n508) );
  NOR2X0 U604 ( .IN1(n510), .IN2(n508), .QN(n378) );
  MUX21X1 U605 ( .IN1(add_result[11]), .IN2(sub_result[11]), .S(n501), .Q(n719) );
  MUX21X1 U606 ( .IN1(add_result[16]), .IN2(sub_result[16]), .S(n20), .Q(n394)
         );
  MUX21X1 U607 ( .IN1(add_result[17]), .IN2(sub_result[17]), .S(n20), .Q(n463)
         );
  MUX21X1 U608 ( .IN1(add_result[20]), .IN2(sub_result[20]), .S(n20), .Q(n397)
         );
  INVX0 U609 ( .INP(n397), .ZN(n490) );
  MUX21X1 U610 ( .IN1(add_result[22]), .IN2(sub_result[22]), .S(n20), .Q(n398)
         );
  INVX0 U611 ( .INP(n398), .ZN(n375) );
  MUX21X1 U612 ( .IN1(add_result[23]), .IN2(sub_result[23]), .S(n20), .Q(n393)
         );
  MUX21X1 U613 ( .IN1(add_result[21]), .IN2(sub_result[21]), .S(n20), .Q(n400)
         );
  NOR2X0 U614 ( .IN1(n401), .IN2(n400), .QN(n402) );
  MUX21X1 U615 ( .IN1(add_result[19]), .IN2(sub_result[19]), .S(n20), .Q(n472)
         );
  NOR2X0 U616 ( .IN1(n376), .IN2(n472), .QN(n399) );
  MUX21X1 U617 ( .IN1(add_result[18]), .IN2(sub_result[18]), .S(n20), .Q(n396)
         );
  NOR2X0 U618 ( .IN1(n463), .IN2(n377), .QN(n395) );
  MUX21X1 U619 ( .IN1(add_result[12]), .IN2(sub_result[12]), .S(n20), .Q(n440)
         );
  NOR4X0 U620 ( .IN1(n378), .IN2(n719), .IN3(n562), .IN4(n440), .QN(n714) );
  MUX21X1 U621 ( .IN1(add_result[8]), .IN2(sub_result[8]), .S(n20), .Q(n743)
         );
  NOR3X0 U622 ( .IN1(n735), .IN2(n559), .IN3(n743), .QN(n515) );
  NOR2X0 U623 ( .IN1(n759), .IN2(n379), .QN(n514) );
  NOR2X0 U624 ( .IN1(n792), .IN2(n380), .QN(n522) );
  NOR2X0 U625 ( .IN1(n791), .IN2(n381), .QN(n516) );
  NAND3X0 U626 ( .IN1(n805), .IN2(n797), .IN3(n516), .QN(n560) );
  NAND4X0 U627 ( .IN1(n633), .IN2(n660), .IN3(n639), .IN4(n654), .QN(n389) );
  OR4X1 U628 ( .IN1(input_factor_02[31]), .IN2(input_factor_02[27]), .IN3(
        input_factor_02[24]), .IN4(input_factor_02[25]), .Q(n388) );
  NAND4X0 U629 ( .IN1(n600), .IN2(n557), .IN3(n594), .IN4(n582), .QN(n387) );
  NOR4X0 U630 ( .IN1(input_factor_02[16]), .IN2(input_factor_02[17]), .IN3(
        input_factor_02[19]), .IN4(input_factor_02[22]), .QN(n385) );
  NOR4X0 U631 ( .IN1(input_factor_02[0]), .IN2(input_factor_02[21]), .IN3(
        input_factor_02[13]), .IN4(input_factor_02[18]), .QN(n384) );
  NOR4X0 U632 ( .IN1(input_factor_02[5]), .IN2(input_factor_02[7]), .IN3(
        input_factor_02[8]), .IN4(input_factor_02[9]), .QN(n383) );
  NOR4X0 U633 ( .IN1(input_factor_02[2]), .IN2(input_factor_02[3]), .IN3(
        input_factor_02[6]), .IN4(input_factor_02[4]), .QN(n382) );
  NAND4X0 U634 ( .IN1(n385), .IN2(n384), .IN3(n383), .IN4(n382), .QN(n386) );
  AO222X1 U635 ( .IN1(input_factor_01[31]), .IN2(n689), .IN3(
        input_factor_01[31]), .IN4(n391), .IN5(n390), .IN6(input_factor_02[31]), .Q(n392) );
  AND2X1 U636 ( .IN1(n560), .IN2(n392), .Q(N211) );
  MUX21X1 U637 ( .IN1(n813), .IN2(n811), .S(add_sub_result_24_), .Q(N226) );
  MUX21X1 U638 ( .IN1(n811), .IN2(n791), .S(add_sub_result_24_), .Q(N227) );
  MUX21X1 U639 ( .IN1(n791), .IN2(n783), .S(add_sub_result_24_), .Q(N228) );
  MUX21X1 U640 ( .IN1(n783), .IN2(n792), .S(add_sub_result_24_), .Q(N229) );
  MUX21X1 U641 ( .IN1(n792), .IN2(n784), .S(add_sub_result_24_), .Q(N230) );
  MUX21X1 U642 ( .IN1(n784), .IN2(n759), .S(add_sub_result_24_), .Q(N231) );
  MUX21X1 U643 ( .IN1(n759), .IN2(n751), .S(add_sub_result_24_), .Q(N232) );
  MUX21X1 U644 ( .IN1(n751), .IN2(n743), .S(add_sub_result_24_), .Q(N233) );
  MUX21X1 U645 ( .IN1(n743), .IN2(n735), .S(add_sub_result_24_), .Q(N234) );
  MUX21X1 U646 ( .IN1(n735), .IN2(n727), .S(add_sub_result_24_), .Q(N235) );
  MUX21X1 U647 ( .IN1(n727), .IN2(n719), .S(add_sub_result_24_), .Q(N236) );
  MUX21X1 U648 ( .IN1(n719), .IN2(n440), .S(add_sub_result_24_), .Q(N237) );
  MUX21X1 U649 ( .IN1(add_result[13]), .IN2(sub_result[13]), .S(n20), .Q(n445)
         );
  MUX21X1 U650 ( .IN1(n440), .IN2(n445), .S(add_sub_result_24_), .Q(N238) );
  MUX21X1 U651 ( .IN1(add_result[14]), .IN2(sub_result[14]), .S(n20), .Q(n499)
         );
  MUX21X1 U652 ( .IN1(n445), .IN2(n499), .S(add_sub_result_24_), .Q(N239) );
  MUX21X1 U653 ( .IN1(add_result[15]), .IN2(sub_result[15]), .S(n20), .Q(n454)
         );
  MUX21X1 U654 ( .IN1(n499), .IN2(n454), .S(add_sub_result_24_), .Q(N240) );
  MUX21X1 U655 ( .IN1(n454), .IN2(n394), .S(add_sub_result_24_), .Q(N241) );
  MUX21X1 U656 ( .IN1(n394), .IN2(n463), .S(add_sub_result_24_), .Q(N242) );
  MUX21X1 U657 ( .IN1(n463), .IN2(n396), .S(add_sub_result_24_), .Q(N243) );
  MUX21X1 U658 ( .IN1(n396), .IN2(n472), .S(add_sub_result_24_), .Q(N244) );
  MUX21X1 U659 ( .IN1(n472), .IN2(n397), .S(add_sub_result_24_), .Q(N245) );
  MUX21X1 U660 ( .IN1(n397), .IN2(n400), .S(add_sub_result_24_), .Q(N246) );
  MUX21X1 U661 ( .IN1(n400), .IN2(n398), .S(add_sub_result_24_), .Q(N247) );
  MUX21X1 U662 ( .IN1(n398), .IN2(n393), .S(add_sub_result_24_), .Q(N248) );
  NAND4X0 U663 ( .IN1(n494), .IN2(n483), .IN3(n487), .IN4(n485), .QN(N256) );
  INVX0 U664 ( .INP(n400), .ZN(n486) );
  NOR2X0 U665 ( .IN1(n486), .IN2(n401), .QN(n417) );
  NAND4X0 U666 ( .IN1(n494), .IN2(n481), .IN3(n487), .IN4(n489), .QN(N257) );
  NAND3X0 U667 ( .IN1(n402), .IN2(n490), .IN3(n472), .QN(n491) );
  NAND4X0 U668 ( .IN1(n494), .IN2(n483), .IN3(n491), .IN4(n481), .QN(N258) );
  NOR2X0 U669 ( .IN1(n805), .IN2(n485), .QN(N260) );
  INVX0 U670 ( .INP(n485), .ZN(n419) );
  AO22X1 U671 ( .IN1(n419), .IN2(n811), .IN3(n417), .IN4(n813), .Q(N261) );
  INVX0 U672 ( .INP(n487), .ZN(n418) );
  AO222X1 U673 ( .IN1(n813), .IN2(n418), .IN3(n811), .IN4(n417), .IN5(n791), 
        .IN6(n419), .Q(N262) );
  OA22X1 U674 ( .IN1(n797), .IN2(n487), .IN3(n805), .IN4(n491), .Q(n404) );
  OA22X1 U675 ( .IN1(n803), .IN2(n489), .IN3(n801), .IN4(n485), .Q(n403) );
  OA22X1 U676 ( .IN1(n781), .IN2(n485), .IN3(n801), .IN4(n489), .Q(n407) );
  OA22X1 U677 ( .IN1(n797), .IN2(n491), .IN3(n805), .IN4(n483), .Q(n406) );
  NAND3X0 U678 ( .IN1(n407), .IN2(n406), .IN3(n405), .QN(N264) );
  OA22X1 U679 ( .IN1(n771), .IN2(n485), .IN3(n801), .IN4(n487), .Q(n411) );
  OA22X1 U680 ( .IN1(n803), .IN2(n491), .IN3(n797), .IN4(n483), .Q(n410) );
  INVX0 U681 ( .INP(n481), .ZN(n412) );
  NAND4X0 U682 ( .IN1(n411), .IN2(n410), .IN3(n409), .IN4(n408), .QN(N265) );
  OA22X1 U683 ( .IN1(n781), .IN2(n487), .IN3(n801), .IN4(n491), .Q(n416) );
  OA22X1 U684 ( .IN1(n772), .IN2(n485), .IN3(n771), .IN4(n489), .Q(n415) );
  OA22X1 U685 ( .IN1(n803), .IN2(n483), .IN3(n805), .IN4(n494), .Q(n414) );
  NAND4X0 U686 ( .IN1(n416), .IN2(n415), .IN3(n414), .IN4(n413), .QN(N266) );
  NOR4X0 U687 ( .IN1(n419), .IN2(n418), .IN3(n417), .IN4(N258), .QN(n561) );
  OA22X1 U688 ( .IN1(n803), .IN2(n481), .IN3(n801), .IN4(n483), .Q(n423) );
  OA22X1 U689 ( .IN1(n764), .IN2(n485), .IN3(n771), .IN4(n487), .Q(n422) );
  OA22X1 U690 ( .IN1(n772), .IN2(n489), .IN3(n781), .IN4(n491), .Q(n421) );
  OA22X1 U691 ( .IN1(n797), .IN2(n494), .IN3(n805), .IN4(n821), .Q(n420) );
  NAND4X0 U692 ( .IN1(n423), .IN2(n422), .IN3(n421), .IN4(n420), .QN(N267) );
  OA22X1 U693 ( .IN1(n781), .IN2(n483), .IN3(n801), .IN4(n481), .Q(n427) );
  OA22X1 U694 ( .IN1(n756), .IN2(n485), .IN3(n772), .IN4(n487), .Q(n426) );
  OA22X1 U695 ( .IN1(n764), .IN2(n489), .IN3(n771), .IN4(n491), .Q(n425) );
  OA22X1 U696 ( .IN1(n803), .IN2(n494), .IN3(n797), .IN4(n821), .Q(n424) );
  NAND4X0 U697 ( .IN1(n427), .IN2(n426), .IN3(n425), .IN4(n424), .QN(N268) );
  OA22X1 U698 ( .IN1(n771), .IN2(n483), .IN3(n781), .IN4(n481), .Q(n431) );
  OA22X1 U699 ( .IN1(n748), .IN2(n485), .IN3(n764), .IN4(n487), .Q(n430) );
  OA22X1 U700 ( .IN1(n756), .IN2(n489), .IN3(n772), .IN4(n491), .Q(n429) );
  OA22X1 U701 ( .IN1(n803), .IN2(n821), .IN3(n801), .IN4(n494), .Q(n428) );
  NAND4X0 U702 ( .IN1(n431), .IN2(n430), .IN3(n429), .IN4(n428), .QN(N269) );
  OA22X1 U703 ( .IN1(n772), .IN2(n483), .IN3(n771), .IN4(n481), .Q(n435) );
  OA22X1 U704 ( .IN1(n756), .IN2(n487), .IN3(n740), .IN4(n485), .Q(n434) );
  OA22X1 U705 ( .IN1(n748), .IN2(n489), .IN3(n764), .IN4(n491), .Q(n433) );
  OA22X1 U706 ( .IN1(n781), .IN2(n494), .IN3(n801), .IN4(n821), .Q(n432) );
  NAND4X0 U707 ( .IN1(n435), .IN2(n434), .IN3(n433), .IN4(n432), .QN(N270) );
  OA22X1 U708 ( .IN1(n764), .IN2(n483), .IN3(n772), .IN4(n481), .Q(n439) );
  OA22X1 U709 ( .IN1(n732), .IN2(n485), .IN3(n748), .IN4(n487), .Q(n438) );
  OA22X1 U710 ( .IN1(n756), .IN2(n491), .IN3(n740), .IN4(n489), .Q(n437) );
  OA22X1 U711 ( .IN1(n771), .IN2(n494), .IN3(n781), .IN4(n821), .Q(n436) );
  NAND4X0 U712 ( .IN1(n439), .IN2(n438), .IN3(n437), .IN4(n436), .QN(N271) );
  OA22X1 U713 ( .IN1(n756), .IN2(n483), .IN3(n764), .IN4(n481), .Q(n444) );
  OA22X1 U714 ( .IN1(n724), .IN2(n485), .IN3(n740), .IN4(n487), .Q(n443) );
  OA22X1 U715 ( .IN1(n732), .IN2(n489), .IN3(n748), .IN4(n491), .Q(n442) );
  OA22X1 U716 ( .IN1(n772), .IN2(n494), .IN3(n771), .IN4(n821), .Q(n441) );
  NAND4X0 U717 ( .IN1(n444), .IN2(n443), .IN3(n442), .IN4(n441), .QN(N272) );
  OA22X1 U718 ( .IN1(n756), .IN2(n481), .IN3(n748), .IN4(n483), .Q(n449) );
  OA22X1 U719 ( .IN1(n732), .IN2(n487), .IN3(n713), .IN4(n485), .Q(n448) );
  OA22X1 U720 ( .IN1(n724), .IN2(n489), .IN3(n740), .IN4(n491), .Q(n447) );
  OA22X1 U721 ( .IN1(n764), .IN2(n494), .IN3(n772), .IN4(n821), .Q(n446) );
  NAND4X0 U722 ( .IN1(n449), .IN2(n448), .IN3(n447), .IN4(n446), .QN(N273) );
  OA22X1 U723 ( .IN1(n740), .IN2(n483), .IN3(n748), .IN4(n481), .Q(n453) );
  INVX0 U724 ( .INP(n499), .ZN(n493) );
  OA22X1 U725 ( .IN1(n493), .IN2(n485), .IN3(n724), .IN4(n487), .Q(n452) );
  OA22X1 U726 ( .IN1(n732), .IN2(n491), .IN3(n713), .IN4(n489), .Q(n451) );
  OA22X1 U727 ( .IN1(n756), .IN2(n494), .IN3(n764), .IN4(n821), .Q(n450) );
  NAND4X0 U728 ( .IN1(n453), .IN2(n452), .IN3(n451), .IN4(n450), .QN(N274) );
  OA22X1 U729 ( .IN1(n732), .IN2(n483), .IN3(n740), .IN4(n481), .Q(n458) );
  OA22X1 U730 ( .IN1(n563), .IN2(n485), .IN3(n713), .IN4(n487), .Q(n457) );
  OA22X1 U731 ( .IN1(n493), .IN2(n489), .IN3(n724), .IN4(n491), .Q(n456) );
  OA22X1 U732 ( .IN1(n756), .IN2(n821), .IN3(n748), .IN4(n494), .Q(n455) );
  NAND4X0 U733 ( .IN1(n458), .IN2(n457), .IN3(n456), .IN4(n455), .QN(N275) );
  OA22X1 U734 ( .IN1(n724), .IN2(n483), .IN3(n732), .IN4(n481), .Q(n462) );
  OA22X1 U735 ( .IN1(n493), .IN2(n487), .IN3(n482), .IN4(n485), .Q(n461) );
  OA22X1 U736 ( .IN1(n563), .IN2(n489), .IN3(n713), .IN4(n491), .Q(n460) );
  OA22X1 U737 ( .IN1(n740), .IN2(n494), .IN3(n748), .IN4(n821), .Q(n459) );
  NAND4X0 U738 ( .IN1(n462), .IN2(n461), .IN3(n460), .IN4(n459), .QN(N276) );
  OA22X1 U739 ( .IN1(n724), .IN2(n481), .IN3(n713), .IN4(n483), .Q(n467) );
  INVX0 U740 ( .INP(n463), .ZN(n484) );
  OA22X1 U741 ( .IN1(n563), .IN2(n487), .IN3(n484), .IN4(n485), .Q(n466) );
  OA22X1 U742 ( .IN1(n493), .IN2(n491), .IN3(n482), .IN4(n489), .Q(n465) );
  OA22X1 U743 ( .IN1(n732), .IN2(n494), .IN3(n740), .IN4(n821), .Q(n464) );
  NAND4X0 U744 ( .IN1(n467), .IN2(n466), .IN3(n465), .IN4(n464), .QN(N277) );
  OA22X1 U745 ( .IN1(n493), .IN2(n483), .IN3(n713), .IN4(n481), .Q(n471) );
  OA22X1 U746 ( .IN1(n492), .IN2(n485), .IN3(n482), .IN4(n487), .Q(n470) );
  OA22X1 U747 ( .IN1(n563), .IN2(n491), .IN3(n484), .IN4(n489), .Q(n469) );
  OA22X1 U748 ( .IN1(n724), .IN2(n494), .IN3(n732), .IN4(n821), .Q(n468) );
  NAND4X0 U749 ( .IN1(n471), .IN2(n470), .IN3(n469), .IN4(n468), .QN(N278) );
  OA22X1 U750 ( .IN1(n563), .IN2(n483), .IN3(n493), .IN4(n481), .Q(n476) );
  INVX0 U751 ( .INP(n472), .ZN(n488) );
  OA22X1 U752 ( .IN1(n484), .IN2(n487), .IN3(n488), .IN4(n485), .Q(n475) );
  OA22X1 U753 ( .IN1(n492), .IN2(n489), .IN3(n482), .IN4(n491), .Q(n474) );
  OA22X1 U754 ( .IN1(n724), .IN2(n821), .IN3(n713), .IN4(n494), .Q(n473) );
  NAND4X0 U755 ( .IN1(n476), .IN2(n475), .IN3(n474), .IN4(n473), .QN(N279) );
  OA22X1 U756 ( .IN1(n563), .IN2(n481), .IN3(n482), .IN4(n483), .Q(n480) );
  OA22X1 U757 ( .IN1(n492), .IN2(n487), .IN3(n490), .IN4(n485), .Q(n479) );
  OA22X1 U758 ( .IN1(n484), .IN2(n491), .IN3(n488), .IN4(n489), .Q(n478) );
  OA22X1 U759 ( .IN1(n493), .IN2(n494), .IN3(n713), .IN4(n821), .Q(n477) );
  NAND4X0 U760 ( .IN1(n480), .IN2(n479), .IN3(n478), .IN4(n477), .QN(N280) );
  OA22X1 U761 ( .IN1(n484), .IN2(n483), .IN3(n482), .IN4(n481), .Q(n498) );
  OA22X1 U762 ( .IN1(n488), .IN2(n487), .IN3(n486), .IN4(n485), .Q(n497) );
  OA22X1 U763 ( .IN1(n492), .IN2(n491), .IN3(n490), .IN4(n489), .Q(n496) );
  OA22X1 U764 ( .IN1(n563), .IN2(n494), .IN3(n493), .IN4(n821), .Q(n495) );
  NAND4X0 U765 ( .IN1(n498), .IN2(n497), .IN3(n496), .IN4(n495), .QN(N281) );
  NAND3X0 U766 ( .IN1(n499), .IN2(n512), .IN3(n563), .QN(n712) );
  AO22X1 U767 ( .IN1(n510), .IN2(add_result[12]), .IN3(n508), .IN4(
        sub_result[12]), .Q(n500) );
  INVX0 U768 ( .INP(n712), .ZN(n506) );
  NOR3X0 U769 ( .IN1(n501), .IN2(add_result[14]), .IN3(add_result[15]), .QN(
        n503) );
  NOR3X0 U770 ( .IN1(sub_result[14]), .IN2(sub_result[15]), .IN3(n21), .QN(
        n502) );
  AO22X1 U771 ( .IN1(n503), .IN2(add_result[13]), .IN3(n502), .IN4(
        sub_result[13]), .Q(n504) );
  NOR2X0 U772 ( .IN1(n506), .IN2(n505), .QN(N308) );
  INVX0 U773 ( .INP(add_result[12]), .ZN(n509) );
  INVX0 U774 ( .INP(sub_result[12]), .ZN(n507) );
  AO22X1 U775 ( .IN1(n510), .IN2(n509), .IN3(n508), .IN4(n507), .Q(n511) );
  NAND3X0 U776 ( .IN1(n512), .IN2(n719), .IN3(n511), .QN(n806) );
  NAND4X0 U777 ( .IN1(N308), .IN2(n806), .IN3(n789), .IN4(n780), .QN(n773) );
  NAND4X0 U778 ( .IN1(n789), .IN2(n712), .IN3(n718), .IN4(n773), .QN(N306) );
  NAND4X0 U779 ( .IN1(n780), .IN2(n711), .IN3(n718), .IN4(n773), .QN(N307) );
  AO22X1 U780 ( .IN1(n698), .IN2(exponent_factor_12[0]), .IN3(n817), .IN4(
        exponent_factor_21[0]), .Q(N34) );
  NAND3X0 U781 ( .IN1(n801), .IN2(n522), .IN3(n791), .QN(n535) );
  NAND3X0 U782 ( .IN1(n771), .IN2(n514), .IN3(n792), .QN(n530) );
  NAND3X0 U783 ( .IN1(n764), .IN2(n515), .IN3(n759), .QN(n531) );
  NAND3X0 U784 ( .IN1(n803), .IN2(n797), .IN3(n801), .QN(n513) );
  AND2X1 U785 ( .IN1(n530), .IN2(n532), .Q(n517) );
  NAND4X0 U786 ( .IN1(n519), .IN2(n517), .IN3(n531), .IN4(n533), .QN(n518) );
  NAND4X0 U787 ( .IN1(n535), .IN2(n530), .IN3(n531), .IN4(n518), .QN(N346) );
  NAND3X0 U788 ( .IN1(n517), .IN2(n534), .IN3(n518), .QN(N347) );
  NOR2X0 U789 ( .IN1(n805), .IN2(n533), .QN(N349) );
  AO22X1 U790 ( .IN1(n698), .IN2(exponent_factor_12[1]), .IN3(n817), .IN4(
        exponent_factor_21[1]), .Q(N35) );
  OAI22X1 U791 ( .IN1(n797), .IN2(n533), .IN3(n805), .IN4(n531), .QN(N350) );
  OAI222X1 U792 ( .IN1(n532), .IN2(n805), .IN3(n531), .IN4(n797), .IN5(n533), 
        .IN6(n803), .QN(N351) );
  OA22X1 U793 ( .IN1(n803), .IN2(n531), .IN3(n801), .IN4(n533), .Q(n521) );
  OA22X1 U794 ( .IN1(n797), .IN2(n532), .IN3(n805), .IN4(n530), .Q(n520) );
  OA22X1 U795 ( .IN1(n781), .IN2(n533), .IN3(n801), .IN4(n531), .Q(n525) );
  OA22X1 U796 ( .IN1(n803), .IN2(n532), .IN3(n797), .IN4(n530), .Q(n524) );
  AND2X1 U797 ( .IN1(n522), .IN2(n783), .Q(n536) );
  NAND3X0 U798 ( .IN1(n525), .IN2(n524), .IN3(n523), .QN(N353) );
  OA22X1 U799 ( .IN1(n771), .IN2(n533), .IN3(n781), .IN4(n531), .Q(n529) );
  OA22X1 U800 ( .IN1(n803), .IN2(n530), .IN3(n805), .IN4(n535), .Q(n528) );
  OR2X1 U801 ( .IN1(n532), .IN2(n801), .Q(n526) );
  NAND4X0 U802 ( .IN1(n529), .IN2(n528), .IN3(n527), .IN4(n526), .QN(N354) );
  OA22X1 U803 ( .IN1(n771), .IN2(n531), .IN3(n801), .IN4(n530), .Q(n540) );
  OA22X1 U804 ( .IN1(n772), .IN2(n533), .IN3(n781), .IN4(n532), .Q(n539) );
  OA22X1 U805 ( .IN1(n797), .IN2(n535), .IN3(n805), .IN4(n534), .Q(n538) );
  NAND4X0 U806 ( .IN1(n540), .IN2(n539), .IN3(n538), .IN4(n537), .QN(N355) );
  AO22X1 U807 ( .IN1(n698), .IN2(exponent_factor_12[2]), .IN3(n817), .IN4(
        exponent_factor_21[2]), .Q(N36) );
  AO22X1 U808 ( .IN1(n698), .IN2(exponent_factor_12[3]), .IN3(n817), .IN4(
        exponent_factor_21[3]), .Q(N37) );
  AO22X1 U809 ( .IN1(n698), .IN2(exponent_factor_12[4]), .IN3(n817), .IN4(
        exponent_factor_21[4]), .Q(N38) );
  NAND4X0 U810 ( .IN1(n542), .IN2(n599), .IN3(n587), .IN4(n541), .QN(n545) );
  INVX0 U811 ( .INP(input_factor_01[23]), .ZN(n556) );
  NAND4X0 U812 ( .IN1(n543), .IN2(n556), .IN3(n593), .IN4(n581), .QN(n544) );
  NOR2X0 U813 ( .IN1(n545), .IN2(n544), .QN(n555) );
  NOR4X0 U814 ( .IN1(input_factor_01[7]), .IN2(input_factor_01[6]), .IN3(
        input_factor_01[5]), .IN4(input_factor_01[4]), .QN(n554) );
  NOR4X0 U815 ( .IN1(input_factor_01[3]), .IN2(input_factor_01[2]), .IN3(
        input_factor_01[1]), .IN4(input_factor_01[0]), .QN(n553) );
  NAND4X0 U816 ( .IN1(n699), .IN2(n692), .IN3(n546), .IN4(n683), .QN(n551) );
  NAND4X0 U817 ( .IN1(n547), .IN2(n677), .IN3(n671), .IN4(n665), .QN(n550) );
  NAND4X0 U818 ( .IN1(n659), .IN2(n653), .IN3(n647), .IN4(n644), .QN(n549) );
  NAND4X0 U819 ( .IN1(n638), .IN2(n632), .IN3(n626), .IN4(n622), .QN(n548) );
  NOR4X0 U820 ( .IN1(n551), .IN2(n550), .IN3(n549), .IN4(n548), .QN(n552) );
  NAND4X0 U821 ( .IN1(n555), .IN2(n554), .IN3(n553), .IN4(n552), .QN(n701) );
  OA22X1 U822 ( .IN1(n557), .IN2(n701), .IN3(n700), .IN4(n556), .Q(n572) );
  INVX0 U823 ( .INP(n773), .ZN(n558) );
  OA21X1 U824 ( .IN1(n756), .IN2(n559), .IN3(n558), .Q(n565) );
  NAND3X0 U825 ( .IN1(n560), .IN2(n700), .IN3(n701), .QN(n567) );
  OA21X1 U826 ( .IN1(n563), .IN2(n562), .IN3(n561), .Q(n564) );
  AOI22X1 U827 ( .IN1(n704), .IN2(add_output_exponent_w3[0]), .IN3(n703), 
        .IN4(add_output_exponent_w2[0]), .QN(n571) );
  INVX0 U828 ( .INP(n567), .ZN(n566) );
  AND4X1 U829 ( .IN1(n568), .IN2(n566), .IN3(n565), .IN4(n564), .Q(n705) );
  NAND4X0 U830 ( .IN1(n572), .IN2(n571), .IN3(n570), .IN4(n569), .QN(N380) );
  INVX0 U831 ( .INP(n701), .ZN(n619) );
  AOI22X1 U832 ( .IN1(input_factor_02[24]), .IN2(n619), .IN3(n689), .IN4(
        input_factor_01[24]), .QN(n576) );
  AOI22X1 U833 ( .IN1(n704), .IN2(add_output_exponent_w3[1]), .IN3(n703), 
        .IN4(add_output_exponent_w2[1]), .QN(n575) );
  NAND4X0 U834 ( .IN1(n576), .IN2(n575), .IN3(n574), .IN4(n573), .QN(N381) );
  AOI22X1 U835 ( .IN1(input_factor_02[25]), .IN2(n619), .IN3(n689), .IN4(
        input_factor_01[25]), .QN(n580) );
  AOI22X1 U836 ( .IN1(n704), .IN2(add_output_exponent_w3[2]), .IN3(n703), 
        .IN4(add_output_exponent_w2[2]), .QN(n579) );
  NAND4X0 U837 ( .IN1(n580), .IN2(n579), .IN3(n578), .IN4(n577), .QN(N382) );
  OA22X1 U838 ( .IN1(n582), .IN2(n701), .IN3(n700), .IN4(n581), .Q(n586) );
  AOI22X1 U839 ( .IN1(n704), .IN2(add_output_exponent_w3[3]), .IN3(n703), 
        .IN4(add_output_exponent_w2[3]), .QN(n585) );
  NAND4X0 U840 ( .IN1(n586), .IN2(n585), .IN3(n584), .IN4(n583), .QN(N383) );
  OA22X1 U841 ( .IN1(n588), .IN2(n701), .IN3(n700), .IN4(n587), .Q(n592) );
  AOI22X1 U842 ( .IN1(n704), .IN2(add_output_exponent_w3[4]), .IN3(n703), 
        .IN4(add_output_exponent_w2[4]), .QN(n591) );
  NAND4X0 U843 ( .IN1(n592), .IN2(n591), .IN3(n590), .IN4(n589), .QN(N384) );
  OA22X1 U844 ( .IN1(n594), .IN2(n701), .IN3(n700), .IN4(n593), .Q(n598) );
  AOI22X1 U845 ( .IN1(n704), .IN2(add_output_exponent_w3[5]), .IN3(n703), 
        .IN4(add_output_exponent_w2[5]), .QN(n597) );
  NAND4X0 U846 ( .IN1(n598), .IN2(n597), .IN3(n596), .IN4(n595), .QN(N385) );
  OA22X1 U847 ( .IN1(n600), .IN2(n701), .IN3(n700), .IN4(n599), .Q(n604) );
  AOI22X1 U848 ( .IN1(n704), .IN2(add_output_exponent_w3[6]), .IN3(n703), 
        .IN4(add_output_exponent_w2[6]), .QN(n603) );
  NAND4X0 U849 ( .IN1(n604), .IN2(n603), .IN3(n602), .IN4(n601), .QN(N386) );
  AO22X1 U851 ( .IN1(n689), .IN2(input_factor_01[30]), .IN3(n706), .IN4(
        add_output_exponent_w1[7]), .Q(n606) );
  AO22X1 U852 ( .IN1(n704), .IN2(add_output_exponent_w3[7]), .IN3(n703), .IN4(
        add_output_exponent_w2[7]), .Q(n605) );
  AO222X1 U853 ( .IN1(input_factor_02[0]), .IN2(n619), .IN3(input_factor_01[0]), .IN4(n689), .IN5(n706), .IN6(pre_sig_res_01[0]), .Q(N388) );
  AO222X1 U854 ( .IN1(n689), .IN2(input_factor_01[1]), .IN3(n703), .IN4(
        pre_sig_res_02[1]), .IN5(pre_sig_res_01[1]), .IN6(n706), .Q(N389) );
  AO22X1 U855 ( .IN1(n698), .IN2(exponent_factor_12[5]), .IN3(n817), .IN4(
        exponent_factor_21[5]), .Q(N39) );
  AOI22X1 U856 ( .IN1(n703), .IN2(pre_sig_res_02[2]), .IN3(n706), .IN4(
        pre_sig_res_01[2]), .QN(n608) );
  AOI22X1 U857 ( .IN1(input_factor_02[2]), .IN2(n619), .IN3(n689), .IN4(
        input_factor_01[2]), .QN(n607) );
  AOI22X1 U858 ( .IN1(n703), .IN2(pre_sig_res_02[3]), .IN3(n706), .IN4(
        pre_sig_res_01[3]), .QN(n610) );
  AOI22X1 U859 ( .IN1(input_factor_02[3]), .IN2(n619), .IN3(n689), .IN4(
        input_factor_01[3]), .QN(n609) );
  AOI22X1 U860 ( .IN1(n703), .IN2(pre_sig_res_02[4]), .IN3(n706), .IN4(
        pre_sig_res_01[4]), .QN(n612) );
  AOI22X1 U861 ( .IN1(input_factor_02[4]), .IN2(n619), .IN3(n689), .IN4(
        input_factor_01[4]), .QN(n611) );
  AOI22X1 U862 ( .IN1(n703), .IN2(pre_sig_res_02[5]), .IN3(n706), .IN4(
        pre_sig_res_01[5]), .QN(n616) );
  OA22X1 U863 ( .IN1(n614), .IN2(n701), .IN3(n700), .IN4(n613), .Q(n615) );
  AOI22X1 U864 ( .IN1(n703), .IN2(pre_sig_res_02[6]), .IN3(n706), .IN4(
        pre_sig_res_01[6]), .QN(n618) );
  AOI22X1 U865 ( .IN1(input_factor_02[6]), .IN2(n619), .IN3(n689), .IN4(
        input_factor_01[6]), .QN(n617) );
  AOI22X1 U866 ( .IN1(n703), .IN2(pre_sig_res_02[7]), .IN3(n706), .IN4(
        pre_sig_res_01[7]), .QN(n621) );
  AOI22X1 U867 ( .IN1(input_factor_02[7]), .IN2(n619), .IN3(n689), .IN4(
        input_factor_01[7]), .QN(n620) );
  AOI22X1 U868 ( .IN1(n703), .IN2(pre_sig_res_02[8]), .IN3(n706), .IN4(
        pre_sig_res_01[8]), .QN(n625) );
  OA22X1 U869 ( .IN1(n623), .IN2(n701), .IN3(n700), .IN4(n622), .Q(n624) );
  OA22X1 U870 ( .IN1(n627), .IN2(n701), .IN3(n700), .IN4(n626), .Q(n631) );
  NAND4X0 U871 ( .IN1(n631), .IN2(n630), .IN3(n629), .IN4(n628), .QN(N397) );
  OA22X1 U872 ( .IN1(n633), .IN2(n701), .IN3(n700), .IN4(n632), .Q(n637) );
  NAND4X0 U873 ( .IN1(n637), .IN2(n636), .IN3(n635), .IN4(n634), .QN(N398) );
  OA22X1 U874 ( .IN1(n639), .IN2(n701), .IN3(n700), .IN4(n638), .Q(n643) );
  NAND4X0 U875 ( .IN1(n643), .IN2(n642), .IN3(n641), .IN4(n640), .QN(N399) );
  AO22X1 U876 ( .IN1(n698), .IN2(exponent_factor_12[6]), .IN3(n817), .IN4(
        exponent_factor_21[6]), .Q(N40) );
  NOR2X0 U877 ( .IN1(n700), .IN2(n644), .QN(n646) );
  AO22X1 U878 ( .IN1(n704), .IN2(pre_sig_res_03[12]), .IN3(n703), .IN4(
        pre_sig_res_02[12]), .Q(n645) );
  OA22X1 U879 ( .IN1(n648), .IN2(n701), .IN3(n700), .IN4(n647), .Q(n652) );
  NAND4X0 U880 ( .IN1(n652), .IN2(n651), .IN3(n650), .IN4(n649), .QN(N401) );
  OA22X1 U881 ( .IN1(n654), .IN2(n701), .IN3(n700), .IN4(n653), .Q(n658) );
  NAND4X0 U882 ( .IN1(n658), .IN2(n657), .IN3(n656), .IN4(n655), .QN(N402) );
  OA22X1 U883 ( .IN1(n660), .IN2(n701), .IN3(n700), .IN4(n659), .Q(n664) );
  NAND4X0 U884 ( .IN1(n664), .IN2(n663), .IN3(n662), .IN4(n661), .QN(N403) );
  OA22X1 U885 ( .IN1(n666), .IN2(n701), .IN3(n700), .IN4(n665), .Q(n670) );
  AOI22X1 U886 ( .IN1(n704), .IN2(pre_sig_res_03[16]), .IN3(n703), .IN4(
        pre_sig_res_02[16]), .QN(n669) );
  NAND4X0 U887 ( .IN1(n670), .IN2(n669), .IN3(n668), .IN4(n667), .QN(N404) );
  OA22X1 U888 ( .IN1(n672), .IN2(n701), .IN3(n700), .IN4(n671), .Q(n676) );
  AOI22X1 U889 ( .IN1(n704), .IN2(pre_sig_res_03[17]), .IN3(n703), .IN4(
        pre_sig_res_02[17]), .QN(n675) );
  NAND4X0 U890 ( .IN1(n676), .IN2(n675), .IN3(n674), .IN4(n673), .QN(N405) );
  OA22X1 U891 ( .IN1(n678), .IN2(n701), .IN3(n700), .IN4(n677), .Q(n682) );
  AOI22X1 U892 ( .IN1(n704), .IN2(pre_sig_res_03[18]), .IN3(n703), .IN4(
        pre_sig_res_02[18]), .QN(n681) );
  NAND4X0 U893 ( .IN1(n682), .IN2(n681), .IN3(n680), .IN4(n679), .QN(N406) );
  OA22X1 U894 ( .IN1(n684), .IN2(n701), .IN3(n700), .IN4(n683), .Q(n688) );
  AOI22X1 U895 ( .IN1(n704), .IN2(pre_sig_res_03[19]), .IN3(n703), .IN4(
        pre_sig_res_02[19]), .QN(n687) );
  NAND4X0 U896 ( .IN1(n688), .IN2(n687), .IN3(n686), .IN4(n685), .QN(N407) );
  AO22X1 U897 ( .IN1(n689), .IN2(input_factor_01[20]), .IN3(n706), .IN4(
        pre_sig_res_01[20]), .Q(n691) );
  AO22X1 U898 ( .IN1(n704), .IN2(pre_sig_res_03[20]), .IN3(n703), .IN4(
        pre_sig_res_02[20]), .Q(n690) );
  OA22X1 U899 ( .IN1(n693), .IN2(n701), .IN3(n700), .IN4(n692), .Q(n697) );
  AOI22X1 U900 ( .IN1(n704), .IN2(pre_sig_res_03[21]), .IN3(n703), .IN4(
        pre_sig_res_02[21]), .QN(n696) );
  NAND4X0 U901 ( .IN1(n697), .IN2(n696), .IN3(n695), .IN4(n694), .QN(N409) );
  AO22X1 U902 ( .IN1(n698), .IN2(exponent_factor_12[7]), .IN3(n817), .IN4(
        exponent_factor_21[7]), .Q(N41) );
  OA22X1 U903 ( .IN1(n702), .IN2(n701), .IN3(n700), .IN4(n699), .Q(n710) );
  AOI22X1 U904 ( .IN1(n704), .IN2(pre_sig_res_03[22]), .IN3(n703), .IN4(
        pre_sig_res_02[22]), .QN(n709) );
  NAND4X0 U905 ( .IN1(n710), .IN2(n709), .IN3(n708), .IN4(n707), .QN(N410) );
  NOR2X0 U906 ( .IN1(n844), .IN2(n711), .QN(n812) );
  NOR2X0 U907 ( .IN1(n712), .IN2(n844), .QN(n814) );
  OA22X1 U908 ( .IN1(n724), .IN2(n802), .IN3(n713), .IN4(n800), .Q(n723) );
  OA22X1 U909 ( .IN1(n740), .IN2(n806), .IN3(n764), .IN4(n773), .Q(n717) );
  INVX0 U910 ( .INP(rst_n), .ZN(n815) );
  NAND3X0 U911 ( .IN1(n715), .IN2(n735), .IN3(n714), .QN(n716) );
  OA22X1 U912 ( .IN1(n844), .IN2(n717), .IN3(n815), .IN4(n716), .Q(n722) );
  NAND4X0 U913 ( .IN1(n723), .IN2(n722), .IN3(n721), .IN4(n720), .QN(n843) );
  OA22X1 U914 ( .IN1(n724), .IN2(n800), .IN3(n732), .IN4(n802), .Q(n731) );
  OA22X1 U915 ( .IN1(n764), .IN2(n780), .IN3(n772), .IN4(n773), .Q(n726) );
  OA22X1 U916 ( .IN1(n756), .IN2(n789), .IN3(n748), .IN4(n806), .Q(n725) );
  AO21X1 U917 ( .IN1(n726), .IN2(n725), .IN3(n844), .Q(n730) );
  NAND4X0 U918 ( .IN1(n731), .IN2(n730), .IN3(n729), .IN4(n728), .QN(n842) );
  OA22X1 U919 ( .IN1(n732), .IN2(n800), .IN3(n740), .IN4(n802), .Q(n739) );
  OA22X1 U920 ( .IN1(n772), .IN2(n780), .IN3(n771), .IN4(n773), .Q(n734) );
  OA22X1 U921 ( .IN1(n756), .IN2(n806), .IN3(n764), .IN4(n789), .Q(n733) );
  AO21X1 U922 ( .IN1(n734), .IN2(n733), .IN3(n844), .Q(n738) );
  NAND4X0 U923 ( .IN1(n739), .IN2(n738), .IN3(n737), .IN4(n736), .QN(n841) );
  OA22X1 U924 ( .IN1(n740), .IN2(n800), .IN3(n748), .IN4(n802), .Q(n747) );
  OA22X1 U925 ( .IN1(n771), .IN2(n780), .IN3(n781), .IN4(n773), .Q(n742) );
  OA22X1 U926 ( .IN1(n764), .IN2(n806), .IN3(n772), .IN4(n789), .Q(n741) );
  AO21X1 U927 ( .IN1(n742), .IN2(n741), .IN3(n844), .Q(n746) );
  NAND4X0 U928 ( .IN1(n747), .IN2(n746), .IN3(n745), .IN4(n744), .QN(n840) );
  OA22X1 U929 ( .IN1(n756), .IN2(n802), .IN3(n748), .IN4(n800), .Q(n755) );
  OA22X1 U930 ( .IN1(n781), .IN2(n780), .IN3(n801), .IN4(n773), .Q(n750) );
  OA22X1 U931 ( .IN1(n772), .IN2(n806), .IN3(n771), .IN4(n789), .Q(n749) );
  AO21X1 U932 ( .IN1(n750), .IN2(n749), .IN3(n844), .Q(n754) );
  NAND4X0 U933 ( .IN1(n755), .IN2(n754), .IN3(n753), .IN4(n752), .QN(n839) );
  OA22X1 U934 ( .IN1(n756), .IN2(n800), .IN3(n764), .IN4(n802), .Q(n763) );
  OA22X1 U935 ( .IN1(n803), .IN2(n773), .IN3(n801), .IN4(n780), .Q(n758) );
  OA22X1 U936 ( .IN1(n771), .IN2(n806), .IN3(n781), .IN4(n789), .Q(n757) );
  AO21X1 U937 ( .IN1(n758), .IN2(n757), .IN3(n844), .Q(n762) );
  NAND4X0 U938 ( .IN1(n763), .IN2(n762), .IN3(n761), .IN4(n760), .QN(n838) );
  OA22X1 U939 ( .IN1(n764), .IN2(n800), .IN3(n772), .IN4(n802), .Q(n770) );
  OA22X1 U940 ( .IN1(n803), .IN2(n780), .IN3(n797), .IN4(n773), .Q(n766) );
  OA22X1 U941 ( .IN1(n781), .IN2(n806), .IN3(n801), .IN4(n789), .Q(n765) );
  AO21X1 U942 ( .IN1(n766), .IN2(n765), .IN3(n844), .Q(n769) );
  NAND4X0 U943 ( .IN1(n770), .IN2(n769), .IN3(n768), .IN4(n767), .QN(n837) );
  OA22X1 U944 ( .IN1(n772), .IN2(n800), .IN3(n771), .IN4(n802), .Q(n779) );
  OA22X1 U945 ( .IN1(n797), .IN2(n780), .IN3(n805), .IN4(n773), .Q(n775) );
  OA22X1 U946 ( .IN1(n803), .IN2(n789), .IN3(n801), .IN4(n806), .Q(n774) );
  AO21X1 U947 ( .IN1(n775), .IN2(n774), .IN3(n844), .Q(n778) );
  NAND4X0 U948 ( .IN1(n779), .IN2(n778), .IN3(n777), .IN4(n776), .QN(n836) );
  OA222X1 U949 ( .IN1(n806), .IN2(n803), .IN3(n780), .IN4(n805), .IN5(n789), 
        .IN6(n797), .Q(n782) );
  OA22X1 U950 ( .IN1(n844), .IN2(n782), .IN3(n781), .IN4(n802), .Q(n788) );
  NAND4X0 U951 ( .IN1(n788), .IN2(n787), .IN3(n786), .IN4(n785), .QN(n835) );
  OA22X1 U952 ( .IN1(n797), .IN2(n806), .IN3(n805), .IN4(n789), .Q(n790) );
  OA22X1 U953 ( .IN1(n801), .IN2(n802), .IN3(n790), .IN4(n815), .Q(n796) );
  NAND4X0 U954 ( .IN1(n796), .IN2(n795), .IN3(n794), .IN4(n793), .QN(n834) );
  AOI22X1 U955 ( .IN1(pre_sig_res_03[11]), .IN2(n815), .IN3(n804), .IN4(n813), 
        .QN(n799) );
  OA22X1 U956 ( .IN1(n803), .IN2(n800), .IN3(n797), .IN4(n802), .Q(n798) );
  OA22X1 U957 ( .IN1(n803), .IN2(n802), .IN3(n801), .IN4(n800), .Q(n810) );
  OR3X1 U958 ( .IN1(n806), .IN2(n815), .IN3(n805), .Q(n808) );
  NAND4X0 U959 ( .IN1(n810), .IN2(n809), .IN3(n808), .IN4(n807), .QN(n832) );
  AO222X1 U960 ( .IN1(n813), .IN2(n812), .IN3(n811), .IN4(n814), .IN5(n815), 
        .IN6(pre_sig_res_03[10]), .Q(n831) );
  AO22X1 U961 ( .IN1(pre_sig_res_03[9]), .IN2(n815), .IN3(n814), .IN4(n813), 
        .Q(n830) );
  AO222X1 U962 ( .IN1(input_factor_02[23]), .IN2(n819), .IN3(
        input_factor_01[23]), .IN4(n818), .IN5(larger_exponent[0]), .IN6(n844), 
        .Q(n829) );
  AO222X1 U963 ( .IN1(input_factor_02[24]), .IN2(n819), .IN3(
        input_factor_01[24]), .IN4(n818), .IN5(n844), .IN6(larger_exponent[1]), 
        .Q(n828) );
  AO222X1 U964 ( .IN1(input_factor_02[25]), .IN2(n819), .IN3(
        input_factor_01[25]), .IN4(n818), .IN5(n844), .IN6(larger_exponent[2]), 
        .Q(n827) );
  AO222X1 U965 ( .IN1(input_factor_02[26]), .IN2(n819), .IN3(
        input_factor_01[26]), .IN4(n818), .IN5(n844), .IN6(larger_exponent[3]), 
        .Q(n826) );
  AO222X1 U966 ( .IN1(input_factor_02[27]), .IN2(n819), .IN3(
        input_factor_01[27]), .IN4(n818), .IN5(n844), .IN6(larger_exponent[4]), 
        .Q(n825) );
  AO222X1 U967 ( .IN1(input_factor_02[28]), .IN2(n819), .IN3(
        input_factor_01[28]), .IN4(n818), .IN5(n844), .IN6(larger_exponent[5]), 
        .Q(n824) );
  AO222X1 U968 ( .IN1(input_factor_02[29]), .IN2(n819), .IN3(
        input_factor_01[29]), .IN4(n818), .IN5(n844), .IN6(larger_exponent[6]), 
        .Q(n823) );
endmodule


module add_593 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_594 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_595 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_596 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_597 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_598 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_599 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_600 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_601 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_602 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_603 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_604 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_605 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_606 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_607 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_608 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_609 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_610 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_611 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_612 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_613 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_614 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_615 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_616 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(b), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(b), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module adder24_11 ( clk, rst_n, a, b, cin, out );
  input [23:0] a;
  input [23:0] b;
  output [24:0] out;
  input clk, rst_n, cin;
  wire   c_tmp;
  wire   [24:0] s;
  wire   [22:0] c;

  add_616 add_01 ( .s(s[0]), .a(a[0]), .b(b[0]), .ci(1'b0), .co(c[0]) );
  add_615 add_02 ( .s(s[1]), .a(a[1]), .b(b[1]), .ci(c[0]), .co(c[1]) );
  add_614 add_03 ( .s(s[2]), .a(a[2]), .b(b[2]), .ci(c[1]), .co(c[2]) );
  add_613 add_04 ( .s(s[3]), .a(a[3]), .b(b[3]), .ci(c[2]), .co(c[3]) );
  add_612 add_05 ( .s(s[4]), .a(a[4]), .b(b[4]), .ci(c[3]), .co(c[4]) );
  add_611 add_06 ( .s(s[5]), .a(a[5]), .b(b[5]), .ci(c[4]), .co(c[5]) );
  add_610 add_07 ( .s(s[6]), .a(a[6]), .b(b[6]), .ci(c[5]), .co(c[6]) );
  add_609 add_08 ( .s(s[7]), .a(a[7]), .b(b[7]), .ci(c[6]), .co(c[7]) );
  add_608 add_09 ( .s(s[8]), .a(a[8]), .b(b[8]), .ci(c[7]), .co(c[8]) );
  add_607 add_10 ( .s(s[9]), .a(a[9]), .b(b[9]), .ci(c[8]), .co(c[9]) );
  add_606 add_11 ( .s(s[10]), .a(a[10]), .b(b[10]), .ci(c[9]), .co(c[10]) );
  add_605 add_12 ( .s(s[11]), .a(a[11]), .b(b[11]), .ci(c_tmp), .co(c[11]) );
  add_604 add_13 ( .s(s[12]), .a(a[12]), .b(b[12]), .ci(c[11]), .co(c[12]) );
  add_603 add_14 ( .s(s[13]), .a(a[13]), .b(b[13]), .ci(c[12]), .co(c[13]) );
  add_602 add_15 ( .s(s[14]), .a(a[14]), .b(b[14]), .ci(c[13]), .co(c[14]) );
  add_601 add_16 ( .s(s[15]), .a(a[15]), .b(b[15]), .ci(c[14]), .co(c[15]) );
  add_600 add_17 ( .s(s[16]), .a(a[16]), .b(b[16]), .ci(c[15]), .co(c[16]) );
  add_599 add_18 ( .s(s[17]), .a(a[17]), .b(b[17]), .ci(c[16]), .co(c[17]) );
  add_598 add_19 ( .s(s[18]), .a(a[18]), .b(b[18]), .ci(c[17]), .co(c[18]) );
  add_597 add_20 ( .s(s[19]), .a(a[19]), .b(b[19]), .ci(c[18]), .co(c[19]) );
  add_596 add_21 ( .s(s[20]), .a(a[20]), .b(b[20]), .ci(c[19]), .co(c[20]) );
  add_595 add_22 ( .s(s[21]), .a(a[21]), .b(b[21]), .ci(c[20]), .co(c[21]) );
  add_594 add_23 ( .s(s[22]), .a(a[22]), .b(b[22]), .ci(c[21]), .co(c[22]) );
  add_593 add_24 ( .s(s[23]), .a(a[23]), .b(b[23]), .ci(c[22]), .co(s[24]) );
  DFFARX1 out_reg_10_ ( .D(s[10]), .CLK(clk), .RSTB(rst_n), .Q(out[10]) );
  DFFARX1 out_reg_9_ ( .D(s[9]), .CLK(clk), .RSTB(rst_n), .Q(out[9]) );
  DFFARX1 out_reg_8_ ( .D(s[8]), .CLK(clk), .RSTB(rst_n), .Q(out[8]) );
  DFFARX1 out_reg_7_ ( .D(s[7]), .CLK(clk), .RSTB(rst_n), .Q(out[7]) );
  DFFARX1 out_reg_6_ ( .D(s[6]), .CLK(clk), .RSTB(rst_n), .Q(out[6]) );
  DFFARX1 out_reg_5_ ( .D(s[5]), .CLK(clk), .RSTB(rst_n), .Q(out[5]) );
  DFFARX1 out_reg_4_ ( .D(s[4]), .CLK(clk), .RSTB(rst_n), .Q(out[4]) );
  DFFARX1 out_reg_3_ ( .D(s[3]), .CLK(clk), .RSTB(rst_n), .Q(out[3]) );
  DFFARX1 out_reg_2_ ( .D(s[2]), .CLK(clk), .RSTB(rst_n), .Q(out[2]) );
  DFFARX1 out_reg_1_ ( .D(s[1]), .CLK(clk), .RSTB(rst_n), .Q(out[1]) );
  DFFARX1 out_reg_0_ ( .D(s[0]), .CLK(clk), .RSTB(rst_n), .Q(out[0]) );
  DFFARX1 c_tmp_reg ( .D(c[10]), .CLK(clk), .RSTB(rst_n), .Q(c_tmp) );
  DFFARX1 out_reg_24_ ( .D(s[24]), .CLK(clk), .RSTB(rst_n), .Q(out[24]) );
  DFFARX1 out_reg_23_ ( .D(s[23]), .CLK(clk), .RSTB(rst_n), .Q(out[23]) );
  DFFARX1 out_reg_22_ ( .D(s[22]), .CLK(clk), .RSTB(rst_n), .Q(out[22]) );
  DFFARX1 out_reg_21_ ( .D(s[21]), .CLK(clk), .RSTB(rst_n), .Q(out[21]) );
  DFFARX1 out_reg_20_ ( .D(s[20]), .CLK(clk), .RSTB(rst_n), .Q(out[20]) );
  DFFARX1 out_reg_19_ ( .D(s[19]), .CLK(clk), .RSTB(rst_n), .Q(out[19]) );
  DFFARX1 out_reg_18_ ( .D(s[18]), .CLK(clk), .RSTB(rst_n), .Q(out[18]) );
  DFFARX1 out_reg_17_ ( .D(s[17]), .CLK(clk), .RSTB(rst_n), .Q(out[17]) );
  DFFARX1 out_reg_16_ ( .D(s[16]), .CLK(clk), .RSTB(rst_n), .Q(out[16]) );
  DFFARX1 out_reg_15_ ( .D(s[15]), .CLK(clk), .RSTB(rst_n), .Q(out[15]) );
  DFFARX1 out_reg_14_ ( .D(s[14]), .CLK(clk), .RSTB(rst_n), .Q(out[14]) );
  DFFARX1 out_reg_13_ ( .D(s[13]), .CLK(clk), .RSTB(rst_n), .Q(out[13]) );
  DFFARX1 out_reg_12_ ( .D(s[12]), .CLK(clk), .RSTB(rst_n), .Q(out[12]) );
  DFFARX1 out_reg_11_ ( .D(s[11]), .CLK(clk), .RSTB(rst_n), .Q(out[11]) );
endmodule


module add_617 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_618 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_619 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_620 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_621 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_622 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_623 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_624 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_625 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_626 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_627 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_628 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_629 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_630 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_631 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_632 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_633 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_634 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_635 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_636 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_637 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_638 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_639 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_640 ( s, a, ci, co, b_BAR );
  input a, ci, b_BAR;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(b_BAR), .IN2(n1), .QN(co) );
  INVX0 U2 ( .INP(a), .ZN(n1) );
  MUX21X1 U3 ( .IN1(a), .IN2(n1), .S(b_BAR), .Q(s) );
endmodule


module adder24_12 ( clk, rst_n, a, b, cin, out );
  input [23:0] a;
  input [23:0] b;
  output [24:0] out;
  input clk, rst_n, cin;
  wire   c_tmp, n_1_net_, n_2_net_, n_3_net_, n_4_net_, n_5_net_, n_6_net_,
         n_7_net_, n_8_net_, n_9_net_, n_10_net_, n_11_net_, n_12_net_,
         n_13_net_, n_14_net_, n_15_net_, n_16_net_, n_17_net_, n_18_net_,
         n_19_net_, n_20_net_, n_21_net_, n_22_net_, n_23_net_;
  wire   [24:0] s;
  wire   [23:0] c;

  add_640 add_01 ( .s(s[0]), .a(a[0]), .ci(1'b1), .co(c[0]), .b_BAR(b[0]) );
  add_639 add_02 ( .s(s[1]), .a(a[1]), .b(n_1_net_), .ci(c[0]), .co(c[1]) );
  add_638 add_03 ( .s(s[2]), .a(a[2]), .b(n_2_net_), .ci(c[1]), .co(c[2]) );
  add_637 add_04 ( .s(s[3]), .a(a[3]), .b(n_3_net_), .ci(c[2]), .co(c[3]) );
  add_636 add_05 ( .s(s[4]), .a(a[4]), .b(n_4_net_), .ci(c[3]), .co(c[4]) );
  add_635 add_06 ( .s(s[5]), .a(a[5]), .b(n_5_net_), .ci(c[4]), .co(c[5]) );
  add_634 add_07 ( .s(s[6]), .a(a[6]), .b(n_6_net_), .ci(c[5]), .co(c[6]) );
  add_633 add_08 ( .s(s[7]), .a(a[7]), .b(n_7_net_), .ci(c[6]), .co(c[7]) );
  add_632 add_09 ( .s(s[8]), .a(a[8]), .b(n_8_net_), .ci(c[7]), .co(c[8]) );
  add_631 add_10 ( .s(s[9]), .a(a[9]), .b(n_9_net_), .ci(c[8]), .co(c[9]) );
  add_630 add_11 ( .s(s[10]), .a(a[10]), .b(n_10_net_), .ci(c[9]), .co(c[10])
         );
  add_629 add_12 ( .s(s[11]), .a(a[11]), .b(n_11_net_), .ci(c_tmp), .co(c[11])
         );
  add_628 add_13 ( .s(s[12]), .a(a[12]), .b(n_12_net_), .ci(c[11]), .co(c[12])
         );
  add_627 add_14 ( .s(s[13]), .a(a[13]), .b(n_13_net_), .ci(c[12]), .co(c[13])
         );
  add_626 add_15 ( .s(s[14]), .a(a[14]), .b(n_14_net_), .ci(c[13]), .co(c[14])
         );
  add_625 add_16 ( .s(s[15]), .a(a[15]), .b(n_15_net_), .ci(c[14]), .co(c[15])
         );
  add_624 add_17 ( .s(s[16]), .a(a[16]), .b(n_16_net_), .ci(c[15]), .co(c[16])
         );
  add_623 add_18 ( .s(s[17]), .a(a[17]), .b(n_17_net_), .ci(c[16]), .co(c[17])
         );
  add_622 add_19 ( .s(s[18]), .a(a[18]), .b(n_18_net_), .ci(c[17]), .co(c[18])
         );
  add_621 add_20 ( .s(s[19]), .a(a[19]), .b(n_19_net_), .ci(c[18]), .co(c[19])
         );
  add_620 add_21 ( .s(s[20]), .a(a[20]), .b(n_20_net_), .ci(c[19]), .co(c[20])
         );
  add_619 add_22 ( .s(s[21]), .a(a[21]), .b(n_21_net_), .ci(c[20]), .co(c[21])
         );
  add_618 add_23 ( .s(s[22]), .a(a[22]), .b(n_22_net_), .ci(c[21]), .co(c[22])
         );
  add_617 add_24 ( .s(s[23]), .a(a[23]), .b(n_23_net_), .ci(c[22]), .co(c[23])
         );
  DFFARX1 out_reg_10_ ( .D(s[10]), .CLK(clk), .RSTB(rst_n), .Q(out[10]) );
  DFFARX1 out_reg_9_ ( .D(s[9]), .CLK(clk), .RSTB(rst_n), .Q(out[9]) );
  DFFARX1 out_reg_8_ ( .D(s[8]), .CLK(clk), .RSTB(rst_n), .Q(out[8]) );
  DFFARX1 out_reg_7_ ( .D(s[7]), .CLK(clk), .RSTB(rst_n), .Q(out[7]) );
  DFFARX1 out_reg_6_ ( .D(s[6]), .CLK(clk), .RSTB(rst_n), .Q(out[6]) );
  DFFARX1 out_reg_5_ ( .D(s[5]), .CLK(clk), .RSTB(rst_n), .Q(out[5]) );
  DFFARX1 out_reg_4_ ( .D(s[4]), .CLK(clk), .RSTB(rst_n), .Q(out[4]) );
  DFFARX1 out_reg_3_ ( .D(s[3]), .CLK(clk), .RSTB(rst_n), .Q(out[3]) );
  DFFARX1 out_reg_2_ ( .D(s[2]), .CLK(clk), .RSTB(rst_n), .Q(out[2]) );
  DFFARX1 out_reg_1_ ( .D(s[1]), .CLK(clk), .RSTB(rst_n), .Q(out[1]) );
  DFFARX1 out_reg_0_ ( .D(s[0]), .CLK(clk), .RSTB(rst_n), .Q(out[0]) );
  DFFARX1 c_tmp_reg ( .D(c[10]), .CLK(clk), .RSTB(rst_n), .Q(c_tmp) );
  DFFARX1 out_reg_24_ ( .D(s[24]), .CLK(clk), .RSTB(rst_n), .Q(out[24]) );
  DFFARX1 out_reg_23_ ( .D(s[23]), .CLK(clk), .RSTB(rst_n), .Q(out[23]) );
  DFFARX1 out_reg_22_ ( .D(s[22]), .CLK(clk), .RSTB(rst_n), .Q(out[22]) );
  DFFARX1 out_reg_21_ ( .D(s[21]), .CLK(clk), .RSTB(rst_n), .Q(out[21]) );
  DFFARX1 out_reg_20_ ( .D(s[20]), .CLK(clk), .RSTB(rst_n), .Q(out[20]) );
  DFFARX1 out_reg_19_ ( .D(s[19]), .CLK(clk), .RSTB(rst_n), .Q(out[19]) );
  DFFARX1 out_reg_18_ ( .D(s[18]), .CLK(clk), .RSTB(rst_n), .Q(out[18]) );
  DFFARX1 out_reg_17_ ( .D(s[17]), .CLK(clk), .RSTB(rst_n), .Q(out[17]) );
  DFFARX1 out_reg_16_ ( .D(s[16]), .CLK(clk), .RSTB(rst_n), .Q(out[16]) );
  DFFARX1 out_reg_15_ ( .D(s[15]), .CLK(clk), .RSTB(rst_n), .Q(out[15]) );
  DFFARX1 out_reg_14_ ( .D(s[14]), .CLK(clk), .RSTB(rst_n), .Q(out[14]) );
  DFFARX1 out_reg_13_ ( .D(s[13]), .CLK(clk), .RSTB(rst_n), .Q(out[13]) );
  DFFARX1 out_reg_12_ ( .D(s[12]), .CLK(clk), .RSTB(rst_n), .Q(out[12]) );
  DFFARX1 out_reg_11_ ( .D(s[11]), .CLK(clk), .RSTB(rst_n), .Q(out[11]) );
  INVX0 U3 ( .INP(b[1]), .ZN(n_1_net_) );
  INVX0 U4 ( .INP(b[2]), .ZN(n_2_net_) );
  INVX0 U5 ( .INP(b[3]), .ZN(n_3_net_) );
  INVX0 U6 ( .INP(b[4]), .ZN(n_4_net_) );
  INVX0 U7 ( .INP(b[5]), .ZN(n_5_net_) );
  INVX0 U8 ( .INP(b[6]), .ZN(n_6_net_) );
  INVX0 U9 ( .INP(b[7]), .ZN(n_7_net_) );
  INVX0 U10 ( .INP(b[8]), .ZN(n_8_net_) );
  INVX0 U11 ( .INP(b[9]), .ZN(n_9_net_) );
  INVX0 U12 ( .INP(b[10]), .ZN(n_10_net_) );
  INVX0 U13 ( .INP(c[23]), .ZN(s[24]) );
  INVX0 U14 ( .INP(b[11]), .ZN(n_11_net_) );
  INVX0 U15 ( .INP(b[12]), .ZN(n_12_net_) );
  INVX0 U16 ( .INP(b[13]), .ZN(n_13_net_) );
  INVX0 U17 ( .INP(b[14]), .ZN(n_14_net_) );
  INVX0 U18 ( .INP(b[15]), .ZN(n_15_net_) );
  INVX0 U19 ( .INP(b[16]), .ZN(n_16_net_) );
  INVX0 U20 ( .INP(b[17]), .ZN(n_17_net_) );
  INVX0 U21 ( .INP(b[18]), .ZN(n_18_net_) );
  INVX0 U22 ( .INP(b[19]), .ZN(n_19_net_) );
  INVX0 U23 ( .INP(b[20]), .ZN(n_20_net_) );
  INVX0 U24 ( .INP(b[21]), .ZN(n_21_net_) );
  INVX0 U25 ( .INP(b[22]), .ZN(n_22_net_) );
  INVX0 U26 ( .INP(b[23]), .ZN(n_23_net_) );
endmodule


module add_561 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  XNOR2X1 U1 ( .IN1(ci), .IN2(a), .Q(s) );
endmodule


module add_562 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_563 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_564 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_565 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_566 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_567 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_568 ( s, a, ci, co, b_BAR );
  input a, ci, b_BAR;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(b_BAR), .IN2(n1), .QN(co) );
  INVX0 U2 ( .INP(a), .ZN(n1) );
  MUX21X1 U3 ( .IN1(a), .IN2(n1), .S(b_BAR), .Q(s) );
endmodule


module adder8_41 ( out, a, b, cin );
  output [7:0] out;
  input [7:0] a;
  input [7:0] b;
  input cin;
  wire   n_1_net_, n_2_net_, n_4_net_;
  wire   [6:0] c;

  add_568 add_01 ( .s(out[0]), .a(a[0]), .ci(1'b1), .co(c[0]), .b_BAR(b[0]) );
  add_567 add_02 ( .s(out[1]), .a(a[1]), .b(n_1_net_), .ci(c[0]), .co(c[1]) );
  add_566 add_03 ( .s(out[2]), .a(a[2]), .b(n_2_net_), .ci(c[1]), .co(c[2]) );
  add_565 add_04 ( .s(out[3]), .a(a[3]), .b(1'b1), .ci(c[2]), .co(c[3]) );
  add_564 add_05 ( .s(out[4]), .a(a[4]), .b(n_4_net_), .ci(c[3]), .co(c[4]) );
  add_563 add_06 ( .s(out[5]), .a(a[5]), .b(1'b1), .ci(c[4]), .co(c[5]) );
  add_562 add_07 ( .s(out[6]), .a(a[6]), .b(1'b1), .ci(c[5]), .co(c[6]) );
  add_561 add_08 ( .s(out[7]), .a(a[7]), .b(1'b1), .ci(c[6]) );
  INVX0 U1 ( .INP(b[1]), .ZN(n_1_net_) );
  INVX0 U2 ( .INP(b[2]), .ZN(n_2_net_) );
  INVX0 U3 ( .INP(b[4]), .ZN(n_4_net_) );
endmodule


module add_569 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  XNOR2X1 U1 ( .IN1(ci), .IN2(a), .Q(s) );
endmodule


module add_570 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_571 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_572 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_573 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_574 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_575 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_576 ( s, a, ci, co, b_BAR );
  input a, ci, b_BAR;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(b_BAR), .IN2(n1), .QN(co) );
  INVX0 U2 ( .INP(a), .ZN(n1) );
  MUX21X1 U3 ( .IN1(a), .IN2(n1), .S(b_BAR), .Q(s) );
endmodule


module adder8_42 ( out, a, b, cin );
  output [7:0] out;
  input [7:0] a;
  input [7:0] b;
  input cin;
  wire   n_1_net_, n_2_net_, n_3_net_;
  wire   [6:0] c;

  add_576 add_01 ( .s(out[0]), .a(a[0]), .ci(1'b1), .co(c[0]), .b_BAR(b[0]) );
  add_575 add_02 ( .s(out[1]), .a(a[1]), .b(n_1_net_), .ci(c[0]), .co(c[1]) );
  add_574 add_03 ( .s(out[2]), .a(a[2]), .b(n_2_net_), .ci(c[1]), .co(c[2]) );
  add_573 add_04 ( .s(out[3]), .a(a[3]), .b(n_3_net_), .ci(c[2]), .co(c[3]) );
  add_572 add_05 ( .s(out[4]), .a(a[4]), .b(1'b1), .ci(c[3]), .co(c[4]) );
  add_571 add_06 ( .s(out[5]), .a(a[5]), .b(1'b1), .ci(c[4]), .co(c[5]) );
  add_570 add_07 ( .s(out[6]), .a(a[6]), .b(1'b1), .ci(c[5]), .co(c[6]) );
  add_569 add_08 ( .s(out[7]), .a(a[7]), .b(1'b1), .ci(c[6]) );
  INVX0 U1 ( .INP(b[1]), .ZN(n_1_net_) );
  INVX0 U2 ( .INP(b[2]), .ZN(n_2_net_) );
  INVX0 U3 ( .INP(b[3]), .ZN(n_3_net_) );
endmodule


module add_577 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  XNOR2X1 U1 ( .IN1(ci), .IN2(a), .Q(s) );
endmodule


module add_578 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_579 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_580 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_581 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_582 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_583 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_584 ( s, a, ci, co, b_BAR );
  input a, ci, b_BAR;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(b_BAR), .IN2(n1), .QN(co) );
  INVX0 U2 ( .INP(a), .ZN(n1) );
  MUX21X1 U3 ( .IN1(a), .IN2(n1), .S(b_BAR), .Q(s) );
endmodule


module adder8_43 ( out, a, b, cin );
  output [7:0] out;
  input [7:0] a;
  input [7:0] b;
  input cin;
  wire   n_1_net_, n_2_net_, n_3_net_;
  wire   [6:0] c;

  add_584 add_01 ( .s(out[0]), .a(a[0]), .ci(1'b1), .co(c[0]), .b_BAR(b[0]) );
  add_583 add_02 ( .s(out[1]), .a(a[1]), .b(n_1_net_), .ci(c[0]), .co(c[1]) );
  add_582 add_03 ( .s(out[2]), .a(a[2]), .b(n_2_net_), .ci(c[1]), .co(c[2]) );
  add_581 add_04 ( .s(out[3]), .a(a[3]), .b(n_3_net_), .ci(c[2]), .co(c[3]) );
  add_580 add_05 ( .s(out[4]), .a(a[4]), .b(1'b1), .ci(c[3]), .co(c[4]) );
  add_579 add_06 ( .s(out[5]), .a(a[5]), .b(1'b1), .ci(c[4]), .co(c[5]) );
  add_578 add_07 ( .s(out[6]), .a(a[6]), .b(1'b1), .ci(c[5]), .co(c[6]) );
  add_577 add_08 ( .s(out[7]), .a(a[7]), .b(1'b1), .ci(c[6]) );
  INVX0 U1 ( .INP(b[1]), .ZN(n_1_net_) );
  INVX0 U2 ( .INP(b[2]), .ZN(n_2_net_) );
  INVX0 U3 ( .INP(b[3]), .ZN(n_3_net_) );
endmodule


module add_585 ( s, a, b, co, ci_BAR );
  input a, b, ci_BAR;
  output s, co;


  XNOR2X1 U1 ( .IN1(a), .IN2(ci_BAR), .Q(s) );
endmodule


module add_586 ( s, a, b, ci, co_BAR );
  input a, b, ci;
  output s, co_BAR;


  NAND2X0 U1 ( .IN1(ci), .IN2(a), .QN(co_BAR) );
  OA21X1 U2 ( .IN1(ci), .IN2(a), .IN3(co_BAR), .Q(s) );
endmodule


module add_587 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_588 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_589 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_590 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_591 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_592 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(b), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(b), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module adder8_44 ( out, a, b, cin );
  output [7:0] out;
  input [7:0] a;
  input [7:0] b;
  input cin;

  wire   [6:0] c;

  add_592 add_01 ( .s(out[0]), .a(a[0]), .b(b[0]), .ci(1'b0), .co(c[0]) );
  add_591 add_02 ( .s(out[1]), .a(a[1]), .b(1'b0), .ci(c[0]), .co(c[1]) );
  add_590 add_03 ( .s(out[2]), .a(a[2]), .b(1'b0), .ci(c[1]), .co(c[2]) );
  add_589 add_04 ( .s(out[3]), .a(a[3]), .b(1'b0), .ci(c[2]), .co(c[3]) );
  add_588 add_05 ( .s(out[4]), .a(a[4]), .b(1'b0), .ci(c[3]), .co(c[4]) );
  add_587 add_06 ( .s(out[5]), .a(a[5]), .b(1'b0), .ci(c[4]), .co(c[5]) );
  add_586 add_07 ( .s(out[6]), .a(a[6]), .b(1'b0), .ci(c[5]), .co_BAR(c[6]) );
  add_585 add_08 ( .s(out[7]), .a(a[7]), .b(1'b0), .ci_BAR(c[6]) );
endmodule


module add_641 ( s, a, ci, co, b_BAR );
  input a, ci, b_BAR;
  output s, co;


  XNOR2X1 U1 ( .IN1(ci), .IN2(a), .Q(s) );
endmodule


module add_642 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_643 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_644 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_645 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_646 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_647 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_648 ( s, a, ci, co, b_BAR );
  input a, ci, b_BAR;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(b_BAR), .IN2(n1), .QN(co) );
  INVX0 U2 ( .INP(a), .ZN(n1) );
  MUX21X1 U3 ( .IN1(a), .IN2(n1), .S(b_BAR), .Q(s) );
endmodule


module adder8_45 ( out, a, b, cin );
  output [7:0] out;
  input [7:0] a;
  input [7:0] b;
  input cin;
  wire   n_1_net_, n_2_net_, n_3_net_, n_4_net_, n_5_net_, n_6_net_;
  wire   [6:0] c;

  add_648 add_01 ( .s(out[0]), .a(a[0]), .ci(1'b1), .co(c[0]), .b_BAR(b[0]) );
  add_647 add_02 ( .s(out[1]), .a(a[1]), .b(n_1_net_), .ci(c[0]), .co(c[1]) );
  add_646 add_03 ( .s(out[2]), .a(a[2]), .b(n_2_net_), .ci(c[1]), .co(c[2]) );
  add_645 add_04 ( .s(out[3]), .a(a[3]), .b(n_3_net_), .ci(c[2]), .co(c[3]) );
  add_644 add_05 ( .s(out[4]), .a(a[4]), .b(n_4_net_), .ci(c[3]), .co(c[4]) );
  add_643 add_06 ( .s(out[5]), .a(a[5]), .b(n_5_net_), .ci(c[4]), .co(c[5]) );
  add_642 add_07 ( .s(out[6]), .a(a[6]), .b(n_6_net_), .ci(c[5]), .co(c[6]) );
  add_641 add_08 ( .s(out[7]), .a(a[7]), .ci(c[6]), .b_BAR(1'b0) );
  INVX0 U1 ( .INP(b[1]), .ZN(n_1_net_) );
  INVX0 U2 ( .INP(b[2]), .ZN(n_2_net_) );
  INVX0 U3 ( .INP(b[3]), .ZN(n_3_net_) );
  INVX0 U4 ( .INP(b[4]), .ZN(n_4_net_) );
  INVX0 U5 ( .INP(b[5]), .ZN(n_5_net_) );
  INVX0 U6 ( .INP(b[6]), .ZN(n_6_net_) );
endmodule


module add_649 ( s, a, ci, co, b_BAR );
  input a, ci, b_BAR;
  output s, co;


  XNOR2X1 U1 ( .IN1(b_BAR), .IN2(ci), .Q(s) );
endmodule


module add_650 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_651 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_652 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_653 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_654 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_655 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_656 ( s, a, ci, co, b_BAR );
  input a, ci, b_BAR;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(b_BAR), .IN2(n1), .QN(co) );
  INVX0 U2 ( .INP(a), .ZN(n1) );
  MUX21X1 U3 ( .IN1(a), .IN2(n1), .S(b_BAR), .Q(s) );
endmodule


module adder8_46 ( out, a, b, cin );
  output [7:0] out;
  input [7:0] a;
  input [7:0] b;
  input cin;
  wire   n_1_net_, n_2_net_, n_3_net_, n_4_net_, n_5_net_, n_6_net_;
  wire   [6:0] c;

  add_656 add_01 ( .s(out[0]), .a(a[0]), .ci(1'b1), .co(c[0]), .b_BAR(b[0]) );
  add_655 add_02 ( .s(out[1]), .a(a[1]), .b(n_1_net_), .ci(c[0]), .co(c[1]) );
  add_654 add_03 ( .s(out[2]), .a(a[2]), .b(n_2_net_), .ci(c[1]), .co(c[2]) );
  add_653 add_04 ( .s(out[3]), .a(a[3]), .b(n_3_net_), .ci(c[2]), .co(c[3]) );
  add_652 add_05 ( .s(out[4]), .a(a[4]), .b(n_4_net_), .ci(c[3]), .co(c[4]) );
  add_651 add_06 ( .s(out[5]), .a(a[5]), .b(n_5_net_), .ci(c[4]), .co(c[5]) );
  add_650 add_07 ( .s(out[6]), .a(a[6]), .b(n_6_net_), .ci(c[5]), .co(c[6]) );
  add_649 add_08 ( .s(out[7]), .a(1'b0), .ci(c[6]), .b_BAR(b[7]) );
  INVX0 U1 ( .INP(b[1]), .ZN(n_1_net_) );
  INVX0 U2 ( .INP(b[2]), .ZN(n_2_net_) );
  INVX0 U3 ( .INP(b[3]), .ZN(n_3_net_) );
  INVX0 U4 ( .INP(b[4]), .ZN(n_4_net_) );
  INVX0 U5 ( .INP(b[5]), .ZN(n_5_net_) );
  INVX0 U6 ( .INP(b[6]), .ZN(n_6_net_) );
endmodule


module floating_point_adder_6 ( clk, rst_n, input_factor_01, input_factor_02, 
        output_adder );
  input [31:0] input_factor_01;
  input [31:0] input_factor_02;
  output [31:0] output_adder;
  input clk, rst_n;
  wire   N34, N35, N36, N37, N38, N39, N40, N41, N152, N153, N154, N155, N156,
         N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, N167,
         N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178,
         N179, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189,
         N190, N191, N192, N193, N194, N195, N196, N197, N198,
         add_sub_result_24_, N211, shift_temp_01_0_, N226, N227, N228, N229,
         N230, N231, N232, N233, N234, N235, N236, N237, N238, N239, N240,
         N241, N242, N243, N244, N245, N246, N247, N248, N256, N257, N258,
         N260, N261, N262, N263, N264, N265, N266, N267, N268, N269, N270,
         N271, N272, N273, N274, N275, N276, N277, N278, N279, N280, N281,
         N306, N307, N308, N346, N347, N348, N349, N350, N351, N352, N353,
         N354, N355, N380, N381, N382, N383, N384, N385, N386, N387, N388,
         N389, N390, N391, N392, N393, N394, N395, N396, N397, N398, N399,
         N400, N401, N402, N403, N404, N405, N406, N407, N408, N409, N410, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848;
  wire   [7:0] exp_diff_value;
  wire   [7:0] exponent_factor_21;
  wire   [7:0] exponent_factor_12;
  wire   [23:0] shift_smaller_factor;
  wire   [22:0] larger_factor;
  wire   [7:0] larger_exponent;
  wire   [24:0] add_result;
  wire   [24:0] sub_result;
  wire   [22:0] pre_sig_res_01;
  wire   [3:0] shift_temp_02;
  wire   [22:1] pre_sig_res_02;
  wire   [2:0] shift_temp_03;
  wire   [22:9] pre_sig_res_03;
  wire   [4:0] shift_temp_04;
  wire   [22:16] pre_sig_res_04;
  wire   [7:0] add_output_exponent_w1;
  wire   [7:0] add_output_exponent_w2;
  wire   [7:0] add_output_exponent_w3;
  wire   [7:0] add_output_exponent_w4;

  adder8_46 adder8_01 ( .out(exponent_factor_21), .a({1'b0, 
        input_factor_02[29:23]}), .b(input_factor_01[30:23]), .cin(1'b1) );
  adder8_45 adder8_02 ( .out(exponent_factor_12), .a(input_factor_01[30:23]), 
        .b({1'b0, input_factor_02[29:23]}), .cin(1'b1) );
  adder24_12 adder24_01 ( .clk(clk), .rst_n(rst_n), .a({shift_temp_04[4], 
        larger_factor}), .b(shift_smaller_factor), .cin(1'b1), .out(sub_result) );
  adder24_11 adder24_02 ( .clk(clk), .rst_n(rst_n), .a({shift_temp_04[4], 
        larger_factor}), .b(shift_smaller_factor), .cin(1'b0), .out(add_result) );
  adder8_44 adder8_03 ( .out(add_output_exponent_w1), .a(larger_exponent), .b(
        {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, shift_temp_01_0_}), .cin(
        1'b0) );
  adder8_43 adder8_04 ( .out(add_output_exponent_w2), .a(larger_exponent), .b(
        {1'b0, 1'b0, 1'b0, 1'b0, shift_temp_02}), .cin(1'b1) );
  adder8_42 adder8_05 ( .out(add_output_exponent_w3), .a(larger_exponent), .b(
        {1'b0, 1'b0, 1'b0, 1'b0, shift_temp_04[4], shift_temp_03}), .cin(1'b1)
         );
  adder8_41 adder8_06 ( .out(add_output_exponent_w4), .a(larger_exponent), .b(
        {1'b0, 1'b0, 1'b0, shift_temp_04[4], 1'b0, shift_temp_04[2:0]}), .cin(
        1'b1) );
  DFFARX1 exp_diff_value_reg_7_ ( .D(N41), .CLK(clk), .RSTB(rst_n), .Q(
        exp_diff_value[7]) );
  DFFARX1 exp_diff_value_reg_6_ ( .D(N40), .CLK(clk), .RSTB(rst_n), .Q(
        exp_diff_value[6]) );
  DFFARX1 exp_diff_value_reg_5_ ( .D(N39), .CLK(clk), .RSTB(rst_n), .Q(
        exp_diff_value[5]) );
  DFFARX1 exp_diff_value_reg_4_ ( .D(N38), .CLK(clk), .RSTB(rst_n), .Q(
        exp_diff_value[4]) );
  DFFARX1 exp_diff_value_reg_3_ ( .D(N37), .CLK(clk), .RSTB(rst_n), .Q(
        exp_diff_value[3]), .QN(n4) );
  DFFARX1 exp_diff_value_reg_2_ ( .D(N36), .CLK(clk), .RSTB(rst_n), .Q(n2), 
        .QN(n5) );
  DFFARX1 exp_diff_value_reg_1_ ( .D(N35), .CLK(clk), .RSTB(rst_n), .Q(
        exp_diff_value[1]), .QN(n3) );
  DFFARX1 exp_diff_value_reg_0_ ( .D(N34), .CLK(clk), .RSTB(rst_n), .Q(
        exp_diff_value[0]), .QN(n1) );
  DFFARX1 larger_factor_reg_22_ ( .D(N198), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[22]) );
  DFFARX1 larger_factor_reg_21_ ( .D(N197), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[21]) );
  DFFARX1 larger_factor_reg_20_ ( .D(N196), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[20]) );
  DFFARX1 larger_factor_reg_19_ ( .D(N195), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[19]) );
  DFFARX1 larger_factor_reg_18_ ( .D(N194), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[18]) );
  DFFARX1 larger_factor_reg_17_ ( .D(N193), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[17]) );
  DFFARX1 larger_factor_reg_16_ ( .D(N192), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[16]) );
  DFFARX1 larger_factor_reg_15_ ( .D(N191), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[15]) );
  DFFARX1 larger_factor_reg_14_ ( .D(N190), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[14]) );
  DFFARX1 larger_factor_reg_13_ ( .D(N189), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[13]) );
  DFFARX1 larger_factor_reg_12_ ( .D(N188), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[12]) );
  DFFARX1 larger_factor_reg_11_ ( .D(N187), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[11]) );
  DFFARX1 larger_factor_reg_10_ ( .D(N186), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[10]) );
  DFFARX1 larger_factor_reg_9_ ( .D(N185), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[9]) );
  DFFARX1 larger_factor_reg_8_ ( .D(N184), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[8]) );
  DFFARX1 larger_factor_reg_7_ ( .D(N183), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[7]) );
  DFFARX1 larger_factor_reg_6_ ( .D(N182), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[6]) );
  DFFARX1 larger_factor_reg_5_ ( .D(N181), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[5]) );
  DFFARX1 larger_factor_reg_4_ ( .D(N180), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[4]) );
  DFFARX1 larger_factor_reg_3_ ( .D(N179), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[3]) );
  DFFARX1 larger_factor_reg_2_ ( .D(N178), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[2]) );
  DFFARX1 larger_factor_reg_1_ ( .D(N177), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[1]) );
  DFFARX1 larger_factor_reg_0_ ( .D(N176), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[0]) );
  DFFARX1 shift_smaller_factor_reg_23_ ( .D(N175), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[23]) );
  DFFARX1 shift_smaller_factor_reg_22_ ( .D(N174), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[22]) );
  DFFARX1 shift_smaller_factor_reg_21_ ( .D(N173), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[21]) );
  DFFARX1 shift_smaller_factor_reg_20_ ( .D(N172), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[20]) );
  DFFARX1 shift_smaller_factor_reg_19_ ( .D(N171), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[19]) );
  DFFARX1 shift_smaller_factor_reg_18_ ( .D(N170), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[18]) );
  DFFARX1 shift_smaller_factor_reg_17_ ( .D(N169), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[17]) );
  DFFARX1 shift_smaller_factor_reg_16_ ( .D(N168), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[16]) );
  DFFARX1 shift_smaller_factor_reg_15_ ( .D(N167), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[15]) );
  DFFARX1 shift_smaller_factor_reg_14_ ( .D(N166), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[14]) );
  DFFARX1 shift_smaller_factor_reg_13_ ( .D(N165), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[13]) );
  DFFARX1 shift_smaller_factor_reg_12_ ( .D(N164), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[12]) );
  DFFARX1 shift_smaller_factor_reg_11_ ( .D(N163), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[11]) );
  DFFARX1 shift_smaller_factor_reg_10_ ( .D(N162), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[10]) );
  DFFARX1 shift_smaller_factor_reg_9_ ( .D(N161), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[9]) );
  DFFARX1 shift_smaller_factor_reg_8_ ( .D(N160), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[8]) );
  DFFARX1 shift_smaller_factor_reg_7_ ( .D(N159), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[7]) );
  DFFARX1 shift_smaller_factor_reg_6_ ( .D(N158), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[6]) );
  DFFARX1 shift_smaller_factor_reg_5_ ( .D(N157), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[5]) );
  DFFARX1 shift_smaller_factor_reg_4_ ( .D(N156), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[4]) );
  DFFARX1 shift_smaller_factor_reg_3_ ( .D(N155), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[3]) );
  DFFARX1 shift_smaller_factor_reg_2_ ( .D(N154), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[2]) );
  DFFARX1 shift_smaller_factor_reg_1_ ( .D(N153), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[1]) );
  DFFARX1 shift_smaller_factor_reg_0_ ( .D(N152), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[0]) );
  DFFX1 larger_exponent_reg_7_ ( .D(n826), .CLK(clk), .Q(larger_exponent[7])
         );
  DFFX1 larger_exponent_reg_6_ ( .D(n827), .CLK(clk), .Q(larger_exponent[6])
         );
  DFFX1 larger_exponent_reg_5_ ( .D(n828), .CLK(clk), .Q(larger_exponent[5])
         );
  DFFX1 larger_exponent_reg_4_ ( .D(n829), .CLK(clk), .Q(larger_exponent[4])
         );
  DFFX1 larger_exponent_reg_3_ ( .D(n830), .CLK(clk), .Q(larger_exponent[3])
         );
  DFFX1 larger_exponent_reg_2_ ( .D(n831), .CLK(clk), .Q(larger_exponent[2])
         );
  DFFX1 larger_exponent_reg_1_ ( .D(n832), .CLK(clk), .Q(larger_exponent[1])
         );
  DFFX1 larger_exponent_reg_0_ ( .D(n833), .CLK(clk), .Q(larger_exponent[0])
         );
  DFFARX1 shift_temp_04_reg_4_ ( .D(1'b1), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_04[4]) );
  DFFARX1 shift_temp_01_reg_0_ ( .D(add_sub_result_24_), .CLK(clk), .RSTB(
        rst_n), .Q(shift_temp_01_0_) );
  DFFARX1 pre_sig_res_02_reg_1_ ( .D(N260), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[1]) );
  DFFARX1 pre_sig_res_02_reg_2_ ( .D(N261), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[2]) );
  DFFARX1 pre_sig_res_02_reg_3_ ( .D(N262), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[3]) );
  DFFARX1 pre_sig_res_02_reg_4_ ( .D(N263), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[4]) );
  DFFARX1 pre_sig_res_02_reg_5_ ( .D(N264), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[5]) );
  DFFARX1 pre_sig_res_02_reg_6_ ( .D(N265), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[6]) );
  DFFARX1 pre_sig_res_02_reg_7_ ( .D(N266), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[7]) );
  DFFARX1 shift_temp_02_reg_2_ ( .D(N258), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_02[2]) );
  DFFASX1 shift_temp_02_reg_3_ ( .D(n825), .CLK(clk), .SETB(rst_n), .QN(
        shift_temp_02[3]) );
  DFFARX1 pre_sig_res_02_reg_8_ ( .D(N267), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[8]) );
  DFFARX1 pre_sig_res_02_reg_9_ ( .D(N268), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[9]) );
  DFFARX1 pre_sig_res_02_reg_10_ ( .D(N269), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[10]) );
  DFFARX1 pre_sig_res_02_reg_11_ ( .D(N270), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[11]) );
  DFFARX1 pre_sig_res_02_reg_12_ ( .D(N271), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[12]) );
  DFFARX1 pre_sig_res_02_reg_13_ ( .D(N272), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[13]) );
  DFFARX1 pre_sig_res_02_reg_14_ ( .D(N273), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[14]) );
  DFFARX1 pre_sig_res_02_reg_15_ ( .D(N274), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[15]) );
  DFFARX1 pre_sig_res_02_reg_16_ ( .D(N275), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[16]) );
  DFFARX1 pre_sig_res_02_reg_17_ ( .D(N276), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[17]) );
  DFFARX1 pre_sig_res_02_reg_18_ ( .D(N277), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[18]) );
  DFFARX1 pre_sig_res_02_reg_19_ ( .D(N278), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[19]) );
  DFFARX1 pre_sig_res_02_reg_20_ ( .D(N279), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[20]) );
  DFFARX1 pre_sig_res_02_reg_21_ ( .D(N280), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[21]) );
  DFFARX1 pre_sig_res_02_reg_22_ ( .D(N281), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[22]) );
  DFFARX1 shift_temp_02_reg_1_ ( .D(N257), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_02[1]) );
  DFFARX1 shift_temp_02_reg_0_ ( .D(N256), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_02[0]) );
  DFFX1 pre_sig_res_03_reg_9_ ( .D(n834), .CLK(clk), .Q(pre_sig_res_03[9]) );
  DFFX1 pre_sig_res_03_reg_10_ ( .D(n835), .CLK(clk), .Q(pre_sig_res_03[10])
         );
  DFFX1 pre_sig_res_03_reg_12_ ( .D(n836), .CLK(clk), .Q(pre_sig_res_03[12])
         );
  DFFX1 pre_sig_res_03_reg_11_ ( .D(n837), .CLK(clk), .Q(pre_sig_res_03[11])
         );
  DFFX1 pre_sig_res_03_reg_13_ ( .D(n838), .CLK(clk), .Q(pre_sig_res_03[13])
         );
  DFFX1 pre_sig_res_03_reg_14_ ( .D(n839), .CLK(clk), .Q(pre_sig_res_03[14])
         );
  DFFARX1 shift_temp_03_reg_2_ ( .D(N308), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_03[2]) );
  DFFARX1 shift_temp_03_reg_0_ ( .D(N306), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_03[0]) );
  DFFARX1 shift_temp_03_reg_1_ ( .D(N307), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_03[1]) );
  DFFX1 pre_sig_res_03_reg_15_ ( .D(n840), .CLK(clk), .Q(pre_sig_res_03[15])
         );
  DFFX1 pre_sig_res_03_reg_16_ ( .D(n841), .CLK(clk), .Q(pre_sig_res_03[16])
         );
  DFFX1 pre_sig_res_03_reg_17_ ( .D(n842), .CLK(clk), .Q(pre_sig_res_03[17])
         );
  DFFX1 pre_sig_res_03_reg_18_ ( .D(n843), .CLK(clk), .Q(pre_sig_res_03[18])
         );
  DFFX1 pre_sig_res_03_reg_19_ ( .D(n844), .CLK(clk), .Q(pre_sig_res_03[19])
         );
  DFFX1 pre_sig_res_03_reg_20_ ( .D(n845), .CLK(clk), .Q(pre_sig_res_03[20])
         );
  DFFX1 pre_sig_res_03_reg_21_ ( .D(n846), .CLK(clk), .Q(pre_sig_res_03[21])
         );
  DFFX1 pre_sig_res_03_reg_22_ ( .D(n847), .CLK(clk), .Q(pre_sig_res_03[22])
         );
  DFFARX1 pre_sig_res_04_reg_16_ ( .D(N349), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_04[16]) );
  DFFARX1 pre_sig_res_04_reg_17_ ( .D(N350), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_04[17]) );
  DFFARX1 pre_sig_res_04_reg_18_ ( .D(N351), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_04[18]) );
  DFFARX1 pre_sig_res_04_reg_19_ ( .D(N352), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_04[19]) );
  DFFARX1 pre_sig_res_04_reg_20_ ( .D(N353), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_04[20]) );
  DFFARX1 pre_sig_res_04_reg_21_ ( .D(N354), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_04[21]) );
  DFFARX1 pre_sig_res_04_reg_22_ ( .D(N355), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_04[22]) );
  DFFARX1 add_output_sign_reg ( .D(N211), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[31]) );
  DFFARX1 pre_sig_res_01_reg_0_ ( .D(N226), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[0]) );
  DFFARX1 pre_sig_res_01_reg_1_ ( .D(N227), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[1]) );
  DFFARX1 pre_sig_res_01_reg_2_ ( .D(N228), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[2]) );
  DFFARX1 pre_sig_res_01_reg_3_ ( .D(N229), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[3]) );
  DFFARX1 pre_sig_res_01_reg_4_ ( .D(N230), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[4]) );
  DFFARX1 pre_sig_res_01_reg_5_ ( .D(N231), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[5]) );
  DFFARX1 pre_sig_res_01_reg_6_ ( .D(N232), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[6]) );
  DFFARX1 pre_sig_res_01_reg_7_ ( .D(N233), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[7]) );
  DFFARX1 pre_sig_res_01_reg_8_ ( .D(N234), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[8]) );
  DFFARX1 pre_sig_res_01_reg_9_ ( .D(N235), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[9]) );
  DFFARX1 pre_sig_res_01_reg_10_ ( .D(N236), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[10]) );
  DFFARX1 pre_sig_res_01_reg_11_ ( .D(N237), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[11]) );
  DFFARX1 pre_sig_res_01_reg_12_ ( .D(N238), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[12]) );
  DFFARX1 pre_sig_res_01_reg_13_ ( .D(N239), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[13]) );
  DFFARX1 pre_sig_res_01_reg_14_ ( .D(N240), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[14]) );
  DFFARX1 pre_sig_res_01_reg_15_ ( .D(N241), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[15]) );
  DFFARX1 pre_sig_res_01_reg_16_ ( .D(N242), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[16]) );
  DFFARX1 pre_sig_res_01_reg_17_ ( .D(N243), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[17]) );
  DFFARX1 pre_sig_res_01_reg_18_ ( .D(N244), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[18]) );
  DFFARX1 pre_sig_res_01_reg_19_ ( .D(N245), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[19]) );
  DFFARX1 pre_sig_res_01_reg_20_ ( .D(N246), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[20]) );
  DFFARX1 pre_sig_res_01_reg_21_ ( .D(N247), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[21]) );
  DFFARX1 pre_sig_res_01_reg_22_ ( .D(N248), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[22]) );
  DFFARX1 shift_temp_04_reg_2_ ( .D(N348), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_04[2]) );
  DFFARX1 shift_temp_04_reg_1_ ( .D(N347), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_04[1]) );
  DFFARX1 shift_temp_04_reg_0_ ( .D(N346), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_04[0]) );
  DFFARX1 add_output_exponent_reg_7_ ( .D(N387), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[30]) );
  DFFARX1 add_output_exponent_reg_6_ ( .D(N386), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[29]) );
  DFFARX1 add_output_exponent_reg_5_ ( .D(N385), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[28]) );
  DFFARX1 add_output_exponent_reg_4_ ( .D(N384), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[27]) );
  DFFARX1 add_output_exponent_reg_3_ ( .D(N383), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[26]) );
  DFFARX1 add_output_exponent_reg_2_ ( .D(N382), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[25]) );
  DFFARX1 add_output_exponent_reg_1_ ( .D(N381), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[24]) );
  DFFARX1 add_output_exponent_reg_0_ ( .D(N380), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[23]) );
  DFFARX1 add_output_significands_reg_22_ ( .D(N410), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[22]) );
  DFFARX1 add_output_significands_reg_21_ ( .D(N409), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[21]) );
  DFFARX1 add_output_significands_reg_20_ ( .D(N408), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[20]) );
  DFFARX1 add_output_significands_reg_19_ ( .D(N407), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[19]) );
  DFFARX1 add_output_significands_reg_18_ ( .D(N406), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[18]) );
  DFFARX1 add_output_significands_reg_17_ ( .D(N405), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[17]) );
  DFFARX1 add_output_significands_reg_16_ ( .D(N404), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[16]) );
  DFFARX1 add_output_significands_reg_15_ ( .D(N403), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[15]) );
  DFFARX1 add_output_significands_reg_14_ ( .D(N402), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[14]) );
  DFFARX1 add_output_significands_reg_13_ ( .D(N401), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[13]) );
  DFFARX1 add_output_significands_reg_12_ ( .D(N400), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[12]) );
  DFFARX1 add_output_significands_reg_11_ ( .D(N399), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[11]) );
  DFFARX1 add_output_significands_reg_10_ ( .D(N398), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[10]) );
  DFFARX1 add_output_significands_reg_9_ ( .D(N397), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[9]) );
  DFFARX1 add_output_significands_reg_8_ ( .D(N396), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[8]) );
  DFFARX1 add_output_significands_reg_7_ ( .D(N395), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[7]) );
  DFFARX1 add_output_significands_reg_6_ ( .D(N394), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[6]) );
  DFFARX1 add_output_significands_reg_5_ ( .D(N393), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[5]) );
  DFFARX1 add_output_significands_reg_4_ ( .D(N392), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[4]) );
  DFFARX1 add_output_significands_reg_3_ ( .D(N391), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[3]) );
  DFFARX1 add_output_significands_reg_2_ ( .D(N390), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[2]) );
  DFFARX1 add_output_significands_reg_1_ ( .D(N389), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[1]) );
  DFFARX1 add_output_significands_reg_0_ ( .D(N388), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[0]) );
  INVX1 U5 ( .INP(rst_n), .ZN(n848) );
  NAND2X0 U3 ( .IN1(n484), .IN2(n397), .QN(n559) );
  NAND2X0 U4 ( .IN1(exp_diff_value[4]), .IN2(n118), .QN(n212) );
  NAND2X0 U6 ( .IN1(input_factor_01[16]), .IN2(n372), .QN(n119) );
  NAND2X0 U7 ( .IN1(input_factor_02[17]), .IN2(n684), .QN(n67) );
  NAND2X0 U8 ( .IN1(n352), .IN2(n356), .QN(n545) );
  NAND2X0 U9 ( .IN1(input_factor_02[24]), .IN2(n543), .QN(n37) );
  NAND2X0 U10 ( .IN1(input_factor_01[27]), .IN2(n585), .QN(n33) );
  NAND2X0 U11 ( .IN1(input_factor_01[26]), .IN2(n579), .QN(n34) );
  NAND2X0 U12 ( .IN1(n23), .IN2(input_factor_02[25]), .QN(n36) );
  NAND2X0 U13 ( .IN1(input_factor_01[28]), .IN2(n591), .QN(n44) );
  NAND2X0 U14 ( .IN1(input_factor_02[28]), .IN2(n590), .QN(n48) );
  NAND2X0 U15 ( .IN1(n806), .IN2(n524), .QN(n382) );
  NAND2X0 U16 ( .IN1(n776), .IN2(n516), .QN(n381) );
  NAND2X0 U17 ( .IN1(n769), .IN2(n517), .QN(n380) );
  NAND2X0 U18 ( .IN1(n745), .IN2(n719), .QN(n556) );
  NAND2X0 U19 ( .IN1(n401), .IN2(n494), .QN(n378) );
  NAND2X0 U20 ( .IN1(n492), .IN2(n404), .QN(n377) );
  NAND2X0 U21 ( .IN1(n376), .IN2(n565), .QN(n403) );
  NAND2X0 U22 ( .IN1(n79), .IN2(n77), .QN(n218) );
  NAND2X0 U23 ( .IN1(n83), .IN2(n82), .QN(n219) );
  NAND2X0 U24 ( .IN1(n129), .IN2(n128), .QN(n240) );
  NAND2X0 U25 ( .IN1(n158), .IN2(n157), .QN(n249) );
  NAND2X0 U26 ( .IN1(n156), .IN2(n155), .QN(n250) );
  NAND2X0 U27 ( .IN1(n183), .IN2(n182), .QN(n269) );
  NAND2X0 U28 ( .IN1(exp_diff_value[1]), .IN2(exp_diff_value[0]), .QN(n184) );
  NAND2X0 U29 ( .IN1(n81), .IN2(n80), .QN(n226) );
  NAND2X0 U30 ( .IN1(n133), .IN2(n132), .QN(n236) );
  NAND2X0 U31 ( .IN1(n160), .IN2(n159), .QN(n257) );
  NAND2X0 U32 ( .IN1(n119), .IN2(n120), .QN(n19) );
  NAND2X0 U33 ( .IN1(input_factor_02[21]), .IN2(n700), .QN(n70) );
  NAND2X0 U34 ( .IN1(input_factor_02[27]), .IN2(n584), .QN(n26) );
  NAND2X0 U35 ( .IN1(input_factor_02[26]), .IN2(n578), .QN(n24) );
  NAND2X0 U36 ( .IN1(input_factor_01[23]), .IN2(n383), .QN(n35) );
  NAND2X0 U37 ( .IN1(n3), .IN2(n1), .QN(n207) );
  NAND2X0 U38 ( .IN1(n373), .IN2(n73), .QN(n72) );
  NAND2X0 U39 ( .IN1(n709), .IN2(pre_sig_res_01[9]), .QN(n640) );
  NAND2X0 U40 ( .IN1(n709), .IN2(pre_sig_res_01[10]), .QN(n646) );
  NAND2X0 U41 ( .IN1(n709), .IN2(pre_sig_res_01[11]), .QN(n652) );
  NAND2X0 U42 ( .IN1(n709), .IN2(pre_sig_res_01[12]), .QN(n658) );
  NAND2X0 U43 ( .IN1(n709), .IN2(pre_sig_res_01[13]), .QN(n664) );
  NAND2X0 U44 ( .IN1(n709), .IN2(pre_sig_res_01[14]), .QN(n670) );
  NAND2X0 U45 ( .IN1(n709), .IN2(pre_sig_res_01[15]), .QN(n676) );
  NAND2X0 U46 ( .IN1(n709), .IN2(pre_sig_res_01[16]), .QN(n680) );
  NAND2X0 U47 ( .IN1(n709), .IN2(pre_sig_res_01[17]), .QN(n686) );
  NAND2X0 U48 ( .IN1(n709), .IN2(pre_sig_res_01[20]), .QN(n696) );
  NAND2X0 U49 ( .IN1(n709), .IN2(pre_sig_res_01[21]), .QN(n704) );
  NAND2X0 U50 ( .IN1(n709), .IN2(add_output_exponent_w1[0]), .QN(n566) );
  NAND2X0 U51 ( .IN1(n709), .IN2(add_output_exponent_w1[1]), .QN(n570) );
  NAND2X0 U52 ( .IN1(n709), .IN2(add_output_exponent_w1[2]), .QN(n574) );
  NAND2X0 U53 ( .IN1(n709), .IN2(add_output_exponent_w1[3]), .QN(n580) );
  NAND2X0 U54 ( .IN1(n709), .IN2(add_output_exponent_w1[4]), .QN(n586) );
  NAND2X0 U55 ( .IN1(n709), .IN2(add_output_exponent_w1[5]), .QN(n592) );
  NAND2X0 U56 ( .IN1(n709), .IN2(add_output_exponent_w1[6]), .QN(n598) );
  NAND2X0 U57 ( .IN1(n518), .IN2(n816), .QN(n536) );
  NAND2X0 U58 ( .IN1(n515), .IN2(n524), .QN(n521) );
  NAND2X0 U59 ( .IN1(n72), .IN2(n367), .QN(n393) );
  NAND2X0 U60 ( .IN1(n516), .IN2(n789), .QN(n534) );
  NAND2X0 U61 ( .IN1(n517), .IN2(n756), .QN(n535) );
  NAND2X0 U62 ( .IN1(n761), .IN2(n745), .QN(n720) );
  NAND2X0 U63 ( .IN1(n719), .IN2(n732), .QN(n794) );
  NAND2X0 U64 ( .IN1(n514), .IN2(n502), .QN(n723) );
  NAND2X0 U65 ( .IN1(n514), .IN2(n506), .QN(n716) );
  NAND2X0 U66 ( .IN1(n397), .IN2(n396), .QN(n496) );
  NAND2X0 U67 ( .IN1(n414), .IN2(n818), .QN(n411) );
  NAND2X0 U68 ( .IN1(n401), .IN2(n398), .QN(n485) );
  NAND2X0 U69 ( .IN1(n404), .IN2(n399), .QN(n489) );
  NAND2X0 U70 ( .IN1(n400), .IN2(n565), .QN(n487) );
  NAND2X0 U71 ( .IN1(n76), .IN2(n75), .QN(n84) );
  NAND2X0 U72 ( .IN1(n135), .IN2(n134), .QN(n136) );
  NAND2X0 U73 ( .IN1(n162), .IN2(n161), .QN(n163) );
  NAND2X0 U74 ( .IN1(n708), .IN2(n370), .QN(n223) );
  NAND2X0 U75 ( .IN1(n370), .IN2(n821), .QN(n199) );
  NAND2X0 U76 ( .IN1(n186), .IN2(n185), .QN(n187) );
  NAND2X0 U77 ( .IN1(n708), .IN2(n122), .QN(n235) );
  NAND2X0 U78 ( .IN1(n821), .IN2(n122), .QN(n208) );
  NAND2X0 U79 ( .IN1(n220), .IN2(n222), .QN(n17) );
  NAND2X0 U80 ( .IN1(n280), .IN2(n240), .QN(n241) );
  NAND2X0 U81 ( .IN1(n131), .IN2(n130), .QN(n244) );
  NAND2X0 U82 ( .IN1(n821), .IN2(n266), .QN(n253) );
  NAND2X0 U83 ( .IN1(n708), .IN2(n266), .QN(n254) );
  NAND2X0 U84 ( .IN1(n271), .IN2(n272), .QN(n15) );
  NAND2X0 U85 ( .IN1(n270), .IN2(n269), .QN(n271) );
  NAND2X0 U86 ( .IN1(n181), .IN2(n180), .QN(n279) );
  NAND2X0 U87 ( .IN1(exp_diff_value[3]), .IN2(n216), .QN(n336) );
  NAND2X0 U88 ( .IN1(exp_diff_value[1]), .IN2(n1), .QN(n310) );
  NAND2X0 U89 ( .IN1(n323), .IN2(n5), .QN(n325) );
  NAND2X0 U90 ( .IN1(n337), .IN2(n336), .QN(n338) );
  NAND2X0 U91 ( .IN1(n4), .IN2(n216), .QN(n354) );
  NAND2X0 U92 ( .IN1(n311), .IN2(n310), .QN(n358) );
  NAND2X0 U93 ( .IN1(n74), .IN2(n123), .QN(n367) );
  NAND2X0 U94 ( .IN1(n371), .IN2(n216), .QN(n364) );
  NAND2X0 U95 ( .IN1(exp_diff_value[0]), .IN2(n3), .QN(n326) );
  NAND2X0 U96 ( .IN1(n607), .IN2(n606), .QN(N389) );
  NAND2X0 U97 ( .IN1(n611), .IN2(n610), .QN(N390) );
  NAND2X0 U98 ( .IN1(n615), .IN2(n614), .QN(N391) );
  NAND2X0 U99 ( .IN1(n619), .IN2(n618), .QN(N392) );
  NAND2X0 U100 ( .IN1(n623), .IN2(n622), .QN(N393) );
  NAND2X0 U101 ( .IN1(n627), .IN2(n626), .QN(N394) );
  NAND2X0 U102 ( .IN1(n631), .IN2(n630), .QN(N395) );
  NAND2X0 U103 ( .IN1(n635), .IN2(n634), .QN(N396) );
  NAND2X0 U104 ( .IN1(n712), .IN2(pre_sig_res_03[9]), .QN(n638) );
  NAND2X0 U105 ( .IN1(n711), .IN2(pre_sig_res_02[9]), .QN(n639) );
  NAND2X0 U106 ( .IN1(n712), .IN2(pre_sig_res_03[10]), .QN(n644) );
  NAND2X0 U107 ( .IN1(n711), .IN2(pre_sig_res_02[10]), .QN(n645) );
  NAND2X0 U108 ( .IN1(n712), .IN2(pre_sig_res_03[11]), .QN(n650) );
  NAND2X0 U109 ( .IN1(n711), .IN2(pre_sig_res_02[11]), .QN(n651) );
  NAND2X0 U110 ( .IN1(n712), .IN2(pre_sig_res_03[12]), .QN(n656) );
  NAND2X0 U111 ( .IN1(n711), .IN2(pre_sig_res_02[12]), .QN(n657) );
  NAND2X0 U112 ( .IN1(n712), .IN2(pre_sig_res_03[13]), .QN(n662) );
  NAND2X0 U113 ( .IN1(n711), .IN2(pre_sig_res_02[13]), .QN(n663) );
  NAND2X0 U114 ( .IN1(n712), .IN2(pre_sig_res_03[14]), .QN(n668) );
  NAND2X0 U115 ( .IN1(n711), .IN2(pre_sig_res_02[14]), .QN(n669) );
  NAND2X0 U116 ( .IN1(n712), .IN2(pre_sig_res_03[15]), .QN(n674) );
  NAND2X0 U117 ( .IN1(n711), .IN2(pre_sig_res_02[15]), .QN(n675) );
  NAND2X0 U118 ( .IN1(n714), .IN2(pre_sig_res_04[16]), .QN(n681) );
  NAND2X0 U119 ( .IN1(n714), .IN2(pre_sig_res_04[17]), .QN(n687) );
  NAND2X0 U120 ( .IN1(n10), .IN2(n11), .QN(N406) );
  NAND2X0 U121 ( .IN1(n714), .IN2(pre_sig_res_04[18]), .QN(n11) );
  NAND2X0 U122 ( .IN1(n8), .IN2(n9), .QN(N407) );
  NAND2X0 U123 ( .IN1(n714), .IN2(pre_sig_res_04[19]), .QN(n9) );
  NAND2X0 U124 ( .IN1(n714), .IN2(pre_sig_res_04[20]), .QN(n697) );
  NAND2X0 U125 ( .IN1(n714), .IN2(pre_sig_res_04[21]), .QN(n705) );
  NAND2X0 U126 ( .IN1(n6), .IN2(n7), .QN(N410) );
  NAND2X0 U127 ( .IN1(n714), .IN2(pre_sig_res_04[22]), .QN(n7) );
  NAND2X0 U128 ( .IN1(n714), .IN2(add_output_exponent_w4[0]), .QN(n567) );
  NAND2X0 U129 ( .IN1(n714), .IN2(add_output_exponent_w4[1]), .QN(n571) );
  NAND2X0 U130 ( .IN1(n714), .IN2(add_output_exponent_w4[2]), .QN(n575) );
  NAND2X0 U131 ( .IN1(n714), .IN2(add_output_exponent_w4[3]), .QN(n581) );
  NAND2X0 U132 ( .IN1(n714), .IN2(add_output_exponent_w4[4]), .QN(n587) );
  NAND2X0 U133 ( .IN1(n714), .IN2(add_output_exponent_w4[5]), .QN(n593) );
  NAND2X0 U134 ( .IN1(n714), .IN2(add_output_exponent_w4[6]), .QN(n599) );
  NAND2X0 U135 ( .IN1(n12), .IN2(n13), .QN(N387) );
  NAND2X0 U136 ( .IN1(n714), .IN2(add_output_exponent_w4[7]), .QN(n13) );
  NAND2X0 U137 ( .IN1(n521), .IN2(n520), .QN(N348) );
  NAND2X0 U138 ( .IN1(n538), .IN2(n796), .QN(n539) );
  NAND2X0 U139 ( .IN1(n538), .IN2(n816), .QN(n529) );
  NAND2X0 U140 ( .IN1(n538), .IN2(n818), .QN(n525) );
  NAND2X0 U141 ( .IN1(n523), .IN2(n522), .QN(N352) );
  NAND2X0 U142 ( .IN1(pre_sig_res_03[22]), .IN2(n820), .QN(n725) );
  NAND2X0 U143 ( .IN1(n809), .IN2(n724), .QN(n726) );
  NAND2X0 U144 ( .IN1(pre_sig_res_03[21]), .IN2(n820), .QN(n733) );
  NAND2X0 U145 ( .IN1(n809), .IN2(n732), .QN(n734) );
  NAND2X0 U146 ( .IN1(pre_sig_res_03[20]), .IN2(n820), .QN(n741) );
  NAND2X0 U147 ( .IN1(n809), .IN2(n740), .QN(n742) );
  NAND2X0 U148 ( .IN1(pre_sig_res_03[19]), .IN2(n820), .QN(n749) );
  NAND2X0 U149 ( .IN1(n809), .IN2(n748), .QN(n750) );
  NAND2X0 U150 ( .IN1(pre_sig_res_03[18]), .IN2(n820), .QN(n757) );
  NAND2X0 U151 ( .IN1(n809), .IN2(n756), .QN(n758) );
  NAND2X0 U152 ( .IN1(pre_sig_res_03[17]), .IN2(n820), .QN(n765) );
  NAND2X0 U153 ( .IN1(n809), .IN2(n764), .QN(n766) );
  NAND2X0 U154 ( .IN1(pre_sig_res_03[16]), .IN2(n820), .QN(n772) );
  NAND2X0 U155 ( .IN1(n809), .IN2(n789), .QN(n773) );
  NAND2X0 U156 ( .IN1(pre_sig_res_03[15]), .IN2(n820), .QN(n781) );
  NAND2X0 U157 ( .IN1(n809), .IN2(n797), .QN(n782) );
  NAND2X0 U158 ( .IN1(n716), .IN2(n723), .QN(n507) );
  NAND2X0 U159 ( .IN1(pre_sig_res_03[14]), .IN2(n848), .QN(n791) );
  NAND2X0 U160 ( .IN1(n819), .IN2(n789), .QN(n790) );
  NAND2X0 U161 ( .IN1(n809), .IN2(n788), .QN(n792) );
  NAND2X0 U162 ( .IN1(pre_sig_res_03[13]), .IN2(n820), .QN(n799) );
  NAND2X0 U163 ( .IN1(n819), .IN2(n797), .QN(n798) );
  NAND2X0 U164 ( .IN1(n809), .IN2(n796), .QN(n800) );
  NAND2X0 U165 ( .IN1(n804), .IN2(n803), .QN(n837) );
  NAND2X0 U166 ( .IN1(pre_sig_res_03[12]), .IN2(n820), .QN(n812) );
  NAND2X0 U167 ( .IN1(n809), .IN2(n816), .QN(n814) );
  NAND2X0 U168 ( .IN1(n414), .IN2(n816), .QN(n415) );
  NAND2X0 U169 ( .IN1(n419), .IN2(n797), .QN(n410) );
  NAND2X0 U170 ( .IN1(n420), .IN2(n796), .QN(n407) );
  NAND2X0 U171 ( .IN1(n406), .IN2(n405), .QN(N263) );
  NAND2X0 U172 ( .IN1(n323), .IN2(n312), .QN(n227) );
  NAND2X0 U173 ( .IN1(n270), .IN2(n244), .QN(n245) );
  NAND2X0 U174 ( .IN1(n313), .IN2(n312), .QN(n314) );
  NAND2X0 U175 ( .IN1(n345), .IN2(n344), .QN(N168) );
  NAND2X0 U176 ( .IN1(n349), .IN2(n348), .QN(N169) );
  NAND2X0 U177 ( .IN1(n361), .IN2(n360), .QN(N172) );
  NAND2X0 U178 ( .IN1(n369), .IN2(n368), .QN(N173) );
  NAND2X0 U179 ( .IN1(n374), .IN2(n373), .QN(N175) );
  INVX0 U180 ( .INP(n393), .ZN(n392) );
  INVX0 U181 ( .INP(n558), .ZN(n825) );
  INVX0 U182 ( .INP(n419), .ZN(n491) );
  NOR2X0 U183 ( .IN1(n821), .IN2(n848), .QN(n822) );
  NOR2X0 U184 ( .IN1(n723), .IN2(n820), .QN(n809) );
  INVX0 U185 ( .INP(n817), .ZN(n807) );
  INVX0 U186 ( .INP(n796), .ZN(n808) );
  INVX0 U187 ( .INP(n797), .ZN(n786) );
  INVX0 U188 ( .INP(n764), .ZN(n777) );
  NOR2X0 U189 ( .IN1(n561), .IN2(n564), .QN(n711) );
  NOR2X0 U190 ( .IN1(n562), .IN2(n564), .QN(n712) );
  INVX0 U191 ( .INP(n740), .ZN(n753) );
  INVX0 U192 ( .INP(n456), .ZN(n560) );
  INVX0 U193 ( .INP(n559), .ZN(n514) );
  INVX0 U194 ( .INP(n748), .ZN(n761) );
  NOR2X0 U195 ( .IN1(n565), .IN2(n564), .QN(n709) );
  NAND4X0 U196 ( .IN1(n554), .IN2(n553), .IN3(n552), .IN4(n551), .QN(n702) );
  INVX0 U197 ( .INP(n710), .ZN(n701) );
  INVX0 U198 ( .INP(n310), .ZN(n203) );
  INVX0 U199 ( .INP(n207), .ZN(n372) );
  NOR2X0 U200 ( .IN1(n74), .IN2(n73), .QN(n821) );
  INVX0 U201 ( .INP(n313), .ZN(n362) );
  INVX0 U202 ( .INP(n72), .ZN(n708) );
  INVX0 U203 ( .INP(n398), .ZN(n494) );
  NOR2X0 U204 ( .IN1(add_sub_result_24_), .IN2(n395), .QN(n565) );
  MUX21X1 U205 ( .IN1(add_result[24]), .IN2(sub_result[24]), .S(n20), .Q(
        add_sub_result_24_) );
  INVX0 U206 ( .INP(n396), .ZN(n484) );
  INVX0 U207 ( .INP(n21), .ZN(n20) );
  INVX0 U208 ( .INP(n503), .ZN(n21) );
  INVX0 U209 ( .INP(n732), .ZN(n745) );
  INVX0 U210 ( .INP(n756), .ZN(n769) );
  INVX0 U211 ( .INP(n789), .ZN(n776) );
  INVX0 U212 ( .INP(n788), .ZN(n806) );
  INVX0 U213 ( .INP(n816), .ZN(n802) );
  INVX0 U214 ( .INP(n818), .ZN(n810) );
  MUX21X1 U215 ( .IN1(input_factor_01[31]), .IN2(n375), .S(input_factor_02[31]), .Q(n503) );
  NAND2X0 U216 ( .IN1(input_factor_02[29]), .IN2(n596), .QN(n49) );
  INVX0 U217 ( .INP(input_factor_02[29]), .ZN(n597) );
  INVX0 U218 ( .INP(input_factor_01[31]), .ZN(n375) );
  NAND4X0 U219 ( .IN1(n32), .IN2(n31), .IN3(n30), .IN4(n35), .QN(n373) );
  INVX0 U220 ( .INP(n447), .ZN(n718) );
  INVX0 U221 ( .INP(n724), .ZN(n737) );
  INVX0 U222 ( .INP(n442), .ZN(n729) );
  INVX0 U223 ( .INP(n819), .ZN(n805) );
  NOR2X0 U224 ( .IN1(n14), .IN2(n15), .QN(n284) );
  NOR2X0 U225 ( .IN1(n336), .IN2(n334), .QN(n14) );
  NOR2X0 U226 ( .IN1(n693), .IN2(n692), .QN(n8) );
  NOR2X0 U227 ( .IN1(n715), .IN2(n713), .QN(n6) );
  NOR2X0 U228 ( .IN1(n603), .IN2(n602), .QN(n12) );
  NOR2X0 U229 ( .IN1(n691), .IN2(n690), .QN(n10) );
  NAND3X0 U230 ( .IN1(n494), .IN2(n401), .IN3(n465), .QN(n483) );
  OR2X1 U231 ( .IN1(n556), .IN2(n753), .Q(n785) );
  NOR2X0 U232 ( .IN1(n16), .IN2(n17), .QN(n228) );
  NOR2X0 U233 ( .IN1(n364), .IN2(n221), .QN(n16) );
  NOR2X0 U234 ( .IN1(n18), .IN2(n19), .QN(n214) );
  NOR2X0 U235 ( .IN1(n356), .IN2(n184), .QN(n18) );
  INVX0 U236 ( .INP(n184), .ZN(n204) );
  INVX0 U237 ( .INP(n326), .ZN(n202) );
  NOR4X0 U238 ( .IN1(n391), .IN2(n390), .IN3(n389), .IN4(n388), .QN(n710) );
  MUX21X1 U239 ( .IN1(add_result[1]), .IN2(sub_result[1]), .S(n503), .Q(n816)
         );
  INVX0 U240 ( .INP(input_factor_02[12]), .ZN(n655) );
  INVX0 U241 ( .INP(input_factor_02[13]), .ZN(n661) );
  INVX0 U242 ( .INP(input_factor_02[14]), .ZN(n667) );
  INVX0 U243 ( .INP(n702), .ZN(n22) );
  INVX0 U244 ( .INP(input_factor_01[29]), .ZN(n596) );
  INVX0 U245 ( .INP(input_factor_02[23]), .ZN(n383) );
  OA222X1 U246 ( .IN1(input_factor_02[29]), .IN2(n596), .IN3(n597), .IN4(
        input_factor_01[29]), .IN5(input_factor_01[23]), .IN6(n383), .Q(n32)
         );
  INVX0 U247 ( .INP(input_factor_01[25]), .ZN(n23) );
  INVX0 U248 ( .INP(n36), .ZN(n29) );
  NOR2X0 U249 ( .IN1(input_factor_02[25]), .IN2(n23), .QN(n41) );
  INVX0 U250 ( .INP(input_factor_02[28]), .ZN(n591) );
  INVX0 U251 ( .INP(input_factor_02[26]), .ZN(n579) );
  INVX0 U252 ( .INP(input_factor_01[28]), .ZN(n590) );
  INVX0 U253 ( .INP(input_factor_01[26]), .ZN(n578) );
  NAND4X0 U254 ( .IN1(n44), .IN2(n34), .IN3(n48), .IN4(n24), .QN(n28) );
  INVX0 U255 ( .INP(input_factor_01[27]), .ZN(n584) );
  INVX0 U256 ( .INP(input_factor_02[27]), .ZN(n585) );
  INVX0 U257 ( .INP(input_factor_01[24]), .ZN(n543) );
  NOR2X0 U258 ( .IN1(n543), .IN2(input_factor_02[24]), .QN(n39) );
  INVX0 U259 ( .INP(n39), .ZN(n25) );
  NAND4X0 U260 ( .IN1(n26), .IN2(n33), .IN3(n37), .IN4(n25), .QN(n27) );
  NOR4X0 U261 ( .IN1(n29), .IN2(n41), .IN3(n28), .IN4(n27), .QN(n31) );
  INVX0 U262 ( .INP(input_factor_01[30]), .ZN(n30) );
  INVX0 U263 ( .INP(n33), .ZN(n47) );
  INVX0 U264 ( .INP(n34), .ZN(n43) );
  INVX0 U265 ( .INP(n35), .ZN(n38) );
  OA221X1 U266 ( .IN1(n39), .IN2(n38), .IN3(n39), .IN4(n37), .IN5(n36), .Q(n40) );
  OA22X1 U267 ( .IN1(n41), .IN2(n40), .IN3(input_factor_01[26]), .IN4(n579), 
        .Q(n42) );
  OA22X1 U268 ( .IN1(n43), .IN2(n42), .IN3(input_factor_01[27]), .IN4(n585), 
        .Q(n46) );
  INVX0 U269 ( .INP(n44), .ZN(n45) );
  AO221X1 U270 ( .IN1(n48), .IN2(n47), .IN3(n48), .IN4(n46), .IN5(n45), .Q(n50) );
  AO221X1 U271 ( .IN1(n50), .IN2(n49), .IN3(n597), .IN4(input_factor_01[29]), 
        .IN5(input_factor_01[30]), .Q(n73) );
  INVX0 U272 ( .INP(n373), .ZN(n74) );
  INVX0 U273 ( .INP(input_factor_02[20]), .ZN(n695) );
  INVX0 U274 ( .INP(input_factor_02[16]), .ZN(n679) );
  INVX0 U275 ( .INP(input_factor_02[15]), .ZN(n673) );
  INVX0 U276 ( .INP(input_factor_02[11]), .ZN(n649) );
  INVX0 U277 ( .INP(input_factor_02[10]), .ZN(n643) );
  INVX0 U278 ( .INP(input_factor_02[9]), .ZN(n637) );
  INVX0 U279 ( .INP(input_factor_02[8]), .ZN(n633) );
  INVX0 U280 ( .INP(input_factor_02[7]), .ZN(n629) );
  INVX0 U281 ( .INP(input_factor_02[6]), .ZN(n625) );
  INVX0 U282 ( .INP(input_factor_02[5]), .ZN(n621) );
  INVX0 U283 ( .INP(input_factor_02[4]), .ZN(n617) );
  INVX0 U284 ( .INP(input_factor_02[3]), .ZN(n613) );
  INVX0 U285 ( .INP(input_factor_02[2]), .ZN(n609) );
  INVX0 U286 ( .INP(input_factor_01[0]), .ZN(n546) );
  NOR2X0 U287 ( .IN1(input_factor_02[0]), .IN2(n546), .QN(n51) );
  INVX0 U288 ( .INP(input_factor_02[1]), .ZN(n605) );
  AO222X1 U289 ( .IN1(input_factor_01[1]), .IN2(n51), .IN3(input_factor_01[1]), 
        .IN4(n605), .IN5(n51), .IN6(n605), .Q(n52) );
  AO222X1 U290 ( .IN1(input_factor_01[2]), .IN2(n609), .IN3(input_factor_01[2]), .IN4(n52), .IN5(n609), .IN6(n52), .Q(n53) );
  AO222X1 U291 ( .IN1(input_factor_01[3]), .IN2(n613), .IN3(input_factor_01[3]), .IN4(n53), .IN5(n613), .IN6(n53), .Q(n54) );
  AO222X1 U292 ( .IN1(input_factor_01[4]), .IN2(n617), .IN3(input_factor_01[4]), .IN4(n54), .IN5(n617), .IN6(n54), .Q(n55) );
  AO222X1 U293 ( .IN1(input_factor_01[5]), .IN2(n621), .IN3(input_factor_01[5]), .IN4(n55), .IN5(n621), .IN6(n55), .Q(n56) );
  AO222X1 U294 ( .IN1(input_factor_01[6]), .IN2(n625), .IN3(input_factor_01[6]), .IN4(n56), .IN5(n625), .IN6(n56), .Q(n57) );
  AO222X1 U295 ( .IN1(input_factor_01[7]), .IN2(n629), .IN3(input_factor_01[7]), .IN4(n57), .IN5(n629), .IN6(n57), .Q(n58) );
  AO222X1 U296 ( .IN1(input_factor_01[8]), .IN2(n633), .IN3(input_factor_01[8]), .IN4(n58), .IN5(n633), .IN6(n58), .Q(n59) );
  AO222X1 U297 ( .IN1(input_factor_01[9]), .IN2(n637), .IN3(input_factor_01[9]), .IN4(n59), .IN5(n637), .IN6(n59), .Q(n60) );
  AO222X1 U298 ( .IN1(input_factor_01[10]), .IN2(n643), .IN3(
        input_factor_01[10]), .IN4(n60), .IN5(n643), .IN6(n60), .Q(n61) );
  AO222X1 U299 ( .IN1(input_factor_01[11]), .IN2(n649), .IN3(
        input_factor_01[11]), .IN4(n61), .IN5(n649), .IN6(n61), .Q(n62) );
  AO222X1 U300 ( .IN1(input_factor_01[12]), .IN2(n655), .IN3(
        input_factor_01[12]), .IN4(n62), .IN5(n655), .IN6(n62), .Q(n63) );
  AO222X1 U301 ( .IN1(input_factor_01[13]), .IN2(n661), .IN3(
        input_factor_01[13]), .IN4(n63), .IN5(n661), .IN6(n63), .Q(n64) );
  AO222X1 U302 ( .IN1(input_factor_01[14]), .IN2(n667), .IN3(
        input_factor_01[14]), .IN4(n64), .IN5(n667), .IN6(n64), .Q(n65) );
  AO222X1 U303 ( .IN1(input_factor_01[15]), .IN2(n673), .IN3(
        input_factor_01[15]), .IN4(n65), .IN5(n673), .IN6(n65), .Q(n66) );
  AO222X1 U304 ( .IN1(input_factor_01[16]), .IN2(n679), .IN3(
        input_factor_01[16]), .IN4(n66), .IN5(n679), .IN6(n66), .Q(n68) );
  INVX0 U305 ( .INP(input_factor_01[17]), .ZN(n684) );
  INVX0 U306 ( .INP(input_factor_02[17]), .ZN(n685) );
  INVX0 U307 ( .INP(input_factor_01[18]), .ZN(n352) );
  INVX0 U308 ( .INP(input_factor_01[19]), .ZN(n356) );
  AO221X1 U309 ( .IN1(n68), .IN2(n67), .IN3(n685), .IN4(input_factor_01[17]), 
        .IN5(n545), .Q(n69) );
  AO222X1 U310 ( .IN1(input_factor_01[20]), .IN2(n695), .IN3(
        input_factor_01[20]), .IN4(n69), .IN5(n695), .IN6(n69), .Q(n71) );
  INVX0 U311 ( .INP(input_factor_01[21]), .ZN(n700) );
  INVX0 U312 ( .INP(input_factor_02[21]), .ZN(n703) );
  AO221X1 U313 ( .IN1(n71), .IN2(n70), .IN3(n703), .IN4(input_factor_01[21]), 
        .IN5(input_factor_01[22]), .Q(n123) );
  NOR2X0 U314 ( .IN1(n392), .IN2(n352), .QN(N194) );
  NOR2X0 U315 ( .IN1(n392), .IN2(n356), .QN(N195) );
  INVX0 U316 ( .INP(input_factor_01[22]), .ZN(n121) );
  NOR2X0 U317 ( .IN1(n392), .IN2(n121), .QN(N198) );
  AO22X1 U318 ( .IN1(input_factor_01[30]), .IN2(rst_n), .IN3(n848), .IN4(
        larger_exponent[7]), .Q(n826) );
  NOR4X0 U319 ( .IN1(exp_diff_value[4]), .IN2(exp_diff_value[5]), .IN3(
        exp_diff_value[6]), .IN4(exp_diff_value[7]), .QN(n370) );
  NOR2X0 U320 ( .IN1(exp_diff_value[3]), .IN2(n2), .QN(n371) );
  INVX0 U321 ( .INP(n371), .ZN(n213) );
  NOR2X0 U322 ( .IN1(n223), .IN2(n213), .QN(n280) );
  INVX0 U323 ( .INP(n280), .ZN(n357) );
  AO21X1 U324 ( .IN1(n121), .IN2(n1), .IN3(exp_diff_value[1]), .Q(n329) );
  INVX0 U325 ( .INP(n199), .ZN(n216) );
  OAI22X1 U326 ( .IN1(n326), .IN2(n357), .IN3(n329), .IN4(n364), .QN(N174) );
  INVX0 U328 ( .INP(input_factor_02[0]), .ZN(n124) );
  OA22X1 U329 ( .IN1(n605), .IN2(n326), .IN3(n124), .IN4(n207), .Q(n76) );
  OA22X1 U330 ( .IN1(n609), .IN2(n310), .IN3(n613), .IN4(n184), .Q(n75) );
  OA22X1 U331 ( .IN1(n633), .IN2(n207), .IN3(n637), .IN4(n326), .Q(n79) );
  OA22X1 U332 ( .IN1(n643), .IN2(n310), .IN3(n649), .IN4(n184), .Q(n77) );
  OA22X1 U333 ( .IN1(n655), .IN2(n207), .IN3(n661), .IN4(n326), .Q(n81) );
  OA22X1 U334 ( .IN1(n673), .IN2(n184), .IN3(n667), .IN4(n310), .Q(n80) );
  MUX21X1 U335 ( .IN1(n218), .IN2(n226), .S(n2), .Q(n285) );
  OA22X1 U336 ( .IN1(n617), .IN2(n207), .IN3(n621), .IN4(n326), .Q(n83) );
  OA22X1 U337 ( .IN1(n625), .IN2(n310), .IN3(n629), .IN4(n184), .Q(n82) );
  NOR2X0 U338 ( .IN1(exp_diff_value[3]), .IN2(n5), .QN(n188) );
  AOI222X1 U339 ( .IN1(n84), .IN2(n371), .IN3(n285), .IN4(exp_diff_value[3]), 
        .IN5(n219), .IN6(n188), .QN(n117) );
  AO22X1 U340 ( .IN1(input_factor_01[9]), .IN2(n202), .IN3(input_factor_01[8]), 
        .IN4(n372), .Q(n86) );
  AO22X1 U341 ( .IN1(input_factor_01[11]), .IN2(n204), .IN3(
        input_factor_01[10]), .IN4(n203), .Q(n85) );
  NOR2X0 U342 ( .IN1(n86), .IN2(n85), .QN(n217) );
  AO22X1 U343 ( .IN1(input_factor_01[13]), .IN2(n202), .IN3(
        input_factor_01[12]), .IN4(n372), .Q(n88) );
  AO22X1 U344 ( .IN1(input_factor_01[15]), .IN2(n204), .IN3(
        input_factor_01[14]), .IN4(n203), .Q(n87) );
  NOR2X0 U345 ( .IN1(n88), .IN2(n87), .QN(n215) );
  MUX21X1 U346 ( .IN1(n217), .IN2(n215), .S(n2), .Q(n287) );
  INVX0 U347 ( .INP(n188), .ZN(n198) );
  AO22X1 U348 ( .IN1(input_factor_01[5]), .IN2(n202), .IN3(input_factor_01[4]), 
        .IN4(n372), .Q(n90) );
  AO22X1 U349 ( .IN1(input_factor_01[7]), .IN2(n204), .IN3(input_factor_01[6]), 
        .IN4(n203), .Q(n89) );
  NOR2X0 U350 ( .IN1(n90), .IN2(n89), .QN(n221) );
  AO22X1 U351 ( .IN1(input_factor_01[0]), .IN2(n372), .IN3(input_factor_01[1]), 
        .IN4(n202), .Q(n92) );
  AO22X1 U352 ( .IN1(input_factor_01[3]), .IN2(n204), .IN3(input_factor_01[2]), 
        .IN4(n203), .Q(n91) );
  NOR2X0 U353 ( .IN1(n92), .IN2(n91), .QN(n93) );
  OA222X1 U354 ( .IN1(n4), .IN2(n287), .IN3(n198), .IN4(n221), .IN5(n213), 
        .IN6(n93), .Q(n116) );
  OA22X1 U355 ( .IN1(n117), .IN2(n223), .IN3(n116), .IN4(n199), .Q(n127) );
  AO221X1 U356 ( .IN1(exp_diff_value[0]), .IN2(n685), .IN3(n1), .IN4(n679), 
        .IN5(exp_diff_value[1]), .Q(n224) );
  OA22X1 U357 ( .IN1(input_factor_02[21]), .IN2(n326), .IN3(
        input_factor_02[20]), .IN4(exp_diff_value[0]), .Q(n311) );
  MUX21X1 U358 ( .IN1(n224), .IN2(n358), .S(n2), .Q(n343) );
  NOR3X0 U359 ( .IN1(exp_diff_value[5]), .IN2(exp_diff_value[6]), .IN3(
        exp_diff_value[7]), .QN(n118) );
  NOR2X0 U360 ( .IN1(exp_diff_value[3]), .IN2(n212), .QN(n122) );
  OA22X1 U361 ( .IN1(n352), .IN2(n310), .IN3(n684), .IN4(n326), .Q(n120) );
  INVX0 U362 ( .INP(input_factor_01[20]), .ZN(n694) );
  AO222X1 U363 ( .IN1(n203), .IN2(n121), .IN3(n202), .IN4(n700), .IN5(n372), 
        .IN6(n694), .Q(n359) );
  MUX21X1 U364 ( .IN1(n214), .IN2(n359), .S(n2), .Q(n342) );
  OA22X1 U365 ( .IN1(n343), .IN2(n235), .IN3(n342), .IN4(n208), .Q(n126) );
  OR2X1 U366 ( .IN1(n373), .IN2(n123), .Q(n366) );
  OA22X1 U367 ( .IN1(n124), .IN2(n367), .IN3(n546), .IN4(n366), .Q(n125) );
  NAND3X0 U368 ( .IN1(n127), .IN2(n126), .IN3(n125), .QN(N152) );
  OA22X1 U369 ( .IN1(n621), .IN2(n207), .IN3(n625), .IN4(n326), .Q(n129) );
  OA22X1 U370 ( .IN1(n633), .IN2(n184), .IN3(n629), .IN4(n310), .Q(n128) );
  OA22X1 U371 ( .IN1(n637), .IN2(n207), .IN3(n643), .IN4(n326), .Q(n131) );
  OA22X1 U372 ( .IN1(n655), .IN2(n184), .IN3(n649), .IN4(n310), .Q(n130) );
  OA22X1 U373 ( .IN1(n661), .IN2(n207), .IN3(n667), .IN4(n326), .Q(n133) );
  OA22X1 U374 ( .IN1(n673), .IN2(n310), .IN3(n679), .IN4(n184), .Q(n132) );
  MUX21X1 U375 ( .IN1(n244), .IN2(n236), .S(n2), .Q(n291) );
  OA22X1 U376 ( .IN1(n605), .IN2(n207), .IN3(n609), .IN4(n326), .Q(n135) );
  OA22X1 U377 ( .IN1(n613), .IN2(n310), .IN3(n617), .IN4(n184), .Q(n134) );
  AOI222X1 U378 ( .IN1(n240), .IN2(n188), .IN3(exp_diff_value[3]), .IN4(n291), 
        .IN5(n136), .IN6(n371), .QN(n148) );
  AO22X1 U379 ( .IN1(input_factor_01[10]), .IN2(n202), .IN3(input_factor_01[9]), .IN4(n372), .Q(n139) );
  AO22X1 U380 ( .IN1(input_factor_01[12]), .IN2(n204), .IN3(
        input_factor_01[11]), .IN4(n203), .Q(n137) );
  NOR2X0 U381 ( .IN1(n139), .IN2(n137), .QN(n239) );
  AO22X1 U382 ( .IN1(input_factor_01[14]), .IN2(n202), .IN3(
        input_factor_01[13]), .IN4(n372), .Q(n141) );
  AO22X1 U383 ( .IN1(input_factor_01[16]), .IN2(n204), .IN3(
        input_factor_01[15]), .IN4(n203), .Q(n140) );
  NOR2X0 U384 ( .IN1(n141), .IN2(n140), .QN(n232) );
  MUX21X1 U385 ( .IN1(n239), .IN2(n232), .S(n2), .Q(n293) );
  AO22X1 U386 ( .IN1(input_factor_01[6]), .IN2(n202), .IN3(input_factor_01[5]), 
        .IN4(n372), .Q(n143) );
  AO22X1 U387 ( .IN1(input_factor_01[8]), .IN2(n204), .IN3(input_factor_01[7]), 
        .IN4(n203), .Q(n142) );
  NOR2X0 U388 ( .IN1(n143), .IN2(n142), .QN(n233) );
  AO22X1 U389 ( .IN1(input_factor_01[2]), .IN2(n202), .IN3(input_factor_01[1]), 
        .IN4(n372), .Q(n145) );
  AO22X1 U390 ( .IN1(input_factor_01[4]), .IN2(n204), .IN3(input_factor_01[3]), 
        .IN4(n203), .Q(n144) );
  NOR2X0 U391 ( .IN1(n145), .IN2(n144), .QN(n146) );
  OA222X1 U392 ( .IN1(n4), .IN2(n293), .IN3(n198), .IN4(n233), .IN5(n213), 
        .IN6(n146), .Q(n147) );
  OA22X1 U393 ( .IN1(n148), .IN2(n223), .IN3(n147), .IN4(n199), .Q(n154) );
  AO22X1 U394 ( .IN1(input_factor_01[18]), .IN2(n202), .IN3(
        input_factor_01[17]), .IN4(n372), .Q(n150) );
  AO22X1 U395 ( .IN1(input_factor_01[20]), .IN2(n204), .IN3(
        input_factor_01[19]), .IN4(n203), .Q(n149) );
  NOR2X0 U396 ( .IN1(n150), .IN2(n149), .QN(n231) );
  AO22X1 U397 ( .IN1(input_factor_01[22]), .IN2(n202), .IN3(
        input_factor_01[21]), .IN4(n1), .Q(n151) );
  NOR2X0 U398 ( .IN1(n203), .IN2(n151), .QN(n365) );
  MUX21X1 U399 ( .IN1(n231), .IN2(n365), .S(n2), .Q(n347) );
  OA22X1 U400 ( .IN1(n685), .IN2(n207), .IN3(n695), .IN4(n184), .Q(n237) );
  AO21X1 U401 ( .IN1(n703), .IN2(n3), .IN3(exp_diff_value[0]), .Q(n234) );
  MUX21X1 U402 ( .IN1(n237), .IN2(n234), .S(n2), .Q(n346) );
  OA22X1 U403 ( .IN1(n208), .IN2(n347), .IN3(n235), .IN4(n346), .Q(n153) );
  INVX0 U404 ( .INP(input_factor_01[1]), .ZN(n604) );
  OA22X1 U405 ( .IN1(n605), .IN2(n367), .IN3(n604), .IN4(n366), .Q(n152) );
  NAND3X0 U406 ( .IN1(n154), .IN2(n153), .IN3(n152), .QN(N153) );
  OA22X1 U407 ( .IN1(n625), .IN2(n207), .IN3(n629), .IN4(n326), .Q(n156) );
  OA22X1 U408 ( .IN1(n633), .IN2(n310), .IN3(n637), .IN4(n184), .Q(n155) );
  OA22X1 U409 ( .IN1(n643), .IN2(n207), .IN3(n649), .IN4(n326), .Q(n158) );
  OA22X1 U410 ( .IN1(n655), .IN2(n310), .IN3(n661), .IN4(n184), .Q(n157) );
  OA22X1 U411 ( .IN1(n673), .IN2(n326), .IN3(n667), .IN4(n207), .Q(n160) );
  OA22X1 U412 ( .IN1(n679), .IN2(n310), .IN3(n685), .IN4(n184), .Q(n159) );
  MUX21X1 U413 ( .IN1(n249), .IN2(n257), .S(n2), .Q(n297) );
  OA22X1 U414 ( .IN1(n609), .IN2(n207), .IN3(n613), .IN4(n326), .Q(n162) );
  OA22X1 U415 ( .IN1(n617), .IN2(n310), .IN3(n621), .IN4(n184), .Q(n161) );
  AOI222X1 U416 ( .IN1(n250), .IN2(n188), .IN3(exp_diff_value[3]), .IN4(n297), 
        .IN5(n163), .IN6(n371), .QN(n174) );
  AO22X1 U417 ( .IN1(input_factor_01[11]), .IN2(n202), .IN3(
        input_factor_01[10]), .IN4(n372), .Q(n165) );
  AO22X1 U418 ( .IN1(input_factor_01[13]), .IN2(n204), .IN3(
        input_factor_01[12]), .IN4(n203), .Q(n164) );
  NOR2X0 U419 ( .IN1(n165), .IN2(n164), .QN(n261) );
  AO22X1 U420 ( .IN1(input_factor_01[15]), .IN2(n202), .IN3(
        input_factor_01[14]), .IN4(n372), .Q(n167) );
  AO22X1 U421 ( .IN1(input_factor_01[17]), .IN2(n204), .IN3(
        input_factor_01[16]), .IN4(n203), .Q(n166) );
  NOR2X0 U422 ( .IN1(n167), .IN2(n166), .QN(n256) );
  MUX21X1 U423 ( .IN1(n261), .IN2(n256), .S(n2), .Q(n299) );
  AO22X1 U424 ( .IN1(input_factor_01[7]), .IN2(n202), .IN3(input_factor_01[6]), 
        .IN4(n372), .Q(n169) );
  AO22X1 U425 ( .IN1(input_factor_01[9]), .IN2(n204), .IN3(input_factor_01[8]), 
        .IN4(n203), .Q(n168) );
  NOR2X0 U426 ( .IN1(n169), .IN2(n168), .QN(n252) );
  AO22X1 U427 ( .IN1(input_factor_01[3]), .IN2(n202), .IN3(input_factor_01[2]), 
        .IN4(n372), .Q(n171) );
  AO22X1 U428 ( .IN1(input_factor_01[5]), .IN2(n204), .IN3(input_factor_01[4]), 
        .IN4(n203), .Q(n170) );
  NOR2X0 U429 ( .IN1(n171), .IN2(n170), .QN(n172) );
  OA222X1 U430 ( .IN1(n4), .IN2(n299), .IN3(n198), .IN4(n252), .IN5(n213), 
        .IN6(n172), .Q(n173) );
  OA22X1 U431 ( .IN1(n174), .IN2(n223), .IN3(n173), .IN4(n199), .Q(n179) );
  AO22X1 U432 ( .IN1(input_factor_01[18]), .IN2(n372), .IN3(
        input_factor_01[19]), .IN4(n202), .Q(n176) );
  AO22X1 U433 ( .IN1(input_factor_01[21]), .IN2(n204), .IN3(
        input_factor_01[20]), .IN4(n203), .Q(n175) );
  NOR2X0 U434 ( .IN1(n176), .IN2(n175), .QN(n255) );
  MUX21X1 U435 ( .IN1(n255), .IN2(n329), .S(n2), .Q(n350) );
  OA22X1 U436 ( .IN1(n695), .IN2(n310), .IN3(n703), .IN4(n184), .Q(n258) );
  MUX21X1 U437 ( .IN1(n258), .IN2(n326), .S(n2), .Q(n351) );
  OA22X1 U438 ( .IN1(n350), .IN2(n208), .IN3(n351), .IN4(n235), .Q(n178) );
  INVX0 U439 ( .INP(input_factor_01[2]), .ZN(n608) );
  OA22X1 U440 ( .IN1(n609), .IN2(n367), .IN3(n608), .IN4(n366), .Q(n177) );
  NAND3X0 U441 ( .IN1(n179), .IN2(n178), .IN3(n177), .QN(N154) );
  OA22X1 U442 ( .IN1(n633), .IN2(n326), .IN3(n629), .IN4(n207), .Q(n181) );
  OA22X1 U443 ( .IN1(n637), .IN2(n310), .IN3(n643), .IN4(n184), .Q(n180) );
  OA22X1 U444 ( .IN1(n655), .IN2(n326), .IN3(n649), .IN4(n207), .Q(n183) );
  OA22X1 U445 ( .IN1(n661), .IN2(n310), .IN3(n667), .IN4(n184), .Q(n182) );
  AO222X1 U446 ( .IN1(input_factor_02[15]), .IN2(n372), .IN3(
        input_factor_02[17]), .IN4(n203), .IN5(input_factor_02[16]), .IN6(n202), .Q(n278) );
  MUX21X1 U447 ( .IN1(n269), .IN2(n278), .S(n2), .Q(n303) );
  OA22X1 U448 ( .IN1(n613), .IN2(n207), .IN3(n617), .IN4(n326), .Q(n186) );
  OA22X1 U449 ( .IN1(n621), .IN2(n310), .IN3(n625), .IN4(n184), .Q(n185) );
  AOI222X1 U450 ( .IN1(n279), .IN2(n188), .IN3(exp_diff_value[3]), .IN4(n303), 
        .IN5(n187), .IN6(n371), .QN(n201) );
  AO22X1 U451 ( .IN1(input_factor_01[12]), .IN2(n202), .IN3(
        input_factor_01[11]), .IN4(n372), .Q(n190) );
  AO22X1 U452 ( .IN1(input_factor_01[14]), .IN2(n204), .IN3(
        input_factor_01[13]), .IN4(n203), .Q(n189) );
  NOR2X0 U453 ( .IN1(n190), .IN2(n189), .QN(n274) );
  AO22X1 U454 ( .IN1(input_factor_01[16]), .IN2(n202), .IN3(
        input_factor_01[15]), .IN4(n372), .Q(n192) );
  AO22X1 U455 ( .IN1(input_factor_01[18]), .IN2(n204), .IN3(
        input_factor_01[17]), .IN4(n203), .Q(n191) );
  NOR2X0 U456 ( .IN1(n192), .IN2(n191), .QN(n268) );
  MUX21X1 U457 ( .IN1(n274), .IN2(n268), .S(n2), .Q(n305) );
  AO22X1 U458 ( .IN1(input_factor_01[8]), .IN2(n202), .IN3(input_factor_01[7]), 
        .IN4(n372), .Q(n194) );
  AO22X1 U459 ( .IN1(input_factor_01[10]), .IN2(n204), .IN3(input_factor_01[9]), .IN4(n203), .Q(n193) );
  NOR2X0 U460 ( .IN1(n194), .IN2(n193), .QN(n275) );
  AO22X1 U461 ( .IN1(input_factor_01[4]), .IN2(n202), .IN3(input_factor_01[3]), 
        .IN4(n372), .Q(n196) );
  AO22X1 U462 ( .IN1(input_factor_01[6]), .IN2(n204), .IN3(input_factor_01[5]), 
        .IN4(n203), .Q(n195) );
  NOR2X0 U463 ( .IN1(n196), .IN2(n195), .QN(n197) );
  OA222X1 U464 ( .IN1(n4), .IN2(n305), .IN3(n198), .IN4(n275), .IN5(n213), 
        .IN6(n197), .Q(n200) );
  OA22X1 U465 ( .IN1(n201), .IN2(n223), .IN3(n200), .IN4(n199), .Q(n211) );
  AO22X1 U466 ( .IN1(input_factor_01[20]), .IN2(n202), .IN3(
        input_factor_01[19]), .IN4(n372), .Q(n206) );
  AO22X1 U467 ( .IN1(input_factor_01[22]), .IN2(n204), .IN3(
        input_factor_01[21]), .IN4(n203), .Q(n205) );
  NOR2X0 U468 ( .IN1(n206), .IN2(n205), .QN(n267) );
  MUX21X1 U469 ( .IN1(n267), .IN2(n207), .S(n2), .Q(n353) );
  OA22X1 U470 ( .IN1(n695), .IN2(n326), .IN3(n703), .IN4(n310), .Q(n276) );
  MUX21X1 U471 ( .IN1(n276), .IN2(n207), .S(n2), .Q(n355) );
  OA22X1 U472 ( .IN1(n353), .IN2(n208), .IN3(n355), .IN4(n235), .Q(n210) );
  INVX0 U473 ( .INP(input_factor_01[3]), .ZN(n612) );
  OA22X1 U474 ( .IN1(n613), .IN2(n367), .IN3(n612), .IN4(n366), .Q(n209) );
  NAND3X0 U475 ( .IN1(n211), .IN2(n210), .IN3(n209), .QN(N155) );
  NOR2X0 U476 ( .IN1(n213), .IN2(n212), .QN(n266) );
  OA22X1 U477 ( .IN1(n359), .IN2(n253), .IN3(n358), .IN4(n254), .Q(n230) );
  OR2X1 U478 ( .IN1(n5), .IN2(n354), .Q(n273) );
  MUX21X1 U479 ( .IN1(n215), .IN2(n214), .S(n2), .Q(n309) );
  OA22X1 U480 ( .IN1(n217), .IN2(n273), .IN3(n309), .IN4(n336), .Q(n229) );
  NOR2X0 U481 ( .IN1(n223), .IN2(exp_diff_value[3]), .QN(n313) );
  NOR2X0 U482 ( .IN1(n5), .IN2(n362), .QN(n270) );
  AOI22X1 U483 ( .IN1(n280), .IN2(n219), .IN3(n270), .IN4(n218), .QN(n222) );
  INVX0 U484 ( .INP(input_factor_01[4]), .ZN(n616) );
  OA22X1 U485 ( .IN1(n617), .IN2(n367), .IN3(n616), .IN4(n366), .Q(n220) );
  NOR2X0 U486 ( .IN1(n223), .IN2(n4), .QN(n323) );
  INVX0 U487 ( .INP(n224), .ZN(n225) );
  MUX21X1 U488 ( .IN1(n226), .IN2(n225), .S(n2), .Q(n312) );
  NAND4X0 U489 ( .IN1(n230), .IN2(n229), .IN3(n228), .IN4(n227), .QN(N156) );
  MUX21X1 U490 ( .IN1(n232), .IN2(n231), .S(n2), .Q(n318) );
  OA22X1 U491 ( .IN1(n233), .IN2(n364), .IN3(n318), .IN4(n336), .Q(n248) );
  OR2X1 U492 ( .IN1(n2), .IN2(n234), .Q(n363) );
  OA22X1 U493 ( .IN1(n365), .IN2(n253), .IN3(n235), .IN4(n363), .Q(n243) );
  INVX0 U494 ( .INP(n236), .ZN(n238) );
  MUX21X1 U495 ( .IN1(n238), .IN2(n237), .S(n2), .Q(n319) );
  INVX0 U496 ( .INP(n323), .ZN(n337) );
  OA22X1 U497 ( .IN1(n239), .IN2(n273), .IN3(n319), .IN4(n337), .Q(n242) );
  AND3X1 U498 ( .IN1(n243), .IN2(n242), .IN3(n241), .Q(n247) );
  INVX0 U499 ( .INP(input_factor_01[5]), .ZN(n620) );
  OA22X1 U500 ( .IN1(n621), .IN2(n367), .IN3(n620), .IN4(n366), .Q(n246) );
  NAND4X0 U501 ( .IN1(n248), .IN2(n247), .IN3(n246), .IN4(n245), .QN(N157) );
  AOI22X1 U502 ( .IN1(n280), .IN2(n250), .IN3(n270), .IN4(n249), .QN(n251) );
  OA21X1 U503 ( .IN1(n252), .IN2(n364), .IN3(n251), .Q(n265) );
  OA22X1 U504 ( .IN1(n326), .IN2(n254), .IN3(n329), .IN4(n253), .Q(n264) );
  MUX21X1 U505 ( .IN1(n256), .IN2(n255), .S(n2), .Q(n327) );
  INVX0 U506 ( .INP(n257), .ZN(n259) );
  MUX21X1 U507 ( .IN1(n259), .IN2(n258), .S(n2), .Q(n324) );
  OA22X1 U508 ( .IN1(n336), .IN2(n327), .IN3(n337), .IN4(n324), .Q(n260) );
  OA21X1 U509 ( .IN1(n261), .IN2(n273), .IN3(n260), .Q(n263) );
  INVX0 U510 ( .INP(input_factor_01[6]), .ZN(n624) );
  OA22X1 U511 ( .IN1(n625), .IN2(n367), .IN3(n624), .IN4(n366), .Q(n262) );
  NAND4X0 U512 ( .IN1(n265), .IN2(n264), .IN3(n263), .IN4(n262), .QN(N158) );
  NAND3X0 U513 ( .IN1(n372), .IN2(n266), .IN3(n373), .QN(n272) );
  MUX21X1 U514 ( .IN1(n268), .IN2(n267), .S(n2), .Q(n334) );
  OA22X1 U515 ( .IN1(n275), .IN2(n364), .IN3(n274), .IN4(n273), .Q(n283) );
  INVX0 U516 ( .INP(n276), .ZN(n277) );
  MUX21X1 U517 ( .IN1(n278), .IN2(n277), .S(n2), .Q(n333) );
  AOI22X1 U518 ( .IN1(n333), .IN2(n323), .IN3(n280), .IN4(n279), .QN(n282) );
  INVX0 U519 ( .INP(input_factor_01[7]), .ZN(n628) );
  OA22X1 U520 ( .IN1(n629), .IN2(n367), .IN3(n628), .IN4(n366), .Q(n281) );
  NAND4X0 U521 ( .IN1(n284), .IN2(n283), .IN3(n282), .IN4(n281), .QN(N159) );
  INVX0 U522 ( .INP(n285), .ZN(n286) );
  OA22X1 U523 ( .IN1(n342), .IN2(n336), .IN3(n286), .IN4(n362), .Q(n290) );
  OA22X1 U524 ( .IN1(n343), .IN2(n337), .IN3(n287), .IN4(n354), .Q(n289) );
  INVX0 U525 ( .INP(input_factor_01[8]), .ZN(n632) );
  OA22X1 U526 ( .IN1(n633), .IN2(n367), .IN3(n632), .IN4(n366), .Q(n288) );
  NAND3X0 U527 ( .IN1(n290), .IN2(n289), .IN3(n288), .QN(N160) );
  INVX0 U528 ( .INP(n291), .ZN(n292) );
  OA22X1 U529 ( .IN1(n292), .IN2(n362), .IN3(n347), .IN4(n336), .Q(n296) );
  OA22X1 U530 ( .IN1(n293), .IN2(n354), .IN3(n346), .IN4(n337), .Q(n295) );
  INVX0 U531 ( .INP(input_factor_01[9]), .ZN(n636) );
  OA22X1 U532 ( .IN1(n637), .IN2(n367), .IN3(n636), .IN4(n366), .Q(n294) );
  NAND3X0 U533 ( .IN1(n296), .IN2(n295), .IN3(n294), .QN(N161) );
  INVX0 U534 ( .INP(n297), .ZN(n298) );
  OA22X1 U535 ( .IN1(n350), .IN2(n336), .IN3(n298), .IN4(n362), .Q(n302) );
  OA22X1 U536 ( .IN1(n351), .IN2(n337), .IN3(n299), .IN4(n354), .Q(n301) );
  INVX0 U537 ( .INP(input_factor_01[10]), .ZN(n642) );
  OA22X1 U538 ( .IN1(n643), .IN2(n367), .IN3(n642), .IN4(n366), .Q(n300) );
  NAND3X0 U539 ( .IN1(n302), .IN2(n301), .IN3(n300), .QN(N162) );
  INVX0 U540 ( .INP(n303), .ZN(n304) );
  OA22X1 U541 ( .IN1(n353), .IN2(n336), .IN3(n304), .IN4(n362), .Q(n308) );
  OA22X1 U542 ( .IN1(n355), .IN2(n337), .IN3(n305), .IN4(n354), .Q(n307) );
  INVX0 U543 ( .INP(input_factor_01[11]), .ZN(n648) );
  OA22X1 U544 ( .IN1(n649), .IN2(n367), .IN3(n648), .IN4(n366), .Q(n306) );
  NAND3X0 U545 ( .IN1(n308), .IN2(n307), .IN3(n306), .QN(N163) );
  OR2X1 U546 ( .IN1(n336), .IN2(n2), .Q(n328) );
  OA22X1 U547 ( .IN1(n359), .IN2(n328), .IN3(n354), .IN4(n309), .Q(n317) );
  INVX0 U548 ( .INP(input_factor_01[12]), .ZN(n654) );
  OA22X1 U549 ( .IN1(n655), .IN2(n367), .IN3(n654), .IN4(n366), .Q(n316) );
  NAND4X0 U550 ( .IN1(n311), .IN2(n323), .IN3(n5), .IN4(n310), .QN(n315) );
  NAND4X0 U551 ( .IN1(n317), .IN2(n316), .IN3(n315), .IN4(n314), .QN(N164) );
  OA22X1 U552 ( .IN1(n362), .IN2(n319), .IN3(n354), .IN4(n318), .Q(n322) );
  OA22X1 U553 ( .IN1(n365), .IN2(n328), .IN3(n363), .IN4(n337), .Q(n321) );
  INVX0 U554 ( .INP(input_factor_01[13]), .ZN(n660) );
  OA22X1 U555 ( .IN1(n661), .IN2(n367), .IN3(n660), .IN4(n366), .Q(n320) );
  NAND3X0 U556 ( .IN1(n322), .IN2(n321), .IN3(n320), .QN(N165) );
  OA22X1 U557 ( .IN1(n326), .IN2(n325), .IN3(n362), .IN4(n324), .Q(n332) );
  OA22X1 U558 ( .IN1(n329), .IN2(n328), .IN3(n354), .IN4(n327), .Q(n331) );
  INVX0 U559 ( .INP(input_factor_01[14]), .ZN(n666) );
  OA22X1 U560 ( .IN1(n667), .IN2(n367), .IN3(n666), .IN4(n366), .Q(n330) );
  NAND3X0 U561 ( .IN1(n332), .IN2(n331), .IN3(n330), .QN(N166) );
  INVX0 U562 ( .INP(n333), .ZN(n335) );
  OA22X1 U563 ( .IN1(n362), .IN2(n335), .IN3(n354), .IN4(n334), .Q(n341) );
  INVX0 U564 ( .INP(input_factor_01[15]), .ZN(n672) );
  OA22X1 U565 ( .IN1(n673), .IN2(n367), .IN3(n672), .IN4(n366), .Q(n340) );
  NAND3X0 U566 ( .IN1(n338), .IN2(n5), .IN3(n372), .QN(n339) );
  NAND3X0 U567 ( .IN1(n341), .IN2(n340), .IN3(n339), .QN(N167) );
  OA22X1 U568 ( .IN1(n343), .IN2(n362), .IN3(n342), .IN4(n354), .Q(n345) );
  INVX0 U569 ( .INP(input_factor_01[16]), .ZN(n678) );
  OA22X1 U570 ( .IN1(n679), .IN2(n367), .IN3(n678), .IN4(n366), .Q(n344) );
  OA22X1 U571 ( .IN1(n347), .IN2(n354), .IN3(n346), .IN4(n362), .Q(n349) );
  OA22X1 U572 ( .IN1(n685), .IN2(n367), .IN3(n684), .IN4(n366), .Q(n348) );
  OAI222X1 U573 ( .IN1(n366), .IN2(n352), .IN3(n362), .IN4(n351), .IN5(n354), 
        .IN6(n350), .QN(N170) );
  OAI222X1 U574 ( .IN1(n366), .IN2(n356), .IN3(n362), .IN4(n355), .IN5(n354), 
        .IN6(n353), .QN(N171) );
  OA22X1 U575 ( .IN1(n359), .IN2(n364), .IN3(n358), .IN4(n357), .Q(n361) );
  OA22X1 U576 ( .IN1(n695), .IN2(n367), .IN3(n694), .IN4(n366), .Q(n360) );
  OA22X1 U577 ( .IN1(n365), .IN2(n364), .IN3(n363), .IN4(n362), .Q(n369) );
  OA22X1 U578 ( .IN1(n703), .IN2(n367), .IN3(n700), .IN4(n366), .Q(n368) );
  NAND3X0 U579 ( .IN1(n372), .IN2(n371), .IN3(n370), .QN(n374) );
  MUX21X1 U580 ( .IN1(input_factor_01[0]), .IN2(input_factor_02[0]), .S(n392), 
        .Q(N176) );
  MUX21X1 U581 ( .IN1(input_factor_01[1]), .IN2(input_factor_02[1]), .S(n392), 
        .Q(N177) );
  MUX21X1 U582 ( .IN1(input_factor_01[2]), .IN2(input_factor_02[2]), .S(n392), 
        .Q(N178) );
  MUX21X1 U583 ( .IN1(input_factor_01[3]), .IN2(input_factor_02[3]), .S(n392), 
        .Q(N179) );
  MUX21X1 U584 ( .IN1(input_factor_01[4]), .IN2(input_factor_02[4]), .S(n392), 
        .Q(N180) );
  MUX21X1 U585 ( .IN1(input_factor_01[5]), .IN2(input_factor_02[5]), .S(n392), 
        .Q(N181) );
  MUX21X1 U586 ( .IN1(input_factor_01[6]), .IN2(input_factor_02[6]), .S(n392), 
        .Q(N182) );
  MUX21X1 U587 ( .IN1(input_factor_01[7]), .IN2(input_factor_02[7]), .S(n392), 
        .Q(N183) );
  MUX21X1 U588 ( .IN1(input_factor_01[8]), .IN2(input_factor_02[8]), .S(n392), 
        .Q(N184) );
  MUX21X1 U589 ( .IN1(input_factor_01[9]), .IN2(input_factor_02[9]), .S(n392), 
        .Q(N185) );
  MUX21X1 U590 ( .IN1(input_factor_01[10]), .IN2(input_factor_02[10]), .S(n392), .Q(N186) );
  MUX21X1 U591 ( .IN1(input_factor_01[11]), .IN2(input_factor_02[11]), .S(n392), .Q(N187) );
  MUX21X1 U592 ( .IN1(input_factor_01[12]), .IN2(input_factor_02[12]), .S(n392), .Q(N188) );
  MUX21X1 U593 ( .IN1(input_factor_01[13]), .IN2(input_factor_02[13]), .S(n392), .Q(N189) );
  MUX21X1 U594 ( .IN1(input_factor_01[14]), .IN2(input_factor_02[14]), .S(n392), .Q(N190) );
  MUX21X1 U595 ( .IN1(input_factor_01[15]), .IN2(input_factor_02[15]), .S(n392), .Q(N191) );
  MUX21X1 U596 ( .IN1(input_factor_01[16]), .IN2(input_factor_02[16]), .S(n392), .Q(N192) );
  MUX21X1 U597 ( .IN1(input_factor_01[17]), .IN2(input_factor_02[17]), .S(n392), .Q(N193) );
  MUX21X1 U598 ( .IN1(input_factor_01[20]), .IN2(input_factor_02[20]), .S(n392), .Q(N196) );
  MUX21X1 U599 ( .IN1(input_factor_01[21]), .IN2(input_factor_02[21]), .S(n392), .Q(N197) );
  MUX21X1 U600 ( .IN1(add_result[0]), .IN2(sub_result[0]), .S(n503), .Q(n818)
         );
  MUX21X1 U601 ( .IN1(add_result[2]), .IN2(sub_result[2]), .S(n503), .Q(n796)
         );
  MUX21X1 U602 ( .IN1(add_result[3]), .IN2(sub_result[3]), .S(n503), .Q(n788)
         );
  MUX21X1 U603 ( .IN1(add_result[4]), .IN2(sub_result[4]), .S(n503), .Q(n797)
         );
  MUX21X1 U604 ( .IN1(add_result[5]), .IN2(sub_result[5]), .S(n503), .Q(n789)
         );
  MUX21X1 U605 ( .IN1(add_result[6]), .IN2(sub_result[6]), .S(n503), .Q(n764)
         );
  MUX21X1 U606 ( .IN1(add_result[7]), .IN2(sub_result[7]), .S(n503), .Q(n756)
         );
  MUX21X1 U607 ( .IN1(add_result[9]), .IN2(sub_result[9]), .S(n503), .Q(n740)
         );
  MUX21X1 U608 ( .IN1(add_result[10]), .IN2(sub_result[10]), .S(n503), .Q(n732) );
  NOR4X0 U609 ( .IN1(n503), .IN2(add_result[14]), .IN3(add_result[15]), .IN4(
        add_result[13]), .QN(n512) );
  NOR4X0 U610 ( .IN1(sub_result[15]), .IN2(sub_result[14]), .IN3(
        sub_result[13]), .IN4(n21), .QN(n510) );
  NOR2X0 U611 ( .IN1(n512), .IN2(n510), .QN(n379) );
  MUX21X1 U612 ( .IN1(add_result[11]), .IN2(sub_result[11]), .S(n503), .Q(n724) );
  MUX21X1 U613 ( .IN1(add_result[16]), .IN2(sub_result[16]), .S(n20), .Q(n396)
         );
  MUX21X1 U614 ( .IN1(add_result[17]), .IN2(sub_result[17]), .S(n20), .Q(n465)
         );
  MUX21X1 U615 ( .IN1(add_result[20]), .IN2(sub_result[20]), .S(n20), .Q(n399)
         );
  INVX0 U616 ( .INP(n399), .ZN(n492) );
  MUX21X1 U617 ( .IN1(add_result[22]), .IN2(sub_result[22]), .S(n20), .Q(n400)
         );
  INVX0 U618 ( .INP(n400), .ZN(n376) );
  MUX21X1 U619 ( .IN1(add_result[23]), .IN2(sub_result[23]), .S(n20), .Q(n395)
         );
  MUX21X1 U620 ( .IN1(add_result[21]), .IN2(sub_result[21]), .S(n20), .Q(n402)
         );
  NOR2X0 U621 ( .IN1(n403), .IN2(n402), .QN(n404) );
  MUX21X1 U622 ( .IN1(add_result[19]), .IN2(sub_result[19]), .S(n20), .Q(n474)
         );
  NOR2X0 U623 ( .IN1(n377), .IN2(n474), .QN(n401) );
  MUX21X1 U624 ( .IN1(add_result[18]), .IN2(sub_result[18]), .S(n20), .Q(n398)
         );
  NOR2X0 U625 ( .IN1(n465), .IN2(n378), .QN(n397) );
  MUX21X1 U626 ( .IN1(add_result[12]), .IN2(sub_result[12]), .S(n20), .Q(n442)
         );
  NOR4X0 U627 ( .IN1(n379), .IN2(n724), .IN3(n559), .IN4(n442), .QN(n719) );
  MUX21X1 U628 ( .IN1(add_result[8]), .IN2(sub_result[8]), .S(n20), .Q(n748)
         );
  NOR3X0 U629 ( .IN1(n740), .IN2(n556), .IN3(n748), .QN(n517) );
  NOR2X0 U630 ( .IN1(n764), .IN2(n380), .QN(n516) );
  NOR2X0 U631 ( .IN1(n797), .IN2(n381), .QN(n524) );
  NOR2X0 U632 ( .IN1(n796), .IN2(n382), .QN(n518) );
  NAND3X0 U633 ( .IN1(n810), .IN2(n802), .IN3(n518), .QN(n557) );
  NAND4X0 U634 ( .IN1(n655), .IN2(n673), .IN3(n661), .IN4(n667), .QN(n391) );
  OR4X1 U635 ( .IN1(input_factor_02[31]), .IN2(input_factor_02[27]), .IN3(
        input_factor_02[24]), .IN4(input_factor_02[25]), .Q(n390) );
  NAND4X0 U636 ( .IN1(n597), .IN2(n383), .IN3(n591), .IN4(n579), .QN(n389) );
  NOR4X0 U637 ( .IN1(input_factor_02[1]), .IN2(input_factor_02[0]), .IN3(
        input_factor_02[2]), .IN4(input_factor_02[3]), .QN(n387) );
  NOR4X0 U638 ( .IN1(input_factor_02[16]), .IN2(input_factor_02[17]), .IN3(
        input_factor_02[20]), .IN4(input_factor_02[21]), .QN(n386) );
  NOR4X0 U639 ( .IN1(input_factor_02[7]), .IN2(input_factor_02[9]), .IN3(
        input_factor_02[10]), .IN4(input_factor_02[11]), .QN(n385) );
  NOR4X0 U640 ( .IN1(input_factor_02[4]), .IN2(input_factor_02[5]), .IN3(
        input_factor_02[8]), .IN4(input_factor_02[6]), .QN(n384) );
  NAND4X0 U641 ( .IN1(n387), .IN2(n386), .IN3(n385), .IN4(n384), .QN(n388) );
  AO222X1 U642 ( .IN1(input_factor_01[31]), .IN2(n710), .IN3(
        input_factor_01[31]), .IN4(n393), .IN5(n392), .IN6(input_factor_02[31]), .Q(n394) );
  AND2X1 U643 ( .IN1(n557), .IN2(n394), .Q(N211) );
  MUX21X1 U644 ( .IN1(n818), .IN2(n816), .S(add_sub_result_24_), .Q(N226) );
  MUX21X1 U645 ( .IN1(n816), .IN2(n796), .S(add_sub_result_24_), .Q(N227) );
  MUX21X1 U646 ( .IN1(n796), .IN2(n788), .S(add_sub_result_24_), .Q(N228) );
  MUX21X1 U647 ( .IN1(n788), .IN2(n797), .S(add_sub_result_24_), .Q(N229) );
  MUX21X1 U648 ( .IN1(n797), .IN2(n789), .S(add_sub_result_24_), .Q(N230) );
  MUX21X1 U649 ( .IN1(n789), .IN2(n764), .S(add_sub_result_24_), .Q(N231) );
  MUX21X1 U650 ( .IN1(n764), .IN2(n756), .S(add_sub_result_24_), .Q(N232) );
  MUX21X1 U651 ( .IN1(n756), .IN2(n748), .S(add_sub_result_24_), .Q(N233) );
  MUX21X1 U652 ( .IN1(n748), .IN2(n740), .S(add_sub_result_24_), .Q(N234) );
  MUX21X1 U653 ( .IN1(n740), .IN2(n732), .S(add_sub_result_24_), .Q(N235) );
  MUX21X1 U654 ( .IN1(n732), .IN2(n724), .S(add_sub_result_24_), .Q(N236) );
  MUX21X1 U655 ( .IN1(n724), .IN2(n442), .S(add_sub_result_24_), .Q(N237) );
  MUX21X1 U656 ( .IN1(add_result[13]), .IN2(sub_result[13]), .S(n20), .Q(n447)
         );
  MUX21X1 U657 ( .IN1(n442), .IN2(n447), .S(add_sub_result_24_), .Q(N238) );
  MUX21X1 U658 ( .IN1(add_result[14]), .IN2(sub_result[14]), .S(n20), .Q(n501)
         );
  MUX21X1 U659 ( .IN1(n447), .IN2(n501), .S(add_sub_result_24_), .Q(N239) );
  MUX21X1 U660 ( .IN1(add_result[15]), .IN2(sub_result[15]), .S(n20), .Q(n456)
         );
  MUX21X1 U661 ( .IN1(n501), .IN2(n456), .S(add_sub_result_24_), .Q(N240) );
  MUX21X1 U662 ( .IN1(n456), .IN2(n396), .S(add_sub_result_24_), .Q(N241) );
  MUX21X1 U663 ( .IN1(n396), .IN2(n465), .S(add_sub_result_24_), .Q(N242) );
  MUX21X1 U664 ( .IN1(n465), .IN2(n398), .S(add_sub_result_24_), .Q(N243) );
  MUX21X1 U665 ( .IN1(n398), .IN2(n474), .S(add_sub_result_24_), .Q(N244) );
  MUX21X1 U666 ( .IN1(n474), .IN2(n399), .S(add_sub_result_24_), .Q(N245) );
  MUX21X1 U667 ( .IN1(n399), .IN2(n402), .S(add_sub_result_24_), .Q(N246) );
  MUX21X1 U668 ( .IN1(n402), .IN2(n400), .S(add_sub_result_24_), .Q(N247) );
  MUX21X1 U669 ( .IN1(n400), .IN2(n395), .S(add_sub_result_24_), .Q(N248) );
  NAND4X0 U670 ( .IN1(n496), .IN2(n485), .IN3(n489), .IN4(n487), .QN(N256) );
  INVX0 U671 ( .INP(n402), .ZN(n488) );
  NOR2X0 U672 ( .IN1(n488), .IN2(n403), .QN(n419) );
  NAND4X0 U673 ( .IN1(n496), .IN2(n483), .IN3(n489), .IN4(n491), .QN(N257) );
  NAND3X0 U674 ( .IN1(n404), .IN2(n492), .IN3(n474), .QN(n493) );
  NAND4X0 U675 ( .IN1(n496), .IN2(n485), .IN3(n493), .IN4(n483), .QN(N258) );
  NOR2X0 U676 ( .IN1(n810), .IN2(n487), .QN(N260) );
  INVX0 U677 ( .INP(n487), .ZN(n421) );
  AO22X1 U678 ( .IN1(n421), .IN2(n816), .IN3(n419), .IN4(n818), .Q(N261) );
  INVX0 U679 ( .INP(n489), .ZN(n420) );
  AO222X1 U680 ( .IN1(n818), .IN2(n420), .IN3(n816), .IN4(n419), .IN5(n796), 
        .IN6(n421), .Q(N262) );
  OA22X1 U681 ( .IN1(n802), .IN2(n489), .IN3(n810), .IN4(n493), .Q(n406) );
  OA22X1 U682 ( .IN1(n808), .IN2(n491), .IN3(n806), .IN4(n487), .Q(n405) );
  OA22X1 U683 ( .IN1(n786), .IN2(n487), .IN3(n806), .IN4(n491), .Q(n409) );
  OA22X1 U684 ( .IN1(n802), .IN2(n493), .IN3(n810), .IN4(n485), .Q(n408) );
  NAND3X0 U685 ( .IN1(n409), .IN2(n408), .IN3(n407), .QN(N264) );
  OA22X1 U686 ( .IN1(n776), .IN2(n487), .IN3(n806), .IN4(n489), .Q(n413) );
  OA22X1 U687 ( .IN1(n808), .IN2(n493), .IN3(n802), .IN4(n485), .Q(n412) );
  INVX0 U688 ( .INP(n483), .ZN(n414) );
  NAND4X0 U689 ( .IN1(n413), .IN2(n412), .IN3(n411), .IN4(n410), .QN(N265) );
  OA22X1 U690 ( .IN1(n786), .IN2(n489), .IN3(n806), .IN4(n493), .Q(n418) );
  OA22X1 U691 ( .IN1(n777), .IN2(n487), .IN3(n776), .IN4(n491), .Q(n417) );
  OA22X1 U692 ( .IN1(n808), .IN2(n485), .IN3(n810), .IN4(n496), .Q(n416) );
  NAND4X0 U693 ( .IN1(n418), .IN2(n417), .IN3(n416), .IN4(n415), .QN(N266) );
  NOR4X0 U694 ( .IN1(n421), .IN2(n420), .IN3(n419), .IN4(N258), .QN(n558) );
  OA22X1 U695 ( .IN1(n808), .IN2(n483), .IN3(n806), .IN4(n485), .Q(n425) );
  OA22X1 U696 ( .IN1(n769), .IN2(n487), .IN3(n776), .IN4(n489), .Q(n424) );
  OA22X1 U697 ( .IN1(n777), .IN2(n491), .IN3(n786), .IN4(n493), .Q(n423) );
  OA22X1 U698 ( .IN1(n802), .IN2(n496), .IN3(n810), .IN4(n825), .Q(n422) );
  NAND4X0 U699 ( .IN1(n425), .IN2(n424), .IN3(n423), .IN4(n422), .QN(N267) );
  OA22X1 U700 ( .IN1(n786), .IN2(n485), .IN3(n806), .IN4(n483), .Q(n429) );
  OA22X1 U701 ( .IN1(n761), .IN2(n487), .IN3(n777), .IN4(n489), .Q(n428) );
  OA22X1 U702 ( .IN1(n769), .IN2(n491), .IN3(n776), .IN4(n493), .Q(n427) );
  OA22X1 U703 ( .IN1(n808), .IN2(n496), .IN3(n802), .IN4(n825), .Q(n426) );
  NAND4X0 U704 ( .IN1(n429), .IN2(n428), .IN3(n427), .IN4(n426), .QN(N268) );
  OA22X1 U705 ( .IN1(n776), .IN2(n485), .IN3(n786), .IN4(n483), .Q(n433) );
  OA22X1 U706 ( .IN1(n753), .IN2(n487), .IN3(n769), .IN4(n489), .Q(n432) );
  OA22X1 U707 ( .IN1(n761), .IN2(n491), .IN3(n777), .IN4(n493), .Q(n431) );
  OA22X1 U708 ( .IN1(n808), .IN2(n825), .IN3(n806), .IN4(n496), .Q(n430) );
  NAND4X0 U709 ( .IN1(n433), .IN2(n432), .IN3(n431), .IN4(n430), .QN(N269) );
  OA22X1 U710 ( .IN1(n777), .IN2(n485), .IN3(n776), .IN4(n483), .Q(n437) );
  OA22X1 U711 ( .IN1(n761), .IN2(n489), .IN3(n745), .IN4(n487), .Q(n436) );
  OA22X1 U712 ( .IN1(n753), .IN2(n491), .IN3(n769), .IN4(n493), .Q(n435) );
  OA22X1 U713 ( .IN1(n786), .IN2(n496), .IN3(n806), .IN4(n825), .Q(n434) );
  NAND4X0 U714 ( .IN1(n437), .IN2(n436), .IN3(n435), .IN4(n434), .QN(N270) );
  OA22X1 U715 ( .IN1(n769), .IN2(n485), .IN3(n777), .IN4(n483), .Q(n441) );
  OA22X1 U716 ( .IN1(n737), .IN2(n487), .IN3(n753), .IN4(n489), .Q(n440) );
  OA22X1 U717 ( .IN1(n761), .IN2(n493), .IN3(n745), .IN4(n491), .Q(n439) );
  OA22X1 U718 ( .IN1(n776), .IN2(n496), .IN3(n786), .IN4(n825), .Q(n438) );
  NAND4X0 U719 ( .IN1(n441), .IN2(n440), .IN3(n439), .IN4(n438), .QN(N271) );
  OA22X1 U720 ( .IN1(n761), .IN2(n485), .IN3(n769), .IN4(n483), .Q(n446) );
  OA22X1 U721 ( .IN1(n729), .IN2(n487), .IN3(n745), .IN4(n489), .Q(n445) );
  OA22X1 U722 ( .IN1(n737), .IN2(n491), .IN3(n753), .IN4(n493), .Q(n444) );
  OA22X1 U723 ( .IN1(n777), .IN2(n496), .IN3(n776), .IN4(n825), .Q(n443) );
  NAND4X0 U724 ( .IN1(n446), .IN2(n445), .IN3(n444), .IN4(n443), .QN(N272) );
  OA22X1 U725 ( .IN1(n761), .IN2(n483), .IN3(n753), .IN4(n485), .Q(n451) );
  OA22X1 U726 ( .IN1(n737), .IN2(n489), .IN3(n718), .IN4(n487), .Q(n450) );
  OA22X1 U727 ( .IN1(n729), .IN2(n491), .IN3(n745), .IN4(n493), .Q(n449) );
  OA22X1 U728 ( .IN1(n769), .IN2(n496), .IN3(n777), .IN4(n825), .Q(n448) );
  NAND4X0 U729 ( .IN1(n451), .IN2(n450), .IN3(n449), .IN4(n448), .QN(N273) );
  OA22X1 U730 ( .IN1(n745), .IN2(n485), .IN3(n753), .IN4(n483), .Q(n455) );
  INVX0 U731 ( .INP(n501), .ZN(n495) );
  OA22X1 U732 ( .IN1(n495), .IN2(n487), .IN3(n729), .IN4(n489), .Q(n454) );
  OA22X1 U733 ( .IN1(n737), .IN2(n493), .IN3(n718), .IN4(n491), .Q(n453) );
  OA22X1 U734 ( .IN1(n761), .IN2(n496), .IN3(n769), .IN4(n825), .Q(n452) );
  NAND4X0 U735 ( .IN1(n455), .IN2(n454), .IN3(n453), .IN4(n452), .QN(N274) );
  OA22X1 U736 ( .IN1(n737), .IN2(n485), .IN3(n745), .IN4(n483), .Q(n460) );
  OA22X1 U737 ( .IN1(n560), .IN2(n487), .IN3(n718), .IN4(n489), .Q(n459) );
  OA22X1 U738 ( .IN1(n495), .IN2(n491), .IN3(n729), .IN4(n493), .Q(n458) );
  OA22X1 U739 ( .IN1(n761), .IN2(n825), .IN3(n753), .IN4(n496), .Q(n457) );
  NAND4X0 U740 ( .IN1(n460), .IN2(n459), .IN3(n458), .IN4(n457), .QN(N275) );
  OA22X1 U741 ( .IN1(n729), .IN2(n485), .IN3(n737), .IN4(n483), .Q(n464) );
  OA22X1 U742 ( .IN1(n495), .IN2(n489), .IN3(n484), .IN4(n487), .Q(n463) );
  OA22X1 U743 ( .IN1(n560), .IN2(n491), .IN3(n718), .IN4(n493), .Q(n462) );
  OA22X1 U744 ( .IN1(n745), .IN2(n496), .IN3(n753), .IN4(n825), .Q(n461) );
  NAND4X0 U745 ( .IN1(n464), .IN2(n463), .IN3(n462), .IN4(n461), .QN(N276) );
  OA22X1 U746 ( .IN1(n729), .IN2(n483), .IN3(n718), .IN4(n485), .Q(n469) );
  INVX0 U747 ( .INP(n465), .ZN(n486) );
  OA22X1 U748 ( .IN1(n560), .IN2(n489), .IN3(n486), .IN4(n487), .Q(n468) );
  OA22X1 U749 ( .IN1(n495), .IN2(n493), .IN3(n484), .IN4(n491), .Q(n467) );
  OA22X1 U750 ( .IN1(n737), .IN2(n496), .IN3(n745), .IN4(n825), .Q(n466) );
  NAND4X0 U751 ( .IN1(n469), .IN2(n468), .IN3(n467), .IN4(n466), .QN(N277) );
  OA22X1 U752 ( .IN1(n495), .IN2(n485), .IN3(n718), .IN4(n483), .Q(n473) );
  OA22X1 U753 ( .IN1(n494), .IN2(n487), .IN3(n484), .IN4(n489), .Q(n472) );
  OA22X1 U754 ( .IN1(n560), .IN2(n493), .IN3(n486), .IN4(n491), .Q(n471) );
  OA22X1 U755 ( .IN1(n729), .IN2(n496), .IN3(n737), .IN4(n825), .Q(n470) );
  NAND4X0 U756 ( .IN1(n473), .IN2(n472), .IN3(n471), .IN4(n470), .QN(N278) );
  OA22X1 U757 ( .IN1(n560), .IN2(n485), .IN3(n495), .IN4(n483), .Q(n478) );
  INVX0 U758 ( .INP(n474), .ZN(n490) );
  OA22X1 U759 ( .IN1(n486), .IN2(n489), .IN3(n490), .IN4(n487), .Q(n477) );
  OA22X1 U760 ( .IN1(n494), .IN2(n491), .IN3(n484), .IN4(n493), .Q(n476) );
  OA22X1 U761 ( .IN1(n729), .IN2(n825), .IN3(n718), .IN4(n496), .Q(n475) );
  NAND4X0 U762 ( .IN1(n478), .IN2(n477), .IN3(n476), .IN4(n475), .QN(N279) );
  OA22X1 U763 ( .IN1(n560), .IN2(n483), .IN3(n484), .IN4(n485), .Q(n482) );
  OA22X1 U764 ( .IN1(n494), .IN2(n489), .IN3(n492), .IN4(n487), .Q(n481) );
  OA22X1 U765 ( .IN1(n486), .IN2(n493), .IN3(n490), .IN4(n491), .Q(n480) );
  OA22X1 U766 ( .IN1(n495), .IN2(n496), .IN3(n718), .IN4(n825), .Q(n479) );
  NAND4X0 U767 ( .IN1(n482), .IN2(n481), .IN3(n480), .IN4(n479), .QN(N280) );
  OA22X1 U768 ( .IN1(n486), .IN2(n485), .IN3(n484), .IN4(n483), .Q(n500) );
  OA22X1 U769 ( .IN1(n490), .IN2(n489), .IN3(n488), .IN4(n487), .Q(n499) );
  OA22X1 U770 ( .IN1(n494), .IN2(n493), .IN3(n492), .IN4(n491), .Q(n498) );
  OA22X1 U771 ( .IN1(n560), .IN2(n496), .IN3(n495), .IN4(n825), .Q(n497) );
  NAND4X0 U772 ( .IN1(n500), .IN2(n499), .IN3(n498), .IN4(n497), .QN(N281) );
  NAND3X0 U773 ( .IN1(n501), .IN2(n514), .IN3(n560), .QN(n717) );
  AO22X1 U774 ( .IN1(n512), .IN2(add_result[12]), .IN3(n510), .IN4(
        sub_result[12]), .Q(n502) );
  INVX0 U775 ( .INP(n717), .ZN(n508) );
  NOR3X0 U776 ( .IN1(n503), .IN2(add_result[14]), .IN3(add_result[15]), .QN(
        n505) );
  NOR3X0 U777 ( .IN1(sub_result[14]), .IN2(sub_result[15]), .IN3(n21), .QN(
        n504) );
  AO22X1 U778 ( .IN1(n505), .IN2(add_result[13]), .IN3(n504), .IN4(
        sub_result[13]), .Q(n506) );
  NOR2X0 U779 ( .IN1(n508), .IN2(n507), .QN(N308) );
  INVX0 U780 ( .INP(add_result[12]), .ZN(n511) );
  INVX0 U781 ( .INP(sub_result[12]), .ZN(n509) );
  AO22X1 U782 ( .IN1(n512), .IN2(n511), .IN3(n510), .IN4(n509), .Q(n513) );
  NAND3X0 U783 ( .IN1(n514), .IN2(n724), .IN3(n513), .QN(n811) );
  NAND4X0 U784 ( .IN1(N308), .IN2(n811), .IN3(n794), .IN4(n785), .QN(n778) );
  NAND4X0 U785 ( .IN1(n794), .IN2(n717), .IN3(n723), .IN4(n778), .QN(N306) );
  NAND4X0 U786 ( .IN1(n785), .IN2(n716), .IN3(n723), .IN4(n778), .QN(N307) );
  AO22X1 U787 ( .IN1(n708), .IN2(exponent_factor_12[0]), .IN3(n821), .IN4(
        exponent_factor_21[0]), .Q(N34) );
  NAND3X0 U788 ( .IN1(n806), .IN2(n524), .IN3(n796), .QN(n537) );
  NAND3X0 U789 ( .IN1(n776), .IN2(n516), .IN3(n797), .QN(n532) );
  NAND3X0 U790 ( .IN1(n769), .IN2(n517), .IN3(n764), .QN(n533) );
  NAND3X0 U791 ( .IN1(n808), .IN2(n802), .IN3(n806), .QN(n515) );
  AND2X1 U792 ( .IN1(n532), .IN2(n534), .Q(n519) );
  NAND4X0 U793 ( .IN1(n521), .IN2(n519), .IN3(n533), .IN4(n535), .QN(n520) );
  NAND4X0 U794 ( .IN1(n537), .IN2(n532), .IN3(n533), .IN4(n520), .QN(N346) );
  NAND3X0 U795 ( .IN1(n519), .IN2(n536), .IN3(n520), .QN(N347) );
  NOR2X0 U796 ( .IN1(n810), .IN2(n535), .QN(N349) );
  AO22X1 U797 ( .IN1(n708), .IN2(exponent_factor_12[1]), .IN3(n821), .IN4(
        exponent_factor_21[1]), .Q(N35) );
  OAI22X1 U798 ( .IN1(n802), .IN2(n535), .IN3(n810), .IN4(n533), .QN(N350) );
  OAI222X1 U799 ( .IN1(n534), .IN2(n810), .IN3(n533), .IN4(n802), .IN5(n535), 
        .IN6(n808), .QN(N351) );
  OA22X1 U800 ( .IN1(n808), .IN2(n533), .IN3(n806), .IN4(n535), .Q(n523) );
  OA22X1 U801 ( .IN1(n802), .IN2(n534), .IN3(n810), .IN4(n532), .Q(n522) );
  OA22X1 U802 ( .IN1(n786), .IN2(n535), .IN3(n806), .IN4(n533), .Q(n527) );
  OA22X1 U803 ( .IN1(n808), .IN2(n534), .IN3(n802), .IN4(n532), .Q(n526) );
  AND2X1 U804 ( .IN1(n524), .IN2(n788), .Q(n538) );
  NAND3X0 U805 ( .IN1(n527), .IN2(n526), .IN3(n525), .QN(N353) );
  OA22X1 U806 ( .IN1(n776), .IN2(n535), .IN3(n786), .IN4(n533), .Q(n531) );
  OA22X1 U807 ( .IN1(n808), .IN2(n532), .IN3(n810), .IN4(n537), .Q(n530) );
  OR2X1 U808 ( .IN1(n534), .IN2(n806), .Q(n528) );
  NAND4X0 U809 ( .IN1(n531), .IN2(n530), .IN3(n529), .IN4(n528), .QN(N354) );
  OA22X1 U810 ( .IN1(n776), .IN2(n533), .IN3(n806), .IN4(n532), .Q(n542) );
  OA22X1 U811 ( .IN1(n777), .IN2(n535), .IN3(n786), .IN4(n534), .Q(n541) );
  OA22X1 U812 ( .IN1(n802), .IN2(n537), .IN3(n810), .IN4(n536), .Q(n540) );
  NAND4X0 U813 ( .IN1(n542), .IN2(n541), .IN3(n540), .IN4(n539), .QN(N355) );
  AO22X1 U814 ( .IN1(n708), .IN2(exponent_factor_12[2]), .IN3(n821), .IN4(
        exponent_factor_21[2]), .Q(N36) );
  AO22X1 U815 ( .IN1(n708), .IN2(exponent_factor_12[3]), .IN3(n821), .IN4(
        exponent_factor_21[3]), .Q(N37) );
  AO22X1 U816 ( .IN1(n708), .IN2(exponent_factor_12[4]), .IN3(n821), .IN4(
        exponent_factor_21[4]), .Q(N38) );
  NAND4X0 U817 ( .IN1(n590), .IN2(n578), .IN3(n584), .IN4(n543), .QN(n544) );
  NOR4X0 U818 ( .IN1(input_factor_01[30]), .IN2(input_factor_01[23]), .IN3(
        n545), .IN4(n544), .QN(n554) );
  NOR4X0 U819 ( .IN1(input_factor_01[22]), .IN2(input_factor_01[21]), .IN3(
        input_factor_01[20]), .IN4(input_factor_01[17]), .QN(n553) );
  NOR4X0 U820 ( .IN1(input_factor_01[31]), .IN2(input_factor_01[25]), .IN3(
        input_factor_01[29]), .IN4(input_factor_01[16]), .QN(n552) );
  NAND4X0 U821 ( .IN1(n628), .IN2(n624), .IN3(n620), .IN4(n616), .QN(n550) );
  NAND4X0 U822 ( .IN1(n612), .IN2(n608), .IN3(n546), .IN4(n604), .QN(n549) );
  NAND4X0 U823 ( .IN1(n672), .IN2(n666), .IN3(n660), .IN4(n654), .QN(n548) );
  NAND4X0 U824 ( .IN1(n648), .IN2(n642), .IN3(n636), .IN4(n632), .QN(n547) );
  NOR4X0 U825 ( .IN1(n550), .IN2(n549), .IN3(n548), .IN4(n547), .QN(n551) );
  AOI22X1 U826 ( .IN1(input_factor_02[23]), .IN2(n22), .IN3(n710), .IN4(
        input_factor_01[23]), .QN(n569) );
  INVX0 U827 ( .INP(n778), .ZN(n555) );
  OA21X1 U828 ( .IN1(n761), .IN2(n556), .IN3(n555), .Q(n562) );
  NAND3X0 U829 ( .IN1(n557), .IN2(n701), .IN3(n702), .QN(n564) );
  OA21X1 U830 ( .IN1(n560), .IN2(n559), .IN3(n558), .Q(n561) );
  AOI22X1 U831 ( .IN1(n712), .IN2(add_output_exponent_w3[0]), .IN3(n711), 
        .IN4(add_output_exponent_w2[0]), .QN(n568) );
  INVX0 U832 ( .INP(n564), .ZN(n563) );
  AND4X1 U833 ( .IN1(n565), .IN2(n563), .IN3(n562), .IN4(n561), .Q(n714) );
  NAND4X0 U834 ( .IN1(n569), .IN2(n568), .IN3(n567), .IN4(n566), .QN(N380) );
  AOI22X1 U835 ( .IN1(input_factor_02[24]), .IN2(n22), .IN3(n710), .IN4(
        input_factor_01[24]), .QN(n573) );
  AOI22X1 U836 ( .IN1(n712), .IN2(add_output_exponent_w3[1]), .IN3(n711), 
        .IN4(add_output_exponent_w2[1]), .QN(n572) );
  NAND4X0 U837 ( .IN1(n573), .IN2(n572), .IN3(n571), .IN4(n570), .QN(N381) );
  AOI22X1 U838 ( .IN1(input_factor_02[25]), .IN2(n22), .IN3(n710), .IN4(
        input_factor_01[25]), .QN(n577) );
  AOI22X1 U839 ( .IN1(n712), .IN2(add_output_exponent_w3[2]), .IN3(n711), 
        .IN4(add_output_exponent_w2[2]), .QN(n576) );
  NAND4X0 U840 ( .IN1(n577), .IN2(n576), .IN3(n575), .IN4(n574), .QN(N382) );
  OA22X1 U841 ( .IN1(n579), .IN2(n702), .IN3(n701), .IN4(n578), .Q(n583) );
  AOI22X1 U842 ( .IN1(n712), .IN2(add_output_exponent_w3[3]), .IN3(n711), 
        .IN4(add_output_exponent_w2[3]), .QN(n582) );
  NAND4X0 U843 ( .IN1(n583), .IN2(n582), .IN3(n581), .IN4(n580), .QN(N383) );
  OA22X1 U844 ( .IN1(n585), .IN2(n702), .IN3(n701), .IN4(n584), .Q(n589) );
  AOI22X1 U845 ( .IN1(n712), .IN2(add_output_exponent_w3[4]), .IN3(n711), 
        .IN4(add_output_exponent_w2[4]), .QN(n588) );
  NAND4X0 U846 ( .IN1(n589), .IN2(n588), .IN3(n587), .IN4(n586), .QN(N384) );
  OA22X1 U847 ( .IN1(n591), .IN2(n702), .IN3(n701), .IN4(n590), .Q(n595) );
  AOI22X1 U848 ( .IN1(n712), .IN2(add_output_exponent_w3[5]), .IN3(n711), 
        .IN4(add_output_exponent_w2[5]), .QN(n594) );
  NAND4X0 U849 ( .IN1(n595), .IN2(n594), .IN3(n593), .IN4(n592), .QN(N385) );
  OA22X1 U850 ( .IN1(n597), .IN2(n702), .IN3(n701), .IN4(n596), .Q(n601) );
  AOI22X1 U851 ( .IN1(n712), .IN2(add_output_exponent_w3[6]), .IN3(n711), 
        .IN4(add_output_exponent_w2[6]), .QN(n600) );
  NAND4X0 U852 ( .IN1(n601), .IN2(n600), .IN3(n599), .IN4(n598), .QN(N386) );
  AO22X1 U854 ( .IN1(n710), .IN2(input_factor_01[30]), .IN3(n709), .IN4(
        add_output_exponent_w1[7]), .Q(n603) );
  AO22X1 U855 ( .IN1(n712), .IN2(add_output_exponent_w3[7]), .IN3(n711), .IN4(
        add_output_exponent_w2[7]), .Q(n602) );
  AO222X1 U856 ( .IN1(input_factor_02[0]), .IN2(n22), .IN3(input_factor_01[0]), 
        .IN4(n710), .IN5(n709), .IN6(pre_sig_res_01[0]), .Q(N388) );
  AOI22X1 U857 ( .IN1(n711), .IN2(pre_sig_res_02[1]), .IN3(n709), .IN4(
        pre_sig_res_01[1]), .QN(n607) );
  OA22X1 U858 ( .IN1(n605), .IN2(n702), .IN3(n701), .IN4(n604), .Q(n606) );
  AO22X1 U859 ( .IN1(n708), .IN2(exponent_factor_12[5]), .IN3(n821), .IN4(
        exponent_factor_21[5]), .Q(N39) );
  AOI22X1 U860 ( .IN1(n711), .IN2(pre_sig_res_02[2]), .IN3(n709), .IN4(
        pre_sig_res_01[2]), .QN(n611) );
  OA22X1 U861 ( .IN1(n609), .IN2(n702), .IN3(n701), .IN4(n608), .Q(n610) );
  AOI22X1 U862 ( .IN1(n711), .IN2(pre_sig_res_02[3]), .IN3(n709), .IN4(
        pre_sig_res_01[3]), .QN(n615) );
  OA22X1 U863 ( .IN1(n613), .IN2(n702), .IN3(n701), .IN4(n612), .Q(n614) );
  AOI22X1 U864 ( .IN1(n711), .IN2(pre_sig_res_02[4]), .IN3(n709), .IN4(
        pre_sig_res_01[4]), .QN(n619) );
  OA22X1 U865 ( .IN1(n617), .IN2(n702), .IN3(n701), .IN4(n616), .Q(n618) );
  AOI22X1 U866 ( .IN1(n711), .IN2(pre_sig_res_02[5]), .IN3(n709), .IN4(
        pre_sig_res_01[5]), .QN(n623) );
  OA22X1 U867 ( .IN1(n621), .IN2(n702), .IN3(n701), .IN4(n620), .Q(n622) );
  AOI22X1 U868 ( .IN1(n711), .IN2(pre_sig_res_02[6]), .IN3(n709), .IN4(
        pre_sig_res_01[6]), .QN(n627) );
  OA22X1 U869 ( .IN1(n625), .IN2(n702), .IN3(n701), .IN4(n624), .Q(n626) );
  AOI22X1 U870 ( .IN1(n711), .IN2(pre_sig_res_02[7]), .IN3(n709), .IN4(
        pre_sig_res_01[7]), .QN(n631) );
  OA22X1 U871 ( .IN1(n629), .IN2(n702), .IN3(n701), .IN4(n628), .Q(n630) );
  AOI22X1 U872 ( .IN1(n711), .IN2(pre_sig_res_02[8]), .IN3(n709), .IN4(
        pre_sig_res_01[8]), .QN(n635) );
  OA22X1 U873 ( .IN1(n633), .IN2(n702), .IN3(n701), .IN4(n632), .Q(n634) );
  OA22X1 U874 ( .IN1(n637), .IN2(n702), .IN3(n701), .IN4(n636), .Q(n641) );
  NAND4X0 U875 ( .IN1(n641), .IN2(n640), .IN3(n639), .IN4(n638), .QN(N397) );
  OA22X1 U876 ( .IN1(n643), .IN2(n702), .IN3(n701), .IN4(n642), .Q(n647) );
  NAND4X0 U877 ( .IN1(n647), .IN2(n646), .IN3(n645), .IN4(n644), .QN(N398) );
  OA22X1 U878 ( .IN1(n649), .IN2(n702), .IN3(n701), .IN4(n648), .Q(n653) );
  NAND4X0 U879 ( .IN1(n653), .IN2(n652), .IN3(n651), .IN4(n650), .QN(N399) );
  AO22X1 U880 ( .IN1(n708), .IN2(exponent_factor_12[6]), .IN3(n821), .IN4(
        exponent_factor_21[6]), .Q(N40) );
  OA22X1 U881 ( .IN1(n655), .IN2(n702), .IN3(n701), .IN4(n654), .Q(n659) );
  NAND4X0 U882 ( .IN1(n659), .IN2(n658), .IN3(n657), .IN4(n656), .QN(N400) );
  OA22X1 U883 ( .IN1(n661), .IN2(n702), .IN3(n701), .IN4(n660), .Q(n665) );
  NAND4X0 U884 ( .IN1(n665), .IN2(n664), .IN3(n663), .IN4(n662), .QN(N401) );
  OA22X1 U885 ( .IN1(n667), .IN2(n702), .IN3(n701), .IN4(n666), .Q(n671) );
  NAND4X0 U886 ( .IN1(n671), .IN2(n670), .IN3(n669), .IN4(n668), .QN(N402) );
  OA22X1 U887 ( .IN1(n673), .IN2(n702), .IN3(n701), .IN4(n672), .Q(n677) );
  NAND4X0 U888 ( .IN1(n677), .IN2(n676), .IN3(n675), .IN4(n674), .QN(N403) );
  OA22X1 U889 ( .IN1(n679), .IN2(n702), .IN3(n701), .IN4(n678), .Q(n683) );
  AOI22X1 U890 ( .IN1(n712), .IN2(pre_sig_res_03[16]), .IN3(n711), .IN4(
        pre_sig_res_02[16]), .QN(n682) );
  NAND4X0 U891 ( .IN1(n683), .IN2(n682), .IN3(n681), .IN4(n680), .QN(N404) );
  OA22X1 U892 ( .IN1(n685), .IN2(n702), .IN3(n701), .IN4(n684), .Q(n689) );
  AOI22X1 U893 ( .IN1(n712), .IN2(pre_sig_res_03[17]), .IN3(n711), .IN4(
        pre_sig_res_02[17]), .QN(n688) );
  NAND4X0 U894 ( .IN1(n689), .IN2(n688), .IN3(n687), .IN4(n686), .QN(N405) );
  AO22X1 U895 ( .IN1(n710), .IN2(input_factor_01[18]), .IN3(n709), .IN4(
        pre_sig_res_01[18]), .Q(n691) );
  AO22X1 U896 ( .IN1(n712), .IN2(pre_sig_res_03[18]), .IN3(n711), .IN4(
        pre_sig_res_02[18]), .Q(n690) );
  AO22X1 U897 ( .IN1(n710), .IN2(input_factor_01[19]), .IN3(n709), .IN4(
        pre_sig_res_01[19]), .Q(n693) );
  AO22X1 U898 ( .IN1(n712), .IN2(pre_sig_res_03[19]), .IN3(n711), .IN4(
        pre_sig_res_02[19]), .Q(n692) );
  OA22X1 U899 ( .IN1(n695), .IN2(n702), .IN3(n701), .IN4(n694), .Q(n699) );
  AOI22X1 U900 ( .IN1(n712), .IN2(pre_sig_res_03[20]), .IN3(n711), .IN4(
        pre_sig_res_02[20]), .QN(n698) );
  NAND4X0 U901 ( .IN1(n699), .IN2(n698), .IN3(n697), .IN4(n696), .QN(N408) );
  OA22X1 U902 ( .IN1(n703), .IN2(n702), .IN3(n701), .IN4(n700), .Q(n707) );
  AOI22X1 U903 ( .IN1(n712), .IN2(pre_sig_res_03[21]), .IN3(n711), .IN4(
        pre_sig_res_02[21]), .QN(n706) );
  NAND4X0 U904 ( .IN1(n707), .IN2(n706), .IN3(n705), .IN4(n704), .QN(N409) );
  AO22X1 U905 ( .IN1(n708), .IN2(exponent_factor_12[7]), .IN3(n821), .IN4(
        exponent_factor_21[7]), .Q(N41) );
  AO22X1 U906 ( .IN1(n710), .IN2(input_factor_01[22]), .IN3(n709), .IN4(
        pre_sig_res_01[22]), .Q(n715) );
  AO22X1 U907 ( .IN1(n712), .IN2(pre_sig_res_03[22]), .IN3(n711), .IN4(
        pre_sig_res_02[22]), .Q(n713) );
  NOR2X0 U908 ( .IN1(n848), .IN2(n716), .QN(n817) );
  NOR2X0 U909 ( .IN1(n717), .IN2(n848), .QN(n819) );
  OA22X1 U910 ( .IN1(n729), .IN2(n807), .IN3(n718), .IN4(n805), .Q(n728) );
  OA22X1 U911 ( .IN1(n745), .IN2(n811), .IN3(n769), .IN4(n778), .Q(n722) );
  INVX0 U912 ( .INP(rst_n), .ZN(n820) );
  NAND3X0 U913 ( .IN1(n720), .IN2(n740), .IN3(n719), .QN(n721) );
  OA22X1 U914 ( .IN1(n848), .IN2(n722), .IN3(n820), .IN4(n721), .Q(n727) );
  NAND4X0 U915 ( .IN1(n728), .IN2(n727), .IN3(n726), .IN4(n725), .QN(n847) );
  OA22X1 U916 ( .IN1(n729), .IN2(n805), .IN3(n737), .IN4(n807), .Q(n736) );
  OA22X1 U917 ( .IN1(n769), .IN2(n785), .IN3(n777), .IN4(n778), .Q(n731) );
  OA22X1 U918 ( .IN1(n761), .IN2(n794), .IN3(n753), .IN4(n811), .Q(n730) );
  AO21X1 U919 ( .IN1(n731), .IN2(n730), .IN3(n848), .Q(n735) );
  NAND4X0 U920 ( .IN1(n736), .IN2(n735), .IN3(n734), .IN4(n733), .QN(n846) );
  OA22X1 U921 ( .IN1(n737), .IN2(n805), .IN3(n745), .IN4(n807), .Q(n744) );
  OA22X1 U922 ( .IN1(n777), .IN2(n785), .IN3(n776), .IN4(n778), .Q(n739) );
  OA22X1 U923 ( .IN1(n761), .IN2(n811), .IN3(n769), .IN4(n794), .Q(n738) );
  AO21X1 U924 ( .IN1(n739), .IN2(n738), .IN3(n848), .Q(n743) );
  NAND4X0 U925 ( .IN1(n744), .IN2(n743), .IN3(n742), .IN4(n741), .QN(n845) );
  OA22X1 U926 ( .IN1(n745), .IN2(n805), .IN3(n753), .IN4(n807), .Q(n752) );
  OA22X1 U927 ( .IN1(n776), .IN2(n785), .IN3(n786), .IN4(n778), .Q(n747) );
  OA22X1 U928 ( .IN1(n769), .IN2(n811), .IN3(n777), .IN4(n794), .Q(n746) );
  AO21X1 U929 ( .IN1(n747), .IN2(n746), .IN3(n848), .Q(n751) );
  NAND4X0 U930 ( .IN1(n752), .IN2(n751), .IN3(n750), .IN4(n749), .QN(n844) );
  OA22X1 U931 ( .IN1(n761), .IN2(n807), .IN3(n753), .IN4(n805), .Q(n760) );
  OA22X1 U932 ( .IN1(n786), .IN2(n785), .IN3(n806), .IN4(n778), .Q(n755) );
  OA22X1 U933 ( .IN1(n777), .IN2(n811), .IN3(n776), .IN4(n794), .Q(n754) );
  AO21X1 U934 ( .IN1(n755), .IN2(n754), .IN3(n848), .Q(n759) );
  NAND4X0 U935 ( .IN1(n760), .IN2(n759), .IN3(n758), .IN4(n757), .QN(n843) );
  OA22X1 U936 ( .IN1(n761), .IN2(n805), .IN3(n769), .IN4(n807), .Q(n768) );
  OA22X1 U937 ( .IN1(n808), .IN2(n778), .IN3(n806), .IN4(n785), .Q(n763) );
  OA22X1 U938 ( .IN1(n776), .IN2(n811), .IN3(n786), .IN4(n794), .Q(n762) );
  AO21X1 U939 ( .IN1(n763), .IN2(n762), .IN3(n848), .Q(n767) );
  NAND4X0 U940 ( .IN1(n768), .IN2(n767), .IN3(n766), .IN4(n765), .QN(n842) );
  OA22X1 U941 ( .IN1(n769), .IN2(n805), .IN3(n777), .IN4(n807), .Q(n775) );
  OA22X1 U942 ( .IN1(n808), .IN2(n785), .IN3(n802), .IN4(n778), .Q(n771) );
  OA22X1 U943 ( .IN1(n786), .IN2(n811), .IN3(n806), .IN4(n794), .Q(n770) );
  AO21X1 U944 ( .IN1(n771), .IN2(n770), .IN3(n848), .Q(n774) );
  NAND4X0 U945 ( .IN1(n775), .IN2(n774), .IN3(n773), .IN4(n772), .QN(n841) );
  OA22X1 U946 ( .IN1(n777), .IN2(n805), .IN3(n776), .IN4(n807), .Q(n784) );
  OA22X1 U947 ( .IN1(n802), .IN2(n785), .IN3(n810), .IN4(n778), .Q(n780) );
  OA22X1 U948 ( .IN1(n808), .IN2(n794), .IN3(n806), .IN4(n811), .Q(n779) );
  AO21X1 U949 ( .IN1(n780), .IN2(n779), .IN3(n848), .Q(n783) );
  NAND4X0 U950 ( .IN1(n784), .IN2(n783), .IN3(n782), .IN4(n781), .QN(n840) );
  OA222X1 U951 ( .IN1(n811), .IN2(n808), .IN3(n785), .IN4(n810), .IN5(n794), 
        .IN6(n802), .Q(n787) );
  OA22X1 U952 ( .IN1(n848), .IN2(n787), .IN3(n786), .IN4(n807), .Q(n793) );
  NAND4X0 U953 ( .IN1(n793), .IN2(n792), .IN3(n791), .IN4(n790), .QN(n839) );
  OA22X1 U954 ( .IN1(n802), .IN2(n811), .IN3(n810), .IN4(n794), .Q(n795) );
  OA22X1 U955 ( .IN1(n806), .IN2(n807), .IN3(n795), .IN4(n820), .Q(n801) );
  NAND4X0 U956 ( .IN1(n801), .IN2(n800), .IN3(n799), .IN4(n798), .QN(n838) );
  AOI22X1 U957 ( .IN1(pre_sig_res_03[11]), .IN2(n820), .IN3(n809), .IN4(n818), 
        .QN(n804) );
  OA22X1 U958 ( .IN1(n808), .IN2(n805), .IN3(n802), .IN4(n807), .Q(n803) );
  OA22X1 U959 ( .IN1(n808), .IN2(n807), .IN3(n806), .IN4(n805), .Q(n815) );
  OR3X1 U960 ( .IN1(n811), .IN2(n820), .IN3(n810), .Q(n813) );
  NAND4X0 U961 ( .IN1(n815), .IN2(n814), .IN3(n813), .IN4(n812), .QN(n836) );
  AO222X1 U962 ( .IN1(n818), .IN2(n817), .IN3(n816), .IN4(n819), .IN5(n820), 
        .IN6(pre_sig_res_03[10]), .Q(n835) );
  AO22X1 U963 ( .IN1(pre_sig_res_03[9]), .IN2(n820), .IN3(n819), .IN4(n818), 
        .Q(n834) );
  AND2X1 U964 ( .IN1(n821), .IN2(rst_n), .Q(n823) );
  AO222X1 U965 ( .IN1(input_factor_02[23]), .IN2(n823), .IN3(
        input_factor_01[23]), .IN4(n822), .IN5(larger_exponent[0]), .IN6(n848), 
        .Q(n833) );
  AO222X1 U966 ( .IN1(input_factor_02[24]), .IN2(n823), .IN3(
        input_factor_01[24]), .IN4(n822), .IN5(n848), .IN6(larger_exponent[1]), 
        .Q(n832) );
  AO222X1 U967 ( .IN1(input_factor_02[25]), .IN2(n823), .IN3(
        input_factor_01[25]), .IN4(n822), .IN5(n848), .IN6(larger_exponent[2]), 
        .Q(n831) );
  AO222X1 U968 ( .IN1(input_factor_02[26]), .IN2(n823), .IN3(
        input_factor_01[26]), .IN4(n822), .IN5(n848), .IN6(larger_exponent[3]), 
        .Q(n830) );
  AO222X1 U969 ( .IN1(input_factor_02[27]), .IN2(n823), .IN3(
        input_factor_01[27]), .IN4(n822), .IN5(n848), .IN6(larger_exponent[4]), 
        .Q(n829) );
  AO222X1 U970 ( .IN1(input_factor_02[28]), .IN2(n823), .IN3(
        input_factor_01[28]), .IN4(n822), .IN5(n848), .IN6(larger_exponent[5]), 
        .Q(n828) );
  AO222X1 U971 ( .IN1(input_factor_02[29]), .IN2(n823), .IN3(
        input_factor_01[29]), .IN4(n822), .IN5(n848), .IN6(larger_exponent[6]), 
        .Q(n827) );
endmodule


module cla51squ_4 ( out, a, b );
  output [50:0] out;
  input [50:0] a;
  input [50:0] b;
  wire   intadd_4_CI, intadd_4_n24, intadd_4_n23, intadd_4_n22, intadd_4_n21,
         intadd_4_n20, intadd_4_n19, intadd_4_n18, intadd_4_n17, intadd_4_n16,
         intadd_4_n15, intadd_4_n14, intadd_4_n13, intadd_4_n12, intadd_4_n11,
         intadd_4_n10, intadd_4_n9, intadd_4_n8, intadd_4_n7, intadd_4_n6,
         intadd_4_n5, intadd_4_n4, intadd_4_n3, intadd_4_n2, intadd_4_n1, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14;

  FADDX1 intadd_4_U25 ( .A(b[23]), .B(a[23]), .CI(intadd_4_CI), .CO(
        intadd_4_n24), .S(out[23]) );
  FADDX1 intadd_4_U24 ( .A(b[24]), .B(a[24]), .CI(intadd_4_n24), .CO(
        intadd_4_n23), .S(out[24]) );
  FADDX1 intadd_4_U23 ( .A(b[25]), .B(a[25]), .CI(intadd_4_n23), .CO(
        intadd_4_n22), .S(out[25]) );
  FADDX1 intadd_4_U22 ( .A(b[26]), .B(a[26]), .CI(intadd_4_n22), .CO(
        intadd_4_n21), .S(out[26]) );
  FADDX1 intadd_4_U21 ( .A(b[27]), .B(a[27]), .CI(intadd_4_n21), .CO(
        intadd_4_n20), .S(out[27]) );
  FADDX1 intadd_4_U20 ( .A(b[28]), .B(a[28]), .CI(intadd_4_n20), .CO(
        intadd_4_n19), .S(out[28]) );
  FADDX1 intadd_4_U19 ( .A(b[29]), .B(a[29]), .CI(intadd_4_n19), .CO(
        intadd_4_n18), .S(out[29]) );
  FADDX1 intadd_4_U18 ( .A(b[30]), .B(a[30]), .CI(intadd_4_n18), .CO(
        intadd_4_n17), .S(out[30]) );
  FADDX1 intadd_4_U17 ( .A(b[31]), .B(a[31]), .CI(intadd_4_n17), .CO(
        intadd_4_n16), .S(out[31]) );
  FADDX1 intadd_4_U16 ( .A(b[32]), .B(a[32]), .CI(intadd_4_n16), .CO(
        intadd_4_n15), .S(out[32]) );
  FADDX1 intadd_4_U15 ( .A(b[33]), .B(a[33]), .CI(intadd_4_n15), .CO(
        intadd_4_n14), .S(out[33]) );
  FADDX1 intadd_4_U14 ( .A(b[34]), .B(a[34]), .CI(intadd_4_n14), .CO(
        intadd_4_n13), .S(out[34]) );
  FADDX1 intadd_4_U13 ( .A(b[35]), .B(a[35]), .CI(intadd_4_n13), .CO(
        intadd_4_n12), .S(out[35]) );
  FADDX1 intadd_4_U12 ( .A(b[36]), .B(a[36]), .CI(intadd_4_n12), .CO(
        intadd_4_n11), .S(out[36]) );
  FADDX1 intadd_4_U11 ( .A(b[37]), .B(a[37]), .CI(intadd_4_n11), .CO(
        intadd_4_n10), .S(out[37]) );
  FADDX1 intadd_4_U10 ( .A(b[38]), .B(a[38]), .CI(intadd_4_n10), .CO(
        intadd_4_n9), .S(out[38]) );
  FADDX1 intadd_4_U9 ( .A(b[39]), .B(a[39]), .CI(intadd_4_n9), .CO(intadd_4_n8), .S(out[39]) );
  FADDX1 intadd_4_U8 ( .A(b[40]), .B(a[40]), .CI(intadd_4_n8), .CO(intadd_4_n7), .S(out[40]) );
  FADDX1 intadd_4_U7 ( .A(b[41]), .B(a[41]), .CI(intadd_4_n7), .CO(intadd_4_n6), .S(out[41]) );
  FADDX1 intadd_4_U6 ( .A(b[42]), .B(a[42]), .CI(intadd_4_n6), .CO(intadd_4_n5), .S(out[42]) );
  FADDX1 intadd_4_U5 ( .A(b[43]), .B(a[43]), .CI(intadd_4_n5), .CO(intadd_4_n4), .S(out[43]) );
  FADDX1 intadd_4_U4 ( .A(b[44]), .B(a[44]), .CI(intadd_4_n4), .CO(intadd_4_n3), .S(out[44]) );
  FADDX1 intadd_4_U3 ( .A(b[45]), .B(a[45]), .CI(intadd_4_n3), .CO(intadd_4_n2), .S(out[45]) );
  FADDX1 intadd_4_U2 ( .A(b[46]), .B(a[46]), .CI(intadd_4_n2), .CO(intadd_4_n1), .S(out[46]) );
  OA21X1 U2 ( .IN1(b[9]), .IN2(a[9]), .IN3(a[8]), .Q(n1) );
  AO22X1 U3 ( .IN1(b[9]), .IN2(a[9]), .IN3(b[8]), .IN4(n1), .Q(n2) );
  AO222X1 U4 ( .IN1(b[10]), .IN2(a[10]), .IN3(b[10]), .IN4(n2), .IN5(a[10]), 
        .IN6(n2), .Q(n3) );
  AO222X1 U5 ( .IN1(b[11]), .IN2(a[11]), .IN3(b[11]), .IN4(n3), .IN5(a[11]), 
        .IN6(n3), .Q(n4) );
  AO222X1 U6 ( .IN1(b[12]), .IN2(a[12]), .IN3(b[12]), .IN4(n4), .IN5(a[12]), 
        .IN6(n4), .Q(n5) );
  AO222X1 U7 ( .IN1(b[13]), .IN2(a[13]), .IN3(b[13]), .IN4(n5), .IN5(a[13]), 
        .IN6(n5), .Q(n6) );
  AO222X1 U8 ( .IN1(b[14]), .IN2(a[14]), .IN3(b[14]), .IN4(n6), .IN5(a[14]), 
        .IN6(n6), .Q(n7) );
  AO222X1 U9 ( .IN1(b[15]), .IN2(a[15]), .IN3(b[15]), .IN4(n7), .IN5(a[15]), 
        .IN6(n7), .Q(n8) );
  AO222X1 U10 ( .IN1(b[16]), .IN2(a[16]), .IN3(b[16]), .IN4(n8), .IN5(a[16]), 
        .IN6(n8), .Q(n9) );
  AO222X1 U11 ( .IN1(b[17]), .IN2(a[17]), .IN3(b[17]), .IN4(n9), .IN5(a[17]), 
        .IN6(n9), .Q(n10) );
  AO222X1 U12 ( .IN1(b[18]), .IN2(a[18]), .IN3(b[18]), .IN4(n10), .IN5(a[18]), 
        .IN6(n10), .Q(n11) );
  AO222X1 U13 ( .IN1(b[19]), .IN2(a[19]), .IN3(b[19]), .IN4(n11), .IN5(a[19]), 
        .IN6(n11), .Q(n12) );
  AO222X1 U14 ( .IN1(b[20]), .IN2(a[20]), .IN3(b[20]), .IN4(n12), .IN5(a[20]), 
        .IN6(n12), .Q(n13) );
  AO222X1 U15 ( .IN1(b[21]), .IN2(a[21]), .IN3(b[21]), .IN4(n13), .IN5(a[21]), 
        .IN6(n13), .Q(n14) );
  AO222X1 U16 ( .IN1(b[22]), .IN2(a[22]), .IN3(b[22]), .IN4(n14), .IN5(a[22]), 
        .IN6(n14), .Q(intadd_4_CI) );
  XOR3X1 U17 ( .IN1(intadd_4_n1), .IN2(a[47]), .IN3(b[47]), .Q(out[47]) );
endmodule


module csa51squ_37 ( sumout, in1, in2, in3, cout_50_, cout_49_, cout_48_, 
        cout_47_, cout_46_, cout_44_, cout_42_, cout_40_, cout_38_, cout_36_, 
        cout_34_, cout_32_, cout_30_, cout_28_, cout_27_, cout_7__BAR, cout_6_, 
        cout_5_, cout_4_, cout_3_, cout_2_, cout_1_, cout_0_, cout_8__BAR, 
        cout_9__BAR, cout_10__BAR, cout_11__BAR, cout_12__BAR, cout_13__BAR, 
        cout_14__BAR, cout_15__BAR, cout_16__BAR, cout_17__BAR, cout_18__BAR, 
        cout_19__BAR, cout_20__BAR, cout_21__BAR, cout_22__BAR, cout_23__BAR, 
        cout_24__BAR, cout_25__BAR, cout_26__BAR, cout_29__BAR, cout_31__BAR, 
        cout_33__BAR, cout_35__BAR, cout_37__BAR, cout_39__BAR, cout_41__BAR, 
        cout_43__BAR, cout_45__BAR );
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  output cout_50_, cout_49_, cout_48_, cout_47_, cout_46_, cout_44_, cout_42_,
         cout_40_, cout_38_, cout_36_, cout_34_, cout_32_, cout_30_, cout_28_,
         cout_27_, cout_7__BAR, cout_6_, cout_5_, cout_4_, cout_3_, cout_2_,
         cout_1_, cout_0_, cout_8__BAR, cout_9__BAR, cout_10__BAR,
         cout_11__BAR, cout_12__BAR, cout_13__BAR, cout_14__BAR, cout_15__BAR,
         cout_16__BAR, cout_17__BAR, cout_18__BAR, cout_19__BAR, cout_20__BAR,
         cout_21__BAR, cout_22__BAR, cout_23__BAR, cout_24__BAR, cout_25__BAR,
         cout_26__BAR, cout_29__BAR, cout_31__BAR, cout_33__BAR, cout_35__BAR,
         cout_37__BAR, cout_39__BAR, cout_41__BAR, cout_43__BAR, cout_45__BAR;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11;

  NAND2X0 U1 ( .IN1(in2[8]), .IN2(in1[8]), .QN(cout_8__BAR) );
  NAND2X0 U2 ( .IN1(in2[9]), .IN2(in1[9]), .QN(cout_9__BAR) );
  NAND2X0 U3 ( .IN1(in2[10]), .IN2(in1[10]), .QN(cout_10__BAR) );
  NAND2X0 U4 ( .IN1(in2[11]), .IN2(in1[11]), .QN(cout_11__BAR) );
  NAND2X0 U5 ( .IN1(in2[12]), .IN2(in1[12]), .QN(cout_12__BAR) );
  NAND2X0 U6 ( .IN1(in2[13]), .IN2(in1[13]), .QN(cout_13__BAR) );
  NAND2X0 U7 ( .IN1(in2[14]), .IN2(in1[14]), .QN(cout_14__BAR) );
  NAND2X0 U8 ( .IN1(in2[15]), .IN2(in1[15]), .QN(cout_15__BAR) );
  NAND2X0 U9 ( .IN1(in2[16]), .IN2(in1[16]), .QN(cout_16__BAR) );
  NAND2X0 U10 ( .IN1(in2[17]), .IN2(in1[17]), .QN(cout_17__BAR) );
  NAND2X0 U11 ( .IN1(in2[18]), .IN2(in1[18]), .QN(cout_18__BAR) );
  NAND2X0 U12 ( .IN1(in2[19]), .IN2(in1[19]), .QN(cout_19__BAR) );
  NAND2X0 U13 ( .IN1(in2[20]), .IN2(in1[20]), .QN(cout_20__BAR) );
  NAND2X0 U14 ( .IN1(in2[21]), .IN2(in1[21]), .QN(cout_21__BAR) );
  NAND2X0 U15 ( .IN1(in2[22]), .IN2(in1[22]), .QN(cout_22__BAR) );
  NAND2X0 U16 ( .IN1(in2[23]), .IN2(in1[23]), .QN(cout_23__BAR) );
  NAND2X0 U17 ( .IN1(in2[24]), .IN2(in1[24]), .QN(cout_24__BAR) );
  NAND2X0 U18 ( .IN1(in2[25]), .IN2(in1[25]), .QN(cout_25__BAR) );
  NAND2X0 U19 ( .IN1(in2[26]), .IN2(in1[26]), .QN(cout_26__BAR) );
  NAND2X0 U20 ( .IN1(in2[29]), .IN2(in1[29]), .QN(cout_29__BAR) );
  NAND2X0 U21 ( .IN1(in2[31]), .IN2(in1[31]), .QN(cout_31__BAR) );
  NAND2X0 U22 ( .IN1(in2[33]), .IN2(in1[33]), .QN(cout_33__BAR) );
  NAND2X0 U23 ( .IN1(in2[35]), .IN2(in1[35]), .QN(cout_35__BAR) );
  NAND2X0 U24 ( .IN1(in2[37]), .IN2(in1[37]), .QN(cout_37__BAR) );
  NAND2X0 U25 ( .IN1(in2[39]), .IN2(in1[39]), .QN(cout_39__BAR) );
  NAND2X0 U26 ( .IN1(in2[41]), .IN2(in1[41]), .QN(cout_41__BAR) );
  NAND2X0 U27 ( .IN1(in2[43]), .IN2(in1[43]), .QN(cout_43__BAR) );
  NAND2X0 U28 ( .IN1(in2[45]), .IN2(in1[45]), .QN(cout_45__BAR) );
  NAND2X0 U29 ( .IN1(in2[7]), .IN2(in1[7]), .QN(cout_7__BAR) );
  NAND2X0 U30 ( .IN1(n1), .IN2(cout_27_), .QN(sumout[27]) );
  NAND2X0 U31 ( .IN1(in1[27]), .IN2(in2[27]), .QN(n1) );
  NAND2X0 U32 ( .IN1(n2), .IN2(cout_28_), .QN(sumout[28]) );
  NAND2X0 U33 ( .IN1(in1[28]), .IN2(in2[28]), .QN(n2) );
  NAND2X0 U34 ( .IN1(n3), .IN2(cout_30_), .QN(sumout[30]) );
  NAND2X0 U35 ( .IN1(in1[30]), .IN2(in2[30]), .QN(n3) );
  NAND2X0 U36 ( .IN1(n4), .IN2(cout_32_), .QN(sumout[32]) );
  NAND2X0 U37 ( .IN1(in1[32]), .IN2(in2[32]), .QN(n4) );
  NAND2X0 U38 ( .IN1(n5), .IN2(cout_34_), .QN(sumout[34]) );
  NAND2X0 U39 ( .IN1(in1[34]), .IN2(in2[34]), .QN(n5) );
  NAND2X0 U40 ( .IN1(n6), .IN2(cout_36_), .QN(sumout[36]) );
  NAND2X0 U41 ( .IN1(in1[36]), .IN2(in2[36]), .QN(n6) );
  NAND2X0 U42 ( .IN1(n7), .IN2(cout_38_), .QN(sumout[38]) );
  NAND2X0 U43 ( .IN1(in1[38]), .IN2(in2[38]), .QN(n7) );
  NAND2X0 U44 ( .IN1(n8), .IN2(cout_40_), .QN(sumout[40]) );
  NAND2X0 U45 ( .IN1(in1[40]), .IN2(in2[40]), .QN(n8) );
  NAND2X0 U46 ( .IN1(n9), .IN2(cout_42_), .QN(sumout[42]) );
  NAND2X0 U47 ( .IN1(in1[42]), .IN2(in2[42]), .QN(n9) );
  NAND2X0 U48 ( .IN1(n10), .IN2(cout_44_), .QN(sumout[44]) );
  NAND2X0 U49 ( .IN1(in1[44]), .IN2(in2[44]), .QN(n10) );
  NAND2X0 U50 ( .IN1(n11), .IN2(cout_46_), .QN(sumout[46]) );
  NAND2X0 U51 ( .IN1(in1[46]), .IN2(in2[46]), .QN(n11) );
  OR2X1 U52 ( .IN1(in2[27]), .IN2(in1[27]), .Q(cout_27_) );
  OR2X1 U53 ( .IN1(in2[28]), .IN2(in1[28]), .Q(cout_28_) );
  OR2X1 U54 ( .IN1(in2[30]), .IN2(in1[30]), .Q(cout_30_) );
  OR2X1 U55 ( .IN1(in2[32]), .IN2(in1[32]), .Q(cout_32_) );
  OR2X1 U56 ( .IN1(in2[34]), .IN2(in1[34]), .Q(cout_34_) );
  OR2X1 U57 ( .IN1(in2[36]), .IN2(in1[36]), .Q(cout_36_) );
  OR2X1 U58 ( .IN1(in2[38]), .IN2(in1[38]), .Q(cout_38_) );
  OR2X1 U59 ( .IN1(in2[40]), .IN2(in1[40]), .Q(cout_40_) );
  OR2X1 U60 ( .IN1(in2[42]), .IN2(in1[42]), .Q(cout_42_) );
  OR2X1 U61 ( .IN1(in2[44]), .IN2(in1[44]), .Q(cout_44_) );
  OR2X1 U62 ( .IN1(in2[46]), .IN2(in1[46]), .Q(cout_46_) );
  OA21X1 U63 ( .IN1(in2[8]), .IN2(in1[8]), .IN3(cout_8__BAR), .Q(sumout[8]) );
  OA21X1 U64 ( .IN1(in2[9]), .IN2(in1[9]), .IN3(cout_9__BAR), .Q(sumout[9]) );
  OA21X1 U65 ( .IN1(in2[10]), .IN2(in1[10]), .IN3(cout_10__BAR), .Q(sumout[10]) );
  OA21X1 U66 ( .IN1(in2[11]), .IN2(in1[11]), .IN3(cout_11__BAR), .Q(sumout[11]) );
  OA21X1 U67 ( .IN1(in2[12]), .IN2(in1[12]), .IN3(cout_12__BAR), .Q(sumout[12]) );
  OA21X1 U68 ( .IN1(in2[13]), .IN2(in1[13]), .IN3(cout_13__BAR), .Q(sumout[13]) );
  OA21X1 U69 ( .IN1(in2[14]), .IN2(in1[14]), .IN3(cout_14__BAR), .Q(sumout[14]) );
  OA21X1 U70 ( .IN1(in2[15]), .IN2(in1[15]), .IN3(cout_15__BAR), .Q(sumout[15]) );
  OA21X1 U71 ( .IN1(in2[16]), .IN2(in1[16]), .IN3(cout_16__BAR), .Q(sumout[16]) );
  OA21X1 U72 ( .IN1(in2[17]), .IN2(in1[17]), .IN3(cout_17__BAR), .Q(sumout[17]) );
  OA21X1 U73 ( .IN1(in2[18]), .IN2(in1[18]), .IN3(cout_18__BAR), .Q(sumout[18]) );
  OA21X1 U74 ( .IN1(in2[19]), .IN2(in1[19]), .IN3(cout_19__BAR), .Q(sumout[19]) );
  OA21X1 U75 ( .IN1(in2[20]), .IN2(in1[20]), .IN3(cout_20__BAR), .Q(sumout[20]) );
  OA21X1 U76 ( .IN1(in2[21]), .IN2(in1[21]), .IN3(cout_21__BAR), .Q(sumout[21]) );
  OA21X1 U77 ( .IN1(in2[22]), .IN2(in1[22]), .IN3(cout_22__BAR), .Q(sumout[22]) );
  OA21X1 U78 ( .IN1(in2[23]), .IN2(in1[23]), .IN3(cout_23__BAR), .Q(sumout[23]) );
  OA21X1 U79 ( .IN1(in2[24]), .IN2(in1[24]), .IN3(cout_24__BAR), .Q(sumout[24]) );
  OA21X1 U80 ( .IN1(in2[25]), .IN2(in1[25]), .IN3(cout_25__BAR), .Q(sumout[25]) );
  OA21X1 U81 ( .IN1(in2[26]), .IN2(in1[26]), .IN3(cout_26__BAR), .Q(sumout[26]) );
  OA21X1 U82 ( .IN1(in2[29]), .IN2(in1[29]), .IN3(cout_29__BAR), .Q(sumout[29]) );
  OA21X1 U83 ( .IN1(in2[31]), .IN2(in1[31]), .IN3(cout_31__BAR), .Q(sumout[31]) );
  OA21X1 U84 ( .IN1(in2[33]), .IN2(in1[33]), .IN3(cout_33__BAR), .Q(sumout[33]) );
  OA21X1 U85 ( .IN1(in2[35]), .IN2(in1[35]), .IN3(cout_35__BAR), .Q(sumout[35]) );
  OA21X1 U86 ( .IN1(in2[37]), .IN2(in1[37]), .IN3(cout_37__BAR), .Q(sumout[37]) );
  OA21X1 U87 ( .IN1(in2[39]), .IN2(in1[39]), .IN3(cout_39__BAR), .Q(sumout[39]) );
  OA21X1 U88 ( .IN1(in2[41]), .IN2(in1[41]), .IN3(cout_41__BAR), .Q(sumout[41]) );
  OA21X1 U89 ( .IN1(in2[43]), .IN2(in1[43]), .IN3(cout_43__BAR), .Q(sumout[43]) );
  OA21X1 U90 ( .IN1(in2[45]), .IN2(in1[45]), .IN3(cout_45__BAR), .Q(sumout[45]) );
  XOR2X1 U91 ( .IN1(in1[47]), .IN2(in2[47]), .Q(sumout[47]) );
endmodule


module csa51squ_38 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;


  AO222X1 U1 ( .IN1(in2[6]), .IN2(in3[6]), .IN3(in2[6]), .IN4(in1[6]), .IN5(
        in3[6]), .IN6(in1[6]), .Q(cout[6]) );
  FADDX1 U2 ( .A(in1[10]), .B(in2[10]), .CI(in3[10]), .CO(cout[10]), .S(
        sumout[10]) );
  FADDX1 U3 ( .A(in1[11]), .B(in2[11]), .CI(in3[11]), .CO(cout[11]), .S(
        sumout[11]) );
  FADDX1 U4 ( .A(in1[12]), .B(in2[12]), .CI(in3[12]), .CO(cout[12]), .S(
        sumout[12]) );
  FADDX1 U5 ( .A(in1[13]), .B(in2[13]), .CI(in3[13]), .CO(cout[13]), .S(
        sumout[13]) );
  FADDX1 U6 ( .A(in1[14]), .B(in2[14]), .CI(in3[14]), .CO(cout[14]), .S(
        sumout[14]) );
  FADDX1 U7 ( .A(in1[15]), .B(in2[15]), .CI(in3[15]), .CO(cout[15]), .S(
        sumout[15]) );
  FADDX1 U8 ( .A(in1[16]), .B(in2[16]), .CI(in3[16]), .CO(cout[16]), .S(
        sumout[16]) );
  FADDX1 U9 ( .A(in1[17]), .B(in2[17]), .CI(in3[17]), .CO(cout[17]), .S(
        sumout[17]) );
  FADDX1 U10 ( .A(in1[18]), .B(in2[18]), .CI(in3[18]), .CO(cout[18]), .S(
        sumout[18]) );
  FADDX1 U11 ( .A(in1[19]), .B(in2[19]), .CI(in3[19]), .CO(cout[19]), .S(
        sumout[19]) );
  FADDX1 U12 ( .A(in1[20]), .B(in2[20]), .CI(in3[20]), .CO(cout[20]), .S(
        sumout[20]) );
  FADDX1 U13 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U14 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U15 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U16 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U17 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U18 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U19 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U20 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U21 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U22 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U23 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U24 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
  FADDX1 U25 ( .A(in1[33]), .B(in2[33]), .CI(in3[33]), .CO(cout[33]), .S(
        sumout[33]) );
  FADDX1 U26 ( .A(in1[34]), .B(in2[34]), .CI(in3[34]), .CO(cout[34]), .S(
        sumout[34]) );
  FADDX1 U27 ( .A(in1[35]), .B(in2[35]), .CI(in3[35]), .CO(cout[35]), .S(
        sumout[35]) );
  FADDX1 U28 ( .A(in1[36]), .B(in2[36]), .CI(in3[36]), .CO(cout[36]), .S(
        sumout[36]) );
  FADDX1 U29 ( .A(in1[37]), .B(in2[37]), .CI(in3[37]), .CO(cout[37]), .S(
        sumout[37]) );
  FADDX1 U30 ( .A(in1[38]), .B(in2[38]), .CI(in3[38]), .CO(cout[38]), .S(
        sumout[38]) );
  FADDX1 U31 ( .A(in1[39]), .B(in2[39]), .CI(in3[39]), .CO(cout[39]), .S(
        sumout[39]) );
  FADDX1 U32 ( .A(in1[40]), .B(in2[40]), .CI(in3[40]), .CO(cout[40]), .S(
        sumout[40]) );
  FADDX1 U33 ( .A(in1[41]), .B(in2[41]), .CI(in3[41]), .CO(cout[41]), .S(
        sumout[41]) );
  FADDX1 U34 ( .A(in1[42]), .B(in2[42]), .CI(in3[42]), .CO(cout[42]), .S(
        sumout[42]) );
  FADDX1 U35 ( .A(in1[43]), .B(in2[43]), .CI(in3[43]), .CO(cout[43]), .S(
        sumout[43]) );
  FADDX1 U36 ( .A(in1[44]), .B(in2[44]), .CI(in3[44]), .CO(cout[44]), .S(
        sumout[44]) );
  FADDX1 U37 ( .A(in1[45]), .B(in2[45]), .CI(in3[45]), .CO(cout[45]), .S(
        sumout[45]) );
  FADDX1 U38 ( .A(in1[46]), .B(in2[46]), .CI(in3[46]), .CO(cout[46]), .S(
        sumout[46]) );
  XOR3X1 U39 ( .IN1(in2[47]), .IN2(in3[47]), .IN3(in1[47]), .Q(sumout[47]) );
  FADDX1 U40 ( .A(in1[7]), .B(in2[7]), .CI(in3[7]), .CO(cout[7]), .S(sumout[7]) );
  FADDX1 U41 ( .A(in1[8]), .B(in2[8]), .CI(in3[8]), .CO(cout[8]), .S(sumout[8]) );
  FADDX1 U42 ( .A(in1[9]), .B(in2[9]), .CI(in3[9]), .CO(cout[9]), .S(sumout[9]) );
endmodule


module csa51squ_39 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14;

  AND2X1 U1 ( .IN1(in2[7]), .IN2(in1[7]), .Q(cout[7]) );
  NOR2X0 U2 ( .IN1(in2[7]), .IN2(in1[7]), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(cout[7]), .QN(sumout[7]) );
  AND2X1 U4 ( .IN1(in2[8]), .IN2(in1[8]), .Q(cout[8]) );
  NOR2X0 U5 ( .IN1(in2[8]), .IN2(in1[8]), .QN(n2) );
  NOR2X0 U6 ( .IN1(n2), .IN2(cout[8]), .QN(sumout[8]) );
  AND2X1 U7 ( .IN1(in2[9]), .IN2(in1[9]), .Q(cout[9]) );
  NOR2X0 U8 ( .IN1(in2[9]), .IN2(in1[9]), .QN(n3) );
  NOR2X0 U9 ( .IN1(n3), .IN2(cout[9]), .QN(sumout[9]) );
  AND2X1 U10 ( .IN1(in2[10]), .IN2(in1[10]), .Q(cout[10]) );
  NOR2X0 U11 ( .IN1(in2[10]), .IN2(in1[10]), .QN(n4) );
  NOR2X0 U12 ( .IN1(n4), .IN2(cout[10]), .QN(sumout[10]) );
  AND2X1 U13 ( .IN1(in2[11]), .IN2(in1[11]), .Q(cout[11]) );
  NOR2X0 U14 ( .IN1(in2[11]), .IN2(in1[11]), .QN(n5) );
  NOR2X0 U15 ( .IN1(n5), .IN2(cout[11]), .QN(sumout[11]) );
  AND2X1 U16 ( .IN1(in2[12]), .IN2(in1[12]), .Q(cout[12]) );
  NOR2X0 U17 ( .IN1(in2[12]), .IN2(in1[12]), .QN(n6) );
  NOR2X0 U18 ( .IN1(n6), .IN2(cout[12]), .QN(sumout[12]) );
  AND2X1 U19 ( .IN1(in3[40]), .IN2(in2[40]), .Q(cout[40]) );
  NOR2X0 U20 ( .IN1(in3[40]), .IN2(in2[40]), .QN(n7) );
  NOR2X0 U21 ( .IN1(n7), .IN2(cout[40]), .QN(sumout[40]) );
  AND2X1 U22 ( .IN1(in3[41]), .IN2(in2[41]), .Q(cout[41]) );
  NOR2X0 U23 ( .IN1(in3[41]), .IN2(in2[41]), .QN(n8) );
  NOR2X0 U24 ( .IN1(n8), .IN2(cout[41]), .QN(sumout[41]) );
  AND2X1 U25 ( .IN1(in3[42]), .IN2(in2[42]), .Q(cout[42]) );
  NOR2X0 U26 ( .IN1(in3[42]), .IN2(in2[42]), .QN(n9) );
  NOR2X0 U27 ( .IN1(n9), .IN2(cout[42]), .QN(sumout[42]) );
  AND2X1 U28 ( .IN1(in3[43]), .IN2(in2[43]), .Q(cout[43]) );
  NOR2X0 U29 ( .IN1(in3[43]), .IN2(in2[43]), .QN(n10) );
  NOR2X0 U30 ( .IN1(n10), .IN2(cout[43]), .QN(sumout[43]) );
  AND2X1 U31 ( .IN1(in3[44]), .IN2(in2[44]), .Q(cout[44]) );
  NOR2X0 U32 ( .IN1(in3[44]), .IN2(in2[44]), .QN(n11) );
  NOR2X0 U33 ( .IN1(n11), .IN2(cout[44]), .QN(sumout[44]) );
  AND2X1 U34 ( .IN1(in3[45]), .IN2(in2[45]), .Q(cout[45]) );
  NOR2X0 U35 ( .IN1(in3[45]), .IN2(in2[45]), .QN(n12) );
  NOR2X0 U36 ( .IN1(n12), .IN2(cout[45]), .QN(sumout[45]) );
  AND2X1 U37 ( .IN1(in3[46]), .IN2(in2[46]), .Q(cout[46]) );
  NOR2X0 U38 ( .IN1(in3[46]), .IN2(in2[46]), .QN(n13) );
  NOR2X0 U39 ( .IN1(n13), .IN2(cout[46]), .QN(sumout[46]) );
  INVX0 U40 ( .INP(in3[47]), .ZN(sumout[47]) );
  AND2X1 U41 ( .IN1(in2[5]), .IN2(in1[5]), .Q(cout[5]) );
  AND2X1 U42 ( .IN1(in2[6]), .IN2(in1[6]), .Q(cout[6]) );
  NOR2X0 U43 ( .IN1(in2[6]), .IN2(in1[6]), .QN(n14) );
  NOR2X0 U44 ( .IN1(n14), .IN2(cout[6]), .QN(sumout[6]) );
  FADDX1 U45 ( .A(in1[13]), .B(in2[13]), .CI(in3[13]), .CO(cout[13]), .S(
        sumout[13]) );
  FADDX1 U46 ( .A(in1[14]), .B(in2[14]), .CI(in3[14]), .CO(cout[14]), .S(
        sumout[14]) );
  FADDX1 U47 ( .A(in1[15]), .B(in2[15]), .CI(in3[15]), .CO(cout[15]), .S(
        sumout[15]) );
  FADDX1 U48 ( .A(in1[16]), .B(in2[16]), .CI(in3[16]), .CO(cout[16]), .S(
        sumout[16]) );
  FADDX1 U49 ( .A(in1[17]), .B(in2[17]), .CI(in3[17]), .CO(cout[17]), .S(
        sumout[17]) );
  FADDX1 U50 ( .A(in1[18]), .B(in2[18]), .CI(in3[18]), .CO(cout[18]), .S(
        sumout[18]) );
  FADDX1 U51 ( .A(in1[19]), .B(in2[19]), .CI(in3[19]), .CO(cout[19]), .S(
        sumout[19]) );
  FADDX1 U52 ( .A(in1[20]), .B(in2[20]), .CI(in3[20]), .CO(cout[20]), .S(
        sumout[20]) );
  FADDX1 U53 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U54 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U55 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U56 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U57 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U58 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U59 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U60 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U61 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U62 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U63 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U64 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
  FADDX1 U65 ( .A(in1[33]), .B(in2[33]), .CI(in3[33]), .CO(cout[33]), .S(
        sumout[33]) );
  FADDX1 U66 ( .A(in1[34]), .B(in2[34]), .CI(in3[34]), .CO(cout[34]), .S(
        sumout[34]) );
  FADDX1 U67 ( .A(in1[35]), .B(in2[35]), .CI(in3[35]), .CO(cout[35]), .S(
        sumout[35]) );
  FADDX1 U68 ( .A(in1[36]), .B(in2[36]), .CI(in3[36]), .CO(cout[36]), .S(
        sumout[36]) );
  FADDX1 U69 ( .A(in1[37]), .B(in2[37]), .CI(in3[37]), .CO(cout[37]), .S(
        sumout[37]) );
  FADDX1 U70 ( .A(in1[38]), .B(in2[38]), .CI(in3[38]), .CO(cout[38]), .S(
        sumout[38]) );
  FADDX1 U71 ( .A(in1[39]), .B(in2[39]), .CI(in3[39]), .CO(cout[39]), .S(
        sumout[39]) );
endmodule


module csa51squ_40 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17;

  NBUFFX2 U1 ( .INP(in1[6]), .Z(sumout[6]) );
  NBUFFX2 U2 ( .INP(in1[7]), .Z(sumout[7]) );
  NBUFFX2 U3 ( .INP(in1[8]), .Z(sumout[8]) );
  NBUFFX2 U4 ( .INP(in1[9]), .Z(sumout[9]) );
  NBUFFX2 U5 ( .INP(in1[10]), .Z(sumout[10]) );
  NBUFFX2 U6 ( .INP(in1[11]), .Z(sumout[11]) );
  AND2X1 U7 ( .IN1(in3[13]), .IN2(in1[13]), .Q(cout[13]) );
  NOR2X0 U8 ( .IN1(in3[13]), .IN2(in1[13]), .QN(n7) );
  NOR2X0 U9 ( .IN1(n7), .IN2(cout[13]), .QN(sumout[13]) );
  AND2X1 U10 ( .IN1(in3[15]), .IN2(in1[15]), .Q(cout[15]) );
  NOR2X0 U11 ( .IN1(in3[15]), .IN2(in1[15]), .QN(n8) );
  NOR2X0 U12 ( .IN1(n8), .IN2(cout[15]), .QN(sumout[15]) );
  AND2X1 U13 ( .IN1(in3[17]), .IN2(in1[17]), .Q(cout[17]) );
  NOR2X0 U14 ( .IN1(in3[17]), .IN2(in1[17]), .QN(n9) );
  NOR2X0 U15 ( .IN1(n9), .IN2(cout[17]), .QN(sumout[17]) );
  AND2X1 U16 ( .IN1(in3[43]), .IN2(in2[43]), .Q(cout[43]) );
  NOR2X0 U17 ( .IN1(in3[43]), .IN2(in2[43]), .QN(n10) );
  NOR2X0 U18 ( .IN1(n10), .IN2(cout[43]), .QN(sumout[43]) );
  AND2X1 U19 ( .IN1(in3[44]), .IN2(in2[44]), .Q(cout[44]) );
  NOR2X0 U20 ( .IN1(in3[44]), .IN2(in2[44]), .QN(n11) );
  NOR2X0 U21 ( .IN1(n11), .IN2(cout[44]), .QN(sumout[44]) );
  AND2X1 U22 ( .IN1(in3[45]), .IN2(in2[45]), .Q(cout[45]) );
  NOR2X0 U23 ( .IN1(in3[45]), .IN2(in2[45]), .QN(n12) );
  NOR2X0 U24 ( .IN1(n12), .IN2(cout[45]), .QN(sumout[45]) );
  AND2X1 U25 ( .IN1(in3[46]), .IN2(in2[46]), .Q(cout[46]) );
  NOR2X0 U26 ( .IN1(in3[46]), .IN2(in2[46]), .QN(n13) );
  NOR2X0 U27 ( .IN1(n13), .IN2(cout[46]), .QN(sumout[46]) );
  XOR2X1 U28 ( .IN1(in3[47]), .IN2(in2[47]), .Q(sumout[47]) );
  AND2X1 U29 ( .IN1(in3[12]), .IN2(in1[12]), .Q(cout[12]) );
  NOR2X0 U30 ( .IN1(in3[12]), .IN2(in1[12]), .QN(n14) );
  NOR2X0 U31 ( .IN1(n14), .IN2(cout[12]), .QN(sumout[12]) );
  AND2X1 U32 ( .IN1(in3[14]), .IN2(in1[14]), .Q(cout[14]) );
  NOR2X0 U33 ( .IN1(in3[14]), .IN2(in1[14]), .QN(n15) );
  NOR2X0 U34 ( .IN1(n15), .IN2(cout[14]), .QN(sumout[14]) );
  AND2X1 U35 ( .IN1(in3[16]), .IN2(in1[16]), .Q(cout[16]) );
  NOR2X0 U36 ( .IN1(in3[16]), .IN2(in1[16]), .QN(n16) );
  NOR2X0 U37 ( .IN1(n16), .IN2(cout[16]), .QN(sumout[16]) );
  AND2X1 U38 ( .IN1(in3[18]), .IN2(in1[18]), .Q(cout[18]) );
  NOR2X0 U39 ( .IN1(in3[18]), .IN2(in1[18]), .QN(n17) );
  NOR2X0 U40 ( .IN1(n17), .IN2(cout[18]), .QN(sumout[18]) );
  FADDX1 U41 ( .A(in1[19]), .B(in2[19]), .CI(in3[19]), .CO(cout[19]), .S(
        sumout[19]) );
  FADDX1 U42 ( .A(in1[20]), .B(in2[20]), .CI(in3[20]), .CO(cout[20]), .S(
        sumout[20]) );
  FADDX1 U43 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U44 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U45 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U46 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U47 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U48 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U49 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U50 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U51 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U52 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U53 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U54 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
  FADDX1 U55 ( .A(in1[33]), .B(in2[33]), .CI(in3[33]), .CO(cout[33]), .S(
        sumout[33]) );
  FADDX1 U56 ( .A(in1[34]), .B(in2[34]), .CI(in3[34]), .CO(cout[34]), .S(
        sumout[34]) );
  FADDX1 U57 ( .A(in1[35]), .B(in2[35]), .CI(in3[35]), .CO(cout[35]), .S(
        sumout[35]) );
  FADDX1 U58 ( .A(in1[36]), .B(in2[36]), .CI(in3[36]), .CO(cout[36]), .S(
        sumout[36]) );
  FADDX1 U59 ( .A(in1[37]), .B(in2[37]), .CI(in3[37]), .CO(cout[37]), .S(
        sumout[37]) );
  FADDX1 U60 ( .A(in1[38]), .B(in2[38]), .CI(in3[38]), .CO(cout[38]), .S(
        sumout[38]) );
  FADDX1 U61 ( .A(in1[39]), .B(in2[39]), .CI(in3[39]), .CO(cout[39]), .S(
        sumout[39]) );
  FADDX1 U62 ( .A(in1[40]), .B(in2[40]), .CI(in3[40]), .CO(cout[40]), .S(
        sumout[40]) );
  FADDX1 U63 ( .A(in1[41]), .B(in2[41]), .CI(in3[41]), .CO(cout[41]), .S(
        sumout[41]) );
  FADDX1 U64 ( .A(in1[42]), .B(in2[42]), .CI(in3[42]), .CO(cout[42]), .S(
        sumout[42]) );
endmodule


module csa51squ_41 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19;

  NBUFFX2 U1 ( .INP(in2[46]), .Z(sumout[46]) );
  NBUFFX2 U2 ( .INP(in2[45]), .Z(sumout[45]) );
  NBUFFX2 U3 ( .INP(in2[44]), .Z(sumout[44]) );
  NBUFFX2 U4 ( .INP(in2[43]), .Z(sumout[43]) );
  NBUFFX2 U5 ( .INP(in2[42]), .Z(sumout[42]) );
  NBUFFX2 U6 ( .INP(in2[41]), .Z(sumout[41]) );
  NBUFFX2 U7 ( .INP(in2[40]), .Z(sumout[40]) );
  NBUFFX2 U8 ( .INP(in2[39]), .Z(sumout[39]) );
  AND2X1 U9 ( .IN1(in2[7]), .IN2(in1[7]), .Q(cout[7]) );
  NOR2X0 U10 ( .IN1(in2[7]), .IN2(in1[7]), .QN(n9) );
  NOR2X0 U11 ( .IN1(n9), .IN2(cout[7]), .QN(sumout[7]) );
  AND2X1 U12 ( .IN1(in2[8]), .IN2(in1[8]), .Q(cout[8]) );
  NOR2X0 U13 ( .IN1(in2[8]), .IN2(in1[8]), .QN(n10) );
  NOR2X0 U14 ( .IN1(n10), .IN2(cout[8]), .QN(sumout[8]) );
  AND2X1 U15 ( .IN1(in2[9]), .IN2(in1[9]), .Q(cout[9]) );
  NOR2X0 U16 ( .IN1(in2[9]), .IN2(in1[9]), .QN(n11) );
  NOR2X0 U17 ( .IN1(n11), .IN2(cout[9]), .QN(sumout[9]) );
  AND2X1 U18 ( .IN1(in3[33]), .IN2(in2[33]), .Q(cout[33]) );
  NOR2X0 U19 ( .IN1(in3[33]), .IN2(in2[33]), .QN(n12) );
  NOR2X0 U20 ( .IN1(n12), .IN2(cout[33]), .QN(sumout[33]) );
  AND2X1 U21 ( .IN1(in3[34]), .IN2(in2[34]), .Q(cout[34]) );
  NOR2X0 U22 ( .IN1(in3[34]), .IN2(in2[34]), .QN(n13) );
  NOR2X0 U23 ( .IN1(n13), .IN2(cout[34]), .QN(sumout[34]) );
  AND2X1 U24 ( .IN1(in3[35]), .IN2(in2[35]), .Q(cout[35]) );
  NOR2X0 U25 ( .IN1(in3[35]), .IN2(in2[35]), .QN(n14) );
  NOR2X0 U26 ( .IN1(n14), .IN2(cout[35]), .QN(sumout[35]) );
  AND2X1 U27 ( .IN1(in3[36]), .IN2(in2[36]), .Q(cout[36]) );
  NOR2X0 U28 ( .IN1(in3[36]), .IN2(in2[36]), .QN(n15) );
  NOR2X0 U29 ( .IN1(n15), .IN2(cout[36]), .QN(sumout[36]) );
  AND2X1 U30 ( .IN1(in3[37]), .IN2(in2[37]), .Q(cout[37]) );
  NOR2X0 U31 ( .IN1(in3[37]), .IN2(in2[37]), .QN(n16) );
  NOR2X0 U32 ( .IN1(n16), .IN2(cout[37]), .QN(sumout[37]) );
  AND2X1 U33 ( .IN1(in3[38]), .IN2(in2[38]), .Q(cout[38]) );
  NOR2X0 U34 ( .IN1(in3[38]), .IN2(in2[38]), .QN(n17) );
  NOR2X0 U35 ( .IN1(n17), .IN2(cout[38]), .QN(sumout[38]) );
  AND2X1 U36 ( .IN1(in2[4]), .IN2(in1[4]), .Q(cout[4]) );
  AND2X1 U37 ( .IN1(in2[5]), .IN2(in1[5]), .Q(cout[5]) );
  NOR2X0 U38 ( .IN1(in2[5]), .IN2(in1[5]), .QN(n18) );
  NOR2X0 U39 ( .IN1(n18), .IN2(cout[5]), .QN(sumout[5]) );
  AND2X1 U40 ( .IN1(in2[6]), .IN2(in1[6]), .Q(cout[6]) );
  NOR2X0 U41 ( .IN1(in2[6]), .IN2(in1[6]), .QN(n19) );
  NOR2X0 U42 ( .IN1(n19), .IN2(cout[6]), .QN(sumout[6]) );
  FADDX1 U43 ( .A(in1[10]), .B(in2[10]), .CI(in3[10]), .CO(cout[10]), .S(
        sumout[10]) );
  FADDX1 U44 ( .A(in1[11]), .B(in2[11]), .CI(in3[11]), .CO(cout[11]), .S(
        sumout[11]) );
  FADDX1 U45 ( .A(in1[12]), .B(in2[12]), .CI(in3[12]), .CO(cout[12]), .S(
        sumout[12]) );
  FADDX1 U46 ( .A(in1[13]), .B(in2[13]), .CI(in3[13]), .CO(cout[13]), .S(
        sumout[13]) );
  FADDX1 U47 ( .A(in1[14]), .B(in2[14]), .CI(in3[14]), .CO(cout[14]), .S(
        sumout[14]) );
  FADDX1 U48 ( .A(in1[15]), .B(in2[15]), .CI(in3[15]), .CO(cout[15]), .S(
        sumout[15]) );
  FADDX1 U49 ( .A(in1[16]), .B(in2[16]), .CI(in3[16]), .CO(cout[16]), .S(
        sumout[16]) );
  FADDX1 U50 ( .A(in1[17]), .B(in2[17]), .CI(in3[17]), .CO(cout[17]), .S(
        sumout[17]) );
  FADDX1 U51 ( .A(in1[18]), .B(in2[18]), .CI(in3[18]), .CO(cout[18]), .S(
        sumout[18]) );
  FADDX1 U52 ( .A(in1[19]), .B(in2[19]), .CI(in3[19]), .CO(cout[19]), .S(
        sumout[19]) );
  FADDX1 U53 ( .A(in1[20]), .B(in2[20]), .CI(in3[20]), .CO(cout[20]), .S(
        sumout[20]) );
  FADDX1 U54 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U55 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U56 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U57 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U58 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U59 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U60 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U61 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U62 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U63 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U64 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U65 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
endmodule


module csa51squ_42 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n7, n8, n9, n10, n11, n12, n13;

  NBUFFX2 U1 ( .INP(in1[12]), .Z(sumout[12]) );
  NBUFFX2 U2 ( .INP(in1[13]), .Z(sumout[13]) );
  NBUFFX2 U3 ( .INP(in1[14]), .Z(sumout[14]) );
  NBUFFX2 U4 ( .INP(in1[15]), .Z(sumout[15]) );
  NBUFFX2 U5 ( .INP(in1[16]), .Z(sumout[16]) );
  NBUFFX2 U6 ( .INP(in1[17]), .Z(sumout[17]) );
  AND2X1 U7 ( .IN1(in3[19]), .IN2(in1[19]), .Q(cout[19]) );
  NOR2X0 U8 ( .IN1(in3[19]), .IN2(in1[19]), .QN(n7) );
  NOR2X0 U9 ( .IN1(n7), .IN2(cout[19]), .QN(sumout[19]) );
  AND2X1 U10 ( .IN1(in3[44]), .IN2(in2[44]), .Q(cout[44]) );
  NOR2X0 U11 ( .IN1(in3[44]), .IN2(in2[44]), .QN(n8) );
  NOR2X0 U12 ( .IN1(n8), .IN2(cout[44]), .QN(sumout[44]) );
  AND2X1 U13 ( .IN1(in3[45]), .IN2(in2[45]), .Q(cout[45]) );
  NOR2X0 U14 ( .IN1(in3[45]), .IN2(in2[45]), .QN(n9) );
  NOR2X0 U15 ( .IN1(n9), .IN2(cout[45]), .QN(sumout[45]) );
  AND2X1 U16 ( .IN1(in3[46]), .IN2(in2[46]), .Q(cout[46]) );
  NOR2X0 U17 ( .IN1(in3[46]), .IN2(in2[46]), .QN(n10) );
  NOR2X0 U18 ( .IN1(n10), .IN2(cout[46]), .QN(sumout[46]) );
  XOR2X1 U19 ( .IN1(in3[47]), .IN2(in2[47]), .Q(sumout[47]) );
  AND2X1 U20 ( .IN1(in3[18]), .IN2(in1[18]), .Q(cout[18]) );
  NOR2X0 U21 ( .IN1(in3[18]), .IN2(in1[18]), .QN(n11) );
  NOR2X0 U22 ( .IN1(n11), .IN2(cout[18]), .QN(sumout[18]) );
  AND2X1 U23 ( .IN1(in3[20]), .IN2(in1[20]), .Q(cout[20]) );
  NOR2X0 U24 ( .IN1(in3[20]), .IN2(in1[20]), .QN(n12) );
  NOR2X0 U25 ( .IN1(n12), .IN2(cout[20]), .QN(sumout[20]) );
  INVX0 U26 ( .INP(in1[42]), .ZN(n13) );
  FADDX1 U27 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U28 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U29 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U30 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U31 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U32 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U33 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U34 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U35 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U36 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U37 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U38 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
  FADDX1 U39 ( .A(in1[33]), .B(in2[33]), .CI(in3[33]), .CO(cout[33]), .S(
        sumout[33]) );
  FADDX1 U40 ( .A(in1[34]), .B(in2[34]), .CI(in3[34]), .CO(cout[34]), .S(
        sumout[34]) );
  FADDX1 U41 ( .A(in1[35]), .B(in2[35]), .CI(in3[35]), .CO(cout[35]), .S(
        sumout[35]) );
  FADDX1 U42 ( .A(in1[36]), .B(in2[36]), .CI(in3[36]), .CO(cout[36]), .S(
        sumout[36]) );
  FADDX1 U43 ( .A(in1[37]), .B(in2[37]), .CI(in3[37]), .CO(cout[37]), .S(
        sumout[37]) );
  FADDX1 U44 ( .A(in1[38]), .B(in2[38]), .CI(in3[38]), .CO(cout[38]), .S(
        sumout[38]) );
  FADDX1 U45 ( .A(in1[39]), .B(in2[39]), .CI(in3[39]), .CO(cout[39]), .S(
        sumout[39]) );
  FADDX1 U46 ( .A(in1[40]), .B(in2[40]), .CI(in3[40]), .CO(cout[40]), .S(
        sumout[40]) );
  FADDX1 U47 ( .A(in1[41]), .B(in2[41]), .CI(in3[41]), .CO(cout[41]), .S(
        sumout[41]) );
  FADDX1 U48 ( .A(in1[42]), .B(in2[42]), .CI(in3[42]), .CO(cout[42]), .S(
        sumout[42]) );
  FADDX1 U49 ( .A(in2[43]), .B(in3[43]), .CI(n13), .CO(cout[43]), .S(
        sumout[43]) );
endmodule


module csa51squ_43 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n9, n10, n11, n12, n13, n14, n15;

  NBUFFX2 U1 ( .INP(in2[6]), .Z(sumout[6]) );
  NBUFFX2 U2 ( .INP(in2[7]), .Z(sumout[7]) );
  NBUFFX2 U3 ( .INP(in2[8]), .Z(sumout[8]) );
  NBUFFX2 U4 ( .INP(in3[42]), .Z(sumout[42]) );
  NBUFFX2 U5 ( .INP(in3[41]), .Z(sumout[41]) );
  NBUFFX2 U6 ( .INP(in3[39]), .Z(sumout[39]) );
  NBUFFX2 U7 ( .INP(in3[38]), .Z(sumout[38]) );
  NBUFFX2 U8 ( .INP(in3[40]), .Z(sumout[40]) );
  AND2X1 U9 ( .IN1(in2[13]), .IN2(in1[13]), .Q(cout[13]) );
  NOR2X0 U10 ( .IN1(in2[13]), .IN2(in1[13]), .QN(n9) );
  NOR2X0 U11 ( .IN1(n9), .IN2(cout[13]), .QN(sumout[13]) );
  AND2X1 U12 ( .IN1(in2[37]), .IN2(in3[37]), .Q(cout[37]) );
  INVX0 U13 ( .INP(in2[37]), .ZN(n15) );
  MUX21X1 U14 ( .IN1(in2[37]), .IN2(n15), .S(in3[37]), .Q(sumout[37]) );
  AND2X1 U15 ( .IN1(in2[9]), .IN2(in1[9]), .Q(cout[9]) );
  NOR2X0 U16 ( .IN1(in2[9]), .IN2(in1[9]), .QN(n10) );
  NOR2X0 U17 ( .IN1(n10), .IN2(cout[9]), .QN(sumout[9]) );
  AND2X1 U18 ( .IN1(in2[10]), .IN2(in1[10]), .Q(cout[10]) );
  NOR2X0 U19 ( .IN1(in2[10]), .IN2(in1[10]), .QN(n11) );
  NOR2X0 U20 ( .IN1(n11), .IN2(cout[10]), .QN(sumout[10]) );
  AND2X1 U21 ( .IN1(in2[11]), .IN2(in1[11]), .Q(cout[11]) );
  NOR2X0 U22 ( .IN1(in2[11]), .IN2(in1[11]), .QN(n12) );
  NOR2X0 U23 ( .IN1(n12), .IN2(cout[11]), .QN(sumout[11]) );
  AND2X1 U24 ( .IN1(in2[12]), .IN2(in1[12]), .Q(cout[12]) );
  NOR2X0 U25 ( .IN1(in2[12]), .IN2(in1[12]), .QN(n13) );
  NOR2X0 U26 ( .IN1(n13), .IN2(cout[12]), .QN(sumout[12]) );
  AND2X1 U27 ( .IN1(in2[14]), .IN2(in1[14]), .Q(cout[14]) );
  NOR2X0 U28 ( .IN1(in2[14]), .IN2(in1[14]), .QN(n14) );
  NOR2X0 U29 ( .IN1(n14), .IN2(cout[14]), .QN(sumout[14]) );
  FADDX1 U30 ( .A(in1[15]), .B(in2[15]), .CI(in3[15]), .CO(cout[15]), .S(
        sumout[15]) );
  FADDX1 U31 ( .A(in1[16]), .B(in2[16]), .CI(in3[16]), .CO(cout[16]), .S(
        sumout[16]) );
  FADDX1 U32 ( .A(in1[17]), .B(in2[17]), .CI(in3[17]), .CO(cout[17]), .S(
        sumout[17]) );
  FADDX1 U33 ( .A(in1[18]), .B(in2[18]), .CI(in3[18]), .CO(cout[18]), .S(
        sumout[18]) );
  FADDX1 U34 ( .A(in1[19]), .B(in2[19]), .CI(in3[19]), .CO(cout[19]), .S(
        sumout[19]) );
  FADDX1 U35 ( .A(in1[20]), .B(in2[20]), .CI(in3[20]), .CO(cout[20]), .S(
        sumout[20]) );
  FADDX1 U36 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U37 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U38 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U39 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U40 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U41 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U42 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U43 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U44 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U45 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U46 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U47 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
  FADDX1 U48 ( .A(in1[33]), .B(in2[33]), .CI(in3[33]), .CO(cout[33]), .S(
        sumout[33]) );
  FADDX1 U49 ( .A(in1[34]), .B(in2[34]), .CI(in3[34]), .CO(cout[34]), .S(
        sumout[34]) );
  FADDX1 U50 ( .A(in1[35]), .B(in2[35]), .CI(in3[35]), .CO(cout[35]), .S(
        sumout[35]) );
  FADDX1 U51 ( .A(in1[36]), .B(in3[36]), .CI(n15), .CO(cout[36]), .S(
        sumout[36]) );
endmodule


module csa51squ_44 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36;

  NBUFFX2 U1 ( .INP(in3[46]), .Z(sumout[46]) );
  NBUFFX2 U2 ( .INP(in3[45]), .Z(sumout[45]) );
  NBUFFX2 U3 ( .INP(in3[44]), .Z(sumout[44]) );
  NBUFFX2 U4 ( .INP(in3[43]), .Z(sumout[43]) );
  NBUFFX2 U5 ( .INP(in3[42]), .Z(sumout[42]) );
  NBUFFX2 U6 ( .INP(in3[33]), .Z(sumout[33]) );
  NBUFFX2 U7 ( .INP(in3[32]), .Z(sumout[32]) );
  NBUFFX2 U8 ( .INP(in3[37]), .Z(sumout[37]) );
  NBUFFX2 U9 ( .INP(in3[36]), .Z(sumout[36]) );
  NBUFFX2 U10 ( .INP(in3[35]), .Z(sumout[35]) );
  NBUFFX2 U11 ( .INP(in3[34]), .Z(sumout[34]) );
  NBUFFX2 U12 ( .INP(in3[41]), .Z(sumout[41]) );
  NBUFFX2 U13 ( .INP(in3[40]), .Z(sumout[40]) );
  NBUFFX2 U14 ( .INP(in3[39]), .Z(sumout[39]) );
  NBUFFX2 U15 ( .INP(in3[38]), .Z(sumout[38]) );
  AND2X1 U16 ( .IN1(in2[31]), .IN2(in3[31]), .Q(cout[31]) );
  INVX0 U17 ( .INP(in2[31]), .ZN(n36) );
  MUX21X1 U18 ( .IN1(in2[31]), .IN2(n36), .S(in3[31]), .Q(sumout[31]) );
  AND2X1 U19 ( .IN1(in2[3]), .IN2(in1[3]), .Q(cout[3]) );
  AND2X1 U20 ( .IN1(in2[4]), .IN2(in1[4]), .Q(cout[4]) );
  NOR2X0 U21 ( .IN1(in2[4]), .IN2(in1[4]), .QN(n16) );
  NOR2X0 U22 ( .IN1(n16), .IN2(cout[4]), .QN(sumout[4]) );
  AND2X1 U23 ( .IN1(in2[5]), .IN2(in1[5]), .Q(cout[5]) );
  NOR2X0 U24 ( .IN1(in2[5]), .IN2(in1[5]), .QN(n17) );
  NOR2X0 U25 ( .IN1(n17), .IN2(cout[5]), .QN(sumout[5]) );
  AND2X1 U26 ( .IN1(in2[6]), .IN2(in1[6]), .Q(cout[6]) );
  NOR2X0 U27 ( .IN1(in2[6]), .IN2(in1[6]), .QN(n18) );
  NOR2X0 U28 ( .IN1(n18), .IN2(cout[6]), .QN(sumout[6]) );
  AND2X1 U29 ( .IN1(in2[7]), .IN2(in1[7]), .Q(cout[7]) );
  NOR2X0 U30 ( .IN1(in2[7]), .IN2(in1[7]), .QN(n19) );
  NOR2X0 U31 ( .IN1(n19), .IN2(cout[7]), .QN(sumout[7]) );
  AND2X1 U32 ( .IN1(in2[8]), .IN2(in1[8]), .Q(cout[8]) );
  NOR2X0 U33 ( .IN1(in2[8]), .IN2(in1[8]), .QN(n20) );
  NOR2X0 U34 ( .IN1(n20), .IN2(cout[8]), .QN(sumout[8]) );
  AND2X1 U35 ( .IN1(in2[9]), .IN2(in1[9]), .Q(cout[9]) );
  NOR2X0 U36 ( .IN1(in2[9]), .IN2(in1[9]), .QN(n21) );
  NOR2X0 U37 ( .IN1(n21), .IN2(cout[9]), .QN(sumout[9]) );
  AND2X1 U38 ( .IN1(in2[10]), .IN2(in1[10]), .Q(cout[10]) );
  NOR2X0 U39 ( .IN1(in2[10]), .IN2(in1[10]), .QN(n22) );
  NOR2X0 U40 ( .IN1(n22), .IN2(cout[10]), .QN(sumout[10]) );
  AND2X1 U41 ( .IN1(in2[11]), .IN2(in1[11]), .Q(cout[11]) );
  NOR2X0 U42 ( .IN1(in2[11]), .IN2(in1[11]), .QN(n23) );
  NOR2X0 U43 ( .IN1(n23), .IN2(cout[11]), .QN(sumout[11]) );
  AND2X1 U44 ( .IN1(in2[12]), .IN2(in1[12]), .Q(cout[12]) );
  NOR2X0 U45 ( .IN1(in2[12]), .IN2(in1[12]), .QN(n24) );
  NOR2X0 U46 ( .IN1(n24), .IN2(cout[12]), .QN(sumout[12]) );
  AND2X1 U47 ( .IN1(in2[13]), .IN2(in1[13]), .Q(cout[13]) );
  NOR2X0 U48 ( .IN1(in2[13]), .IN2(in1[13]), .QN(n25) );
  NOR2X0 U49 ( .IN1(n25), .IN2(cout[13]), .QN(sumout[13]) );
  AND2X1 U50 ( .IN1(in2[14]), .IN2(in1[14]), .Q(cout[14]) );
  NOR2X0 U51 ( .IN1(in2[14]), .IN2(in1[14]), .QN(n26) );
  NOR2X0 U52 ( .IN1(n26), .IN2(cout[14]), .QN(sumout[14]) );
  AND2X1 U53 ( .IN1(in2[15]), .IN2(in1[15]), .Q(cout[15]) );
  NOR2X0 U54 ( .IN1(in2[15]), .IN2(in1[15]), .QN(n27) );
  NOR2X0 U55 ( .IN1(n27), .IN2(cout[15]), .QN(sumout[15]) );
  AND2X1 U56 ( .IN1(in2[16]), .IN2(in1[16]), .Q(cout[16]) );
  NOR2X0 U57 ( .IN1(in2[16]), .IN2(in1[16]), .QN(n28) );
  NOR2X0 U58 ( .IN1(n28), .IN2(cout[16]), .QN(sumout[16]) );
  AND2X1 U59 ( .IN1(in2[17]), .IN2(in1[17]), .Q(cout[17]) );
  NOR2X0 U60 ( .IN1(in2[17]), .IN2(in1[17]), .QN(n29) );
  NOR2X0 U61 ( .IN1(n29), .IN2(cout[17]), .QN(sumout[17]) );
  AND2X1 U62 ( .IN1(in2[18]), .IN2(in1[18]), .Q(cout[18]) );
  NOR2X0 U63 ( .IN1(in2[18]), .IN2(in1[18]), .QN(n30) );
  NOR2X0 U64 ( .IN1(n30), .IN2(cout[18]), .QN(sumout[18]) );
  AND2X1 U65 ( .IN1(in2[19]), .IN2(in1[19]), .Q(cout[19]) );
  NOR2X0 U66 ( .IN1(in2[19]), .IN2(in1[19]), .QN(n31) );
  NOR2X0 U67 ( .IN1(n31), .IN2(cout[19]), .QN(sumout[19]) );
  AND2X1 U68 ( .IN1(in2[20]), .IN2(in1[20]), .Q(cout[20]) );
  NOR2X0 U69 ( .IN1(in2[20]), .IN2(in1[20]), .QN(n32) );
  NOR2X0 U70 ( .IN1(n32), .IN2(cout[20]), .QN(sumout[20]) );
  AND2X1 U71 ( .IN1(in2[21]), .IN2(in1[21]), .Q(cout[21]) );
  NOR2X0 U72 ( .IN1(in2[21]), .IN2(in1[21]), .QN(n33) );
  NOR2X0 U73 ( .IN1(n33), .IN2(cout[21]), .QN(sumout[21]) );
  AND2X1 U74 ( .IN1(in2[22]), .IN2(in1[22]), .Q(cout[22]) );
  NOR2X0 U75 ( .IN1(in2[22]), .IN2(in1[22]), .QN(n34) );
  NOR2X0 U76 ( .IN1(n34), .IN2(cout[22]), .QN(sumout[22]) );
  AND2X1 U77 ( .IN1(in2[23]), .IN2(in1[23]), .Q(cout[23]) );
  NOR2X0 U78 ( .IN1(in2[23]), .IN2(in1[23]), .QN(n35) );
  NOR2X0 U79 ( .IN1(n35), .IN2(cout[23]), .QN(sumout[23]) );
  FADDX1 U80 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U81 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U82 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U83 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U84 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U85 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U86 ( .A(in1[30]), .B(in3[30]), .CI(n36), .CO(cout[30]), .S(
        sumout[30]) );
endmodule


module csa51squ_45 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n3, n4, n5, n6, n7;

  NBUFFX2 U1 ( .INP(in1[18]), .Z(sumout[18]) );
  NBUFFX2 U2 ( .INP(in1[19]), .Z(sumout[19]) );
  AND2X1 U3 ( .IN1(in2[20]), .IN2(in1[20]), .Q(cout[20]) );
  NOR2X0 U4 ( .IN1(in2[20]), .IN2(in1[20]), .QN(n3) );
  NOR2X0 U5 ( .IN1(n3), .IN2(cout[20]), .QN(sumout[20]) );
  AND2X1 U6 ( .IN1(in2[21]), .IN2(in1[21]), .Q(cout[21]) );
  NOR2X0 U7 ( .IN1(in2[21]), .IN2(in1[21]), .QN(n4) );
  NOR2X0 U8 ( .IN1(n4), .IN2(cout[21]), .QN(sumout[21]) );
  AND2X1 U9 ( .IN1(in2[46]), .IN2(in3[46]), .Q(cout[46]) );
  NOR2X0 U10 ( .IN1(in2[46]), .IN2(in3[46]), .QN(n5) );
  NOR2X0 U11 ( .IN1(n5), .IN2(cout[46]), .QN(sumout[46]) );
  INVX0 U12 ( .INP(in2[46]), .ZN(n6) );
  MUX21X1 U13 ( .IN1(n6), .IN2(in2[46]), .S(in3[47]), .Q(sumout[47]) );
  INVX0 U14 ( .INP(in1[44]), .ZN(n7) );
  FADDX1 U15 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U16 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U17 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U18 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U19 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U20 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U21 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U22 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U23 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U24 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U25 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
  FADDX1 U26 ( .A(in1[33]), .B(in2[33]), .CI(in3[33]), .CO(cout[33]), .S(
        sumout[33]) );
  FADDX1 U27 ( .A(in1[34]), .B(in2[34]), .CI(in3[34]), .CO(cout[34]), .S(
        sumout[34]) );
  FADDX1 U28 ( .A(in1[35]), .B(in2[35]), .CI(in3[35]), .CO(cout[35]), .S(
        sumout[35]) );
  FADDX1 U29 ( .A(in1[36]), .B(in2[36]), .CI(in3[36]), .CO(cout[36]), .S(
        sumout[36]) );
  FADDX1 U30 ( .A(in1[37]), .B(in2[37]), .CI(in3[37]), .CO(cout[37]), .S(
        sumout[37]) );
  FADDX1 U31 ( .A(in1[38]), .B(in2[38]), .CI(in3[38]), .CO(cout[38]), .S(
        sumout[38]) );
  FADDX1 U32 ( .A(in1[39]), .B(in2[39]), .CI(in3[39]), .CO(cout[39]), .S(
        sumout[39]) );
  FADDX1 U33 ( .A(in1[40]), .B(in2[40]), .CI(in3[40]), .CO(cout[40]), .S(
        sumout[40]) );
  FADDX1 U34 ( .A(in1[41]), .B(in2[41]), .CI(in3[41]), .CO(cout[41]), .S(
        sumout[41]) );
  FADDX1 U35 ( .A(in1[42]), .B(in2[42]), .CI(in3[42]), .CO(cout[42]), .S(
        sumout[42]) );
  FADDX1 U36 ( .A(in1[43]), .B(in2[43]), .CI(in3[43]), .CO(cout[43]), .S(
        sumout[43]) );
  FADDX1 U37 ( .A(in1[44]), .B(in2[44]), .CI(in3[44]), .CO(cout[44]), .S(
        sumout[44]) );
  FADDX1 U38 ( .A(in2[45]), .B(in3[45]), .CI(n7), .CO(cout[45]), .S(sumout[45]) );
endmodule


module csa51squ_46 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n4, n5, n6, n7, n8;

  NBUFFX2 U1 ( .INP(in1[12]), .Z(sumout[12]) );
  NBUFFX2 U2 ( .INP(in1[13]), .Z(sumout[13]) );
  NBUFFX2 U3 ( .INP(in3[42]), .Z(sumout[42]) );
  AND2X1 U4 ( .IN1(in2[14]), .IN2(in1[14]), .Q(cout[14]) );
  NOR2X0 U5 ( .IN1(in2[14]), .IN2(in1[14]), .QN(n4) );
  NOR2X0 U6 ( .IN1(n4), .IN2(cout[14]), .QN(sumout[14]) );
  AND2X1 U7 ( .IN1(in2[15]), .IN2(in1[15]), .Q(cout[15]) );
  NOR2X0 U8 ( .IN1(in2[15]), .IN2(in1[15]), .QN(n5) );
  NOR2X0 U9 ( .IN1(n5), .IN2(cout[15]), .QN(sumout[15]) );
  AND2X1 U10 ( .IN1(in2[40]), .IN2(in3[40]), .Q(cout[40]) );
  NOR2X0 U11 ( .IN1(in2[40]), .IN2(in3[40]), .QN(n6) );
  NOR2X0 U12 ( .IN1(n6), .IN2(cout[40]), .QN(sumout[40]) );
  INVX0 U13 ( .INP(in3[41]), .ZN(n7) );
  NOR2X0 U14 ( .IN1(in2[40]), .IN2(n7), .QN(cout[41]) );
  MUX21X1 U15 ( .IN1(n7), .IN2(in3[41]), .S(in2[40]), .Q(sumout[41]) );
  INVX0 U16 ( .INP(in1[38]), .ZN(n8) );
  FADDX1 U17 ( .A(in1[16]), .B(in2[16]), .CI(in3[16]), .CO(cout[16]), .S(
        sumout[16]) );
  FADDX1 U18 ( .A(in1[17]), .B(in2[17]), .CI(in3[17]), .CO(cout[17]), .S(
        sumout[17]) );
  FADDX1 U19 ( .A(in1[18]), .B(in2[18]), .CI(in3[18]), .CO(cout[18]), .S(
        sumout[18]) );
  FADDX1 U20 ( .A(in1[19]), .B(in2[19]), .CI(in3[19]), .CO(cout[19]), .S(
        sumout[19]) );
  FADDX1 U21 ( .A(in1[20]), .B(in2[20]), .CI(in3[20]), .CO(cout[20]), .S(
        sumout[20]) );
  FADDX1 U22 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U23 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U24 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U25 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U26 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U27 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U28 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U29 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U30 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U31 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U32 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U33 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
  FADDX1 U34 ( .A(in1[33]), .B(in2[33]), .CI(in3[33]), .CO(cout[33]), .S(
        sumout[33]) );
  FADDX1 U35 ( .A(in1[34]), .B(in2[34]), .CI(in3[34]), .CO(cout[34]), .S(
        sumout[34]) );
  FADDX1 U36 ( .A(in1[35]), .B(in2[35]), .CI(in3[35]), .CO(cout[35]), .S(
        sumout[35]) );
  FADDX1 U37 ( .A(in1[36]), .B(in2[36]), .CI(in3[36]), .CO(cout[36]), .S(
        sumout[36]) );
  FADDX1 U38 ( .A(in1[37]), .B(in2[37]), .CI(in3[37]), .CO(cout[37]), .S(
        sumout[37]) );
  FADDX1 U39 ( .A(in1[38]), .B(in2[38]), .CI(in3[38]), .CO(cout[38]), .S(
        sumout[38]) );
  FADDX1 U40 ( .A(in2[39]), .B(in3[39]), .CI(n8), .CO(cout[39]), .S(sumout[39]) );
endmodule


module csa51squ_47 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n4, n5, n6, n7, n8;

  NBUFFX2 U1 ( .INP(in1[6]), .Z(sumout[6]) );
  NBUFFX2 U2 ( .INP(in1[7]), .Z(sumout[7]) );
  NBUFFX2 U3 ( .INP(in3[37]), .Z(sumout[37]) );
  AND2X1 U4 ( .IN1(in2[8]), .IN2(in1[8]), .Q(cout[8]) );
  NOR2X0 U5 ( .IN1(in2[8]), .IN2(in1[8]), .QN(n4) );
  NOR2X0 U6 ( .IN1(n4), .IN2(cout[8]), .QN(sumout[8]) );
  AND2X1 U7 ( .IN1(in2[9]), .IN2(in1[9]), .Q(cout[9]) );
  NOR2X0 U8 ( .IN1(in2[9]), .IN2(in1[9]), .QN(n5) );
  NOR2X0 U9 ( .IN1(n5), .IN2(cout[9]), .QN(sumout[9]) );
  AND2X1 U10 ( .IN1(in2[34]), .IN2(in3[34]), .Q(cout[34]) );
  NOR2X0 U11 ( .IN1(in2[34]), .IN2(in3[34]), .QN(n6) );
  NOR2X0 U12 ( .IN1(n6), .IN2(cout[34]), .QN(sumout[34]) );
  INVX0 U13 ( .INP(in3[35]), .ZN(n7) );
  NOR2X0 U14 ( .IN1(in2[34]), .IN2(n7), .QN(cout[35]) );
  MUX21X1 U15 ( .IN1(n7), .IN2(in3[35]), .S(in2[34]), .Q(sumout[35]) );
  INVX0 U16 ( .INP(in1[32]), .ZN(n8) );
  FADDX1 U17 ( .A(in1[10]), .B(in2[10]), .CI(in3[10]), .CO(cout[10]), .S(
        sumout[10]) );
  FADDX1 U18 ( .A(in1[11]), .B(in2[11]), .CI(in3[11]), .CO(cout[11]), .S(
        sumout[11]) );
  FADDX1 U19 ( .A(in1[12]), .B(in2[12]), .CI(in3[12]), .CO(cout[12]), .S(
        sumout[12]) );
  FADDX1 U20 ( .A(in1[13]), .B(in2[13]), .CI(in3[13]), .CO(cout[13]), .S(
        sumout[13]) );
  FADDX1 U21 ( .A(in1[14]), .B(in2[14]), .CI(in3[14]), .CO(cout[14]), .S(
        sumout[14]) );
  FADDX1 U22 ( .A(in1[15]), .B(in2[15]), .CI(in3[15]), .CO(cout[15]), .S(
        sumout[15]) );
  FADDX1 U23 ( .A(in1[16]), .B(in2[16]), .CI(in3[16]), .CO(cout[16]), .S(
        sumout[16]) );
  FADDX1 U24 ( .A(in1[17]), .B(in2[17]), .CI(in3[17]), .CO(cout[17]), .S(
        sumout[17]) );
  FADDX1 U25 ( .A(in1[18]), .B(in2[18]), .CI(in3[18]), .CO(cout[18]), .S(
        sumout[18]) );
  FADDX1 U26 ( .A(in1[19]), .B(in2[19]), .CI(in3[19]), .CO(cout[19]), .S(
        sumout[19]) );
  FADDX1 U27 ( .A(in1[20]), .B(in2[20]), .CI(in3[20]), .CO(cout[20]), .S(
        sumout[20]) );
  FADDX1 U28 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U29 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U30 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U31 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U32 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U33 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U34 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U35 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U36 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U37 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U38 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U39 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
  FADDX1 U40 ( .A(in2[33]), .B(in3[33]), .CI(n8), .CO(cout[33]), .S(sumout[33]) );
endmodule


module csa51squ_48 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n2, n3, n4, n5;

  NBUFFX2 U1 ( .INP(in3[31]), .Z(sumout[31]) );
  AND2X1 U2 ( .IN1(in2[2]), .IN2(in1[2]), .Q(cout[2]) );
  AND2X1 U3 ( .IN1(in2[3]), .IN2(in1[3]), .Q(cout[3]) );
  NOR2X0 U4 ( .IN1(in2[3]), .IN2(in1[3]), .QN(n2) );
  NOR2X0 U5 ( .IN1(n2), .IN2(cout[3]), .QN(sumout[3]) );
  AND2X1 U6 ( .IN1(in2[28]), .IN2(in3[28]), .Q(cout[28]) );
  NOR2X0 U7 ( .IN1(in2[28]), .IN2(in3[28]), .QN(n3) );
  NOR2X0 U8 ( .IN1(n3), .IN2(cout[28]), .QN(sumout[28]) );
  INVX0 U9 ( .INP(in3[29]), .ZN(n4) );
  NOR2X0 U10 ( .IN1(in2[28]), .IN2(n4), .QN(cout[29]) );
  MUX21X1 U11 ( .IN1(n4), .IN2(in3[29]), .S(in2[28]), .Q(sumout[29]) );
  INVX0 U12 ( .INP(in1[26]), .ZN(n5) );
  FADDX1 U13 ( .A(in1[10]), .B(in2[10]), .CI(in3[10]), .CO(cout[10]), .S(
        sumout[10]) );
  FADDX1 U14 ( .A(in1[11]), .B(in2[11]), .CI(in3[11]), .CO(cout[11]), .S(
        sumout[11]) );
  FADDX1 U15 ( .A(in1[12]), .B(in2[12]), .CI(in3[12]), .CO(cout[12]), .S(
        sumout[12]) );
  FADDX1 U16 ( .A(in1[13]), .B(in2[13]), .CI(in3[13]), .CO(cout[13]), .S(
        sumout[13]) );
  FADDX1 U17 ( .A(in1[14]), .B(in2[14]), .CI(in3[14]), .CO(cout[14]), .S(
        sumout[14]) );
  FADDX1 U18 ( .A(in1[15]), .B(in2[15]), .CI(in3[15]), .CO(cout[15]), .S(
        sumout[15]) );
  FADDX1 U19 ( .A(in1[16]), .B(in2[16]), .CI(in3[16]), .CO(cout[16]), .S(
        sumout[16]) );
  FADDX1 U20 ( .A(in1[17]), .B(in2[17]), .CI(in3[17]), .CO(cout[17]), .S(
        sumout[17]) );
  FADDX1 U21 ( .A(in1[18]), .B(in2[18]), .CI(in3[18]), .CO(cout[18]), .S(
        sumout[18]) );
  FADDX1 U22 ( .A(in1[19]), .B(in2[19]), .CI(in3[19]), .CO(cout[19]), .S(
        sumout[19]) );
  FADDX1 U23 ( .A(in1[20]), .B(in2[20]), .CI(in3[20]), .CO(cout[20]), .S(
        sumout[20]) );
  FADDX1 U24 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U25 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U26 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U27 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U28 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U29 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U30 ( .A(in2[27]), .B(in3[27]), .CI(n5), .CO(cout[27]), .S(sumout[27]) );
  FADDX1 U31 ( .A(in1[4]), .B(in2[4]), .CI(in3[4]), .CO(cout[4]), .S(sumout[4]) );
  FADDX1 U32 ( .A(in1[5]), .B(in2[5]), .CI(in3[5]), .CO(cout[5]), .S(sumout[5]) );
  FADDX1 U33 ( .A(in1[6]), .B(in2[6]), .CI(in3[6]), .CO(cout[6]), .S(sumout[6]) );
  FADDX1 U34 ( .A(in1[7]), .B(in2[7]), .CI(in3[7]), .CO(cout[7]), .S(sumout[7]) );
  FADDX1 U35 ( .A(in1[8]), .B(in2[8]), .CI(in3[8]), .CO(cout[8]), .S(sumout[8]) );
  FADDX1 U36 ( .A(in1[9]), .B(in2[9]), .CI(in3[9]), .CO(cout[9]), .S(sumout[9]) );
endmodule


module booth27_40 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;


  NBUFFX2 U3 ( .INP(in2[22]), .Z(out1[22]) );
  NBUFFX2 U4 ( .INP(in2[21]), .Z(out1[21]) );
  NBUFFX2 U5 ( .INP(in2[20]), .Z(out1[20]) );
  NBUFFX2 U6 ( .INP(in2[0]), .Z(out1[0]) );
  NBUFFX2 U7 ( .INP(in2[19]), .Z(out1[19]) );
  NBUFFX2 U8 ( .INP(in2[18]), .Z(out1[18]) );
  NBUFFX2 U9 ( .INP(in2[2]), .Z(out1[2]) );
  NBUFFX2 U10 ( .INP(in2[1]), .Z(out1[1]) );
  NBUFFX2 U11 ( .INP(in2[4]), .Z(out1[4]) );
  NBUFFX2 U12 ( .INP(in2[3]), .Z(out1[3]) );
  NBUFFX2 U13 ( .INP(in2[6]), .Z(out1[6]) );
  NBUFFX2 U14 ( .INP(in2[5]), .Z(out1[5]) );
  NBUFFX2 U15 ( .INP(in2[9]), .Z(out1[9]) );
  NBUFFX2 U16 ( .INP(in2[8]), .Z(out1[8]) );
  NBUFFX2 U17 ( .INP(in2[7]), .Z(out1[7]) );
  NBUFFX2 U18 ( .INP(in2[13]), .Z(out1[13]) );
  NBUFFX2 U19 ( .INP(in2[12]), .Z(out1[12]) );
  NBUFFX2 U20 ( .INP(in2[11]), .Z(out1[11]) );
  NBUFFX2 U21 ( .INP(in2[10]), .Z(out1[10]) );
  NBUFFX2 U22 ( .INP(in2[17]), .Z(out1[17]) );
  NBUFFX2 U23 ( .INP(in2[16]), .Z(out1[16]) );
  NBUFFX2 U24 ( .INP(in2[15]), .Z(out1[15]) );
  NBUFFX2 U25 ( .INP(in2[14]), .Z(out1[14]) );
endmodule


module booth27_41 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76;

  NAND2X0 U3 ( .IN1(n1), .IN2(n2), .QN(n8) );
  NAND2X0 U4 ( .IN1(n71), .IN2(in2[0]), .QN(n15) );
  NAND2X0 U5 ( .IN1(n19), .IN2(in2[5]), .QN(n20) );
  NAND2X0 U6 ( .IN1(n25), .IN2(in2[7]), .QN(n26) );
  NAND2X0 U7 ( .IN1(n31), .IN2(in2[9]), .QN(n32) );
  NAND2X0 U8 ( .IN1(n37), .IN2(in2[11]), .QN(n38) );
  NAND2X0 U9 ( .IN1(n43), .IN2(in2[13]), .QN(n44) );
  NAND2X0 U10 ( .IN1(n46), .IN2(in2[14]), .QN(n47) );
  NAND2X0 U11 ( .IN1(n49), .IN2(in2[15]), .QN(n50) );
  NAND2X0 U12 ( .IN1(n52), .IN2(in2[16]), .QN(n53) );
  NAND2X0 U13 ( .IN1(n55), .IN2(in2[17]), .QN(n56) );
  NAND2X0 U14 ( .IN1(n7), .IN2(n15), .QN(out1[1]) );
  NAND2X0 U15 ( .IN1(n10), .IN2(n9), .QN(out1[2]) );
  NAND2X0 U16 ( .IN1(n58), .IN2(in2[18]), .QN(n59) );
  NAND2X0 U17 ( .IN1(n61), .IN2(in2[19]), .QN(n62) );
  NAND2X0 U18 ( .IN1(in1[1]), .IN2(in1[0]), .QN(out1[25]) );
  NOR2X0 U19 ( .IN1(in1[1]), .IN2(in1[0]), .QN(n71) );
  INVX0 U20 ( .INP(in2[0]), .ZN(n1) );
  INVX0 U21 ( .INP(in2[1]), .ZN(n2) );
  INVX0 U22 ( .INP(in2[3]), .ZN(n3) );
  INVX0 U23 ( .INP(in2[21]), .ZN(n4) );
  INVX0 U24 ( .INP(in2[22]), .ZN(n5) );
  INVX0 U25 ( .INP(in1[1]), .ZN(n6) );
  MUX21X1 U26 ( .IN1(in1[1]), .IN2(n6), .S(in1[0]), .Q(n74) );
  INVX0 U27 ( .INP(n74), .ZN(n76) );
  AO221X1 U28 ( .IN1(in2[0]), .IN2(in2[1]), .IN3(n1), .IN4(n2), .IN5(n76), .Q(
        n7) );
  MUX21X1 U29 ( .IN1(n2), .IN2(n8), .S(in2[2]), .Q(n12) );
  AO221X1 U30 ( .IN1(n12), .IN2(in2[2]), .IN3(n12), .IN4(n1), .IN5(n76), .Q(
        n10) );
  INVX0 U31 ( .INP(n71), .ZN(n13) );
  AO221X1 U32 ( .IN1(in2[0]), .IN2(in2[1]), .IN3(n1), .IN4(n2), .IN5(n13), .Q(
        n9) );
  NOR3X0 U33 ( .IN1(in2[0]), .IN2(in2[2]), .IN3(in2[1]), .QN(n11) );
  OR4X1 U34 ( .IN1(in2[3]), .IN2(in2[0]), .IN3(in2[2]), .IN4(in2[1]), .Q(n16)
         );
  OA21X1 U35 ( .IN1(n11), .IN2(n3), .IN3(n16), .Q(n18) );
  INVX0 U36 ( .INP(n18), .ZN(n14) );
  OAI222X1 U37 ( .IN1(n15), .IN2(in2[2]), .IN3(n14), .IN4(n76), .IN5(n13), 
        .IN6(n12), .QN(out1[3]) );
  OR2X1 U38 ( .IN1(in2[4]), .IN2(n16), .Q(n19) );
  NAND2X0 U39 ( .IN1(n16), .IN2(in2[4]), .QN(n17) );
  AND2X1 U40 ( .IN1(n19), .IN2(n17), .Q(n21) );
  AO22X1 U41 ( .IN1(n71), .IN2(n18), .IN3(n21), .IN4(n74), .Q(out1[4]) );
  OR2X1 U42 ( .IN1(in2[5]), .IN2(n19), .Q(n22) );
  AND2X1 U43 ( .IN1(n22), .IN2(n20), .Q(n24) );
  AO22X1 U44 ( .IN1(n71), .IN2(n21), .IN3(n24), .IN4(n74), .Q(out1[5]) );
  OR2X1 U45 ( .IN1(in2[6]), .IN2(n22), .Q(n25) );
  NAND2X0 U46 ( .IN1(n22), .IN2(in2[6]), .QN(n23) );
  AND2X1 U47 ( .IN1(n25), .IN2(n23), .Q(n27) );
  AO22X1 U48 ( .IN1(n71), .IN2(n24), .IN3(n27), .IN4(n74), .Q(out1[6]) );
  OR2X1 U49 ( .IN1(in2[7]), .IN2(n25), .Q(n28) );
  AND2X1 U50 ( .IN1(n28), .IN2(n26), .Q(n30) );
  AO22X1 U51 ( .IN1(n71), .IN2(n27), .IN3(n30), .IN4(n74), .Q(out1[7]) );
  OR2X1 U52 ( .IN1(in2[8]), .IN2(n28), .Q(n31) );
  NAND2X0 U53 ( .IN1(n28), .IN2(in2[8]), .QN(n29) );
  AND2X1 U54 ( .IN1(n31), .IN2(n29), .Q(n33) );
  AO22X1 U55 ( .IN1(n71), .IN2(n30), .IN3(n33), .IN4(n74), .Q(out1[8]) );
  OR2X1 U56 ( .IN1(in2[9]), .IN2(n31), .Q(n34) );
  AND2X1 U57 ( .IN1(n34), .IN2(n32), .Q(n36) );
  AO22X1 U58 ( .IN1(n71), .IN2(n33), .IN3(n36), .IN4(n74), .Q(out1[9]) );
  OR2X1 U59 ( .IN1(in2[10]), .IN2(n34), .Q(n37) );
  NAND2X0 U60 ( .IN1(n34), .IN2(in2[10]), .QN(n35) );
  AND2X1 U61 ( .IN1(n37), .IN2(n35), .Q(n39) );
  AO22X1 U62 ( .IN1(n71), .IN2(n36), .IN3(n39), .IN4(n74), .Q(out1[10]) );
  OR2X1 U63 ( .IN1(in2[11]), .IN2(n37), .Q(n40) );
  AND2X1 U64 ( .IN1(n40), .IN2(n38), .Q(n42) );
  AO22X1 U65 ( .IN1(n71), .IN2(n39), .IN3(n42), .IN4(n74), .Q(out1[11]) );
  OR2X1 U66 ( .IN1(in2[12]), .IN2(n40), .Q(n43) );
  NAND2X0 U67 ( .IN1(n40), .IN2(in2[12]), .QN(n41) );
  AND2X1 U68 ( .IN1(n43), .IN2(n41), .Q(n45) );
  AO22X1 U69 ( .IN1(n71), .IN2(n42), .IN3(n45), .IN4(n74), .Q(out1[12]) );
  OR2X1 U70 ( .IN1(in2[13]), .IN2(n43), .Q(n46) );
  AND2X1 U71 ( .IN1(n46), .IN2(n44), .Q(n48) );
  AO22X1 U72 ( .IN1(n71), .IN2(n45), .IN3(n48), .IN4(n74), .Q(out1[13]) );
  OR2X1 U73 ( .IN1(in2[14]), .IN2(n46), .Q(n49) );
  AND2X1 U74 ( .IN1(n49), .IN2(n47), .Q(n51) );
  AO22X1 U75 ( .IN1(n71), .IN2(n48), .IN3(n51), .IN4(n74), .Q(out1[14]) );
  OR2X1 U76 ( .IN1(in2[15]), .IN2(n49), .Q(n52) );
  AND2X1 U77 ( .IN1(n52), .IN2(n50), .Q(n54) );
  AO22X1 U78 ( .IN1(n71), .IN2(n51), .IN3(n54), .IN4(n74), .Q(out1[15]) );
  OR2X1 U79 ( .IN1(in2[16]), .IN2(n52), .Q(n55) );
  AND2X1 U80 ( .IN1(n55), .IN2(n53), .Q(n57) );
  AO22X1 U81 ( .IN1(n71), .IN2(n54), .IN3(n57), .IN4(n74), .Q(out1[16]) );
  OR2X1 U82 ( .IN1(in2[17]), .IN2(n55), .Q(n58) );
  AND2X1 U83 ( .IN1(n58), .IN2(n56), .Q(n60) );
  AO22X1 U84 ( .IN1(n71), .IN2(n57), .IN3(n60), .IN4(n74), .Q(out1[17]) );
  OR2X1 U85 ( .IN1(in2[18]), .IN2(n58), .Q(n61) );
  AND2X1 U86 ( .IN1(n61), .IN2(n59), .Q(n63) );
  AO22X1 U87 ( .IN1(n71), .IN2(n60), .IN3(n63), .IN4(n74), .Q(out1[18]) );
  OR2X1 U88 ( .IN1(in2[19]), .IN2(n61), .Q(n64) );
  AND2X1 U89 ( .IN1(n64), .IN2(n62), .Q(n65) );
  AO22X1 U90 ( .IN1(n71), .IN2(n63), .IN3(n65), .IN4(n74), .Q(out1[19]) );
  NOR2X0 U91 ( .IN1(in2[20]), .IN2(n64), .QN(n72) );
  AOI21X1 U92 ( .IN1(in2[20]), .IN2(n64), .IN3(n72), .QN(n66) );
  AO22X1 U93 ( .IN1(n71), .IN2(n65), .IN3(n66), .IN4(n74), .Q(out1[20]) );
  MUX21X1 U94 ( .IN1(n4), .IN2(in2[21]), .S(n72), .Q(n69) );
  AO22X1 U95 ( .IN1(n71), .IN2(n66), .IN3(n69), .IN4(n74), .Q(out1[21]) );
  INVX0 U96 ( .INP(n72), .ZN(n67) );
  NOR2X0 U97 ( .IN1(in2[21]), .IN2(n67), .QN(n70) );
  MUX21X1 U98 ( .IN1(n5), .IN2(in2[22]), .S(n70), .Q(n68) );
  AO22X1 U99 ( .IN1(n71), .IN2(n69), .IN3(n68), .IN4(n74), .Q(out1[22]) );
  MUX21X1 U100 ( .IN1(n71), .IN2(n74), .S(n70), .Q(n73) );
  AND3X1 U101 ( .IN1(n72), .IN2(n71), .IN3(n4), .Q(n75) );
  MUX21X1 U102 ( .IN1(n73), .IN2(n75), .S(in2[22]), .Q(out1[23]) );
  AO21X1 U103 ( .IN1(n75), .IN2(n5), .IN3(n74), .Q(out1[24]) );
  NOR2X0 U104 ( .IN1(n76), .IN2(n1), .QN(out1[0]) );
endmodule


module booth27_42 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n25), .IN2(n6), .QN(n30) );
  NAND2X0 U4 ( .IN1(n33), .IN2(n7), .QN(n37) );
  NAND2X0 U5 ( .IN1(n41), .IN2(n8), .QN(n45) );
  NAND2X0 U6 ( .IN1(n49), .IN2(n9), .QN(n53) );
  NAND2X0 U7 ( .IN1(n57), .IN2(n10), .QN(n61) );
  NAND2X0 U8 ( .IN1(n65), .IN2(n11), .QN(n77) );
  NAND2X0 U9 ( .IN1(n81), .IN2(n13), .QN(n89) );
  NAND2X0 U10 ( .IN1(n93), .IN2(n15), .QN(n101) );
  NAND2X0 U11 ( .IN1(n105), .IN2(n17), .QN(n114) );
  NAND2X0 U12 ( .IN1(n27), .IN2(n132), .QN(n4) );
  NAND2X0 U13 ( .IN1(in1[2]), .IN2(n77), .QN(n71) );
  NAND2X0 U14 ( .IN1(n70), .IN2(n132), .QN(n74) );
  NAND2X0 U15 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U16 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U17 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U18 ( .IN1(n118), .IN2(n19), .QN(n125) );
  NAND2X0 U19 ( .IN1(n141), .IN2(n130), .QN(n24) );
  NAND2X0 U20 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NAND2X0 U21 ( .IN1(n32), .IN2(n31), .QN(out1[3]) );
  NAND2X0 U22 ( .IN1(n36), .IN2(n35), .QN(out1[4]) );
  NAND2X0 U23 ( .IN1(n40), .IN2(n39), .QN(out1[5]) );
  NAND2X0 U24 ( .IN1(n44), .IN2(n43), .QN(out1[6]) );
  NAND2X0 U25 ( .IN1(n48), .IN2(n47), .QN(out1[7]) );
  NAND2X0 U26 ( .IN1(n52), .IN2(n51), .QN(out1[8]) );
  NAND2X0 U27 ( .IN1(n56), .IN2(n55), .QN(out1[9]) );
  NAND2X0 U28 ( .IN1(n60), .IN2(n59), .QN(out1[10]) );
  NAND2X0 U29 ( .IN1(n64), .IN2(n63), .QN(out1[11]) );
  NAND2X0 U30 ( .IN1(n69), .IN2(n68), .QN(out1[12]) );
  NAND2X0 U31 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U32 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U33 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U34 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U35 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U36 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U37 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U38 ( .IN1(n23), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U39 ( .IN1(in1[2]), .IN2(n22), .QN(n23) );
  NOR2X0 U40 ( .IN1(n28), .IN2(n26), .QN(n3) );
  NOR2X0 U41 ( .IN1(n142), .IN2(n21), .QN(n1) );
  NOR2X0 U42 ( .IN1(n142), .IN2(n111), .QN(n138) );
  INVX0 U43 ( .INP(n130), .ZN(n137) );
  INVX0 U44 ( .INP(n132), .ZN(n141) );
  NOR3X0 U45 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  NAND3X0 U46 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  MUX21X1 U47 ( .IN1(n22), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  INVX0 U48 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U49 ( .INP(in2[2]), .ZN(n6) );
  INVX0 U50 ( .INP(in2[4]), .ZN(n7) );
  INVX0 U51 ( .INP(in2[6]), .ZN(n8) );
  INVX0 U52 ( .INP(in2[8]), .ZN(n9) );
  INVX0 U53 ( .INP(in2[10]), .ZN(n10) );
  INVX0 U54 ( .INP(in2[12]), .ZN(n11) );
  INVX0 U55 ( .INP(in2[13]), .ZN(n12) );
  INVX0 U56 ( .INP(in2[14]), .ZN(n13) );
  INVX0 U57 ( .INP(in2[15]), .ZN(n14) );
  INVX0 U58 ( .INP(in2[16]), .ZN(n15) );
  INVX0 U59 ( .INP(in2[17]), .ZN(n16) );
  INVX0 U60 ( .INP(in2[18]), .ZN(n17) );
  INVX0 U61 ( .INP(in2[19]), .ZN(n18) );
  INVX0 U62 ( .INP(in2[20]), .ZN(n19) );
  INVX0 U63 ( .INP(in2[21]), .ZN(n20) );
  INVX0 U64 ( .INP(in2[22]), .ZN(n21) );
  INVX0 U65 ( .INP(in1[1]), .ZN(n22) );
  INVX0 U66 ( .INP(in1[2]), .ZN(n111) );
  INVX0 U67 ( .INP(n138), .ZN(n140) );
  NOR2X0 U68 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n25) );
  AOI21X1 U69 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n25), .QN(n27) );
  NOR2X0 U70 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U71 ( .IN1(n24), .IN2(in2[0]), .IN3(n138), .IN4(n27), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U72 ( .INP(n133), .ZN(n67) );
  NOR2X0 U73 ( .IN1(n67), .IN2(n6), .QN(n28) );
  OA21X1 U74 ( .IN1(n25), .IN2(n6), .IN3(n30), .Q(n29) );
  AO22X1 U75 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n29), .Q(n26) );
  AOI22X1 U76 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n29), .QN(n32) );
  NOR2X0 U77 ( .IN1(in2[3]), .IN2(n30), .QN(n33) );
  AO21X1 U78 ( .IN1(in2[3]), .IN2(n30), .IN3(n33), .Q(n34) );
  OA22X1 U79 ( .IN1(n6), .IN2(n130), .IN3(n140), .IN4(n34), .Q(n31) );
  OA21X1 U80 ( .IN1(n33), .IN2(n7), .IN3(n37), .Q(n38) );
  AOI22X1 U81 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n38), .QN(n36) );
  OA22X1 U82 ( .IN1(n67), .IN2(n7), .IN3(n141), .IN4(n34), .Q(n35) );
  NOR2X0 U83 ( .IN1(in2[5]), .IN2(n37), .QN(n41) );
  AO21X1 U84 ( .IN1(in2[5]), .IN2(n37), .IN3(n41), .Q(n42) );
  OA22X1 U85 ( .IN1(n7), .IN2(n130), .IN3(n140), .IN4(n42), .Q(n40) );
  AOI22X1 U86 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n38), .QN(n39) );
  OA21X1 U87 ( .IN1(n41), .IN2(n8), .IN3(n45), .Q(n46) );
  AOI22X1 U88 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n46), .QN(n44) );
  OA22X1 U89 ( .IN1(n67), .IN2(n8), .IN3(n141), .IN4(n42), .Q(n43) );
  NOR2X0 U90 ( .IN1(in2[7]), .IN2(n45), .QN(n49) );
  AO21X1 U91 ( .IN1(in2[7]), .IN2(n45), .IN3(n49), .Q(n50) );
  OA22X1 U92 ( .IN1(n8), .IN2(n130), .IN3(n140), .IN4(n50), .Q(n48) );
  AOI22X1 U93 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n46), .QN(n47) );
  OA21X1 U94 ( .IN1(n49), .IN2(n9), .IN3(n53), .Q(n54) );
  AOI22X1 U95 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n54), .QN(n52) );
  OA22X1 U96 ( .IN1(n67), .IN2(n9), .IN3(n141), .IN4(n50), .Q(n51) );
  NOR2X0 U97 ( .IN1(in2[9]), .IN2(n53), .QN(n57) );
  AO21X1 U98 ( .IN1(in2[9]), .IN2(n53), .IN3(n57), .Q(n58) );
  OA22X1 U99 ( .IN1(n9), .IN2(n130), .IN3(n140), .IN4(n58), .Q(n56) );
  AOI22X1 U100 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n54), .QN(n55) );
  OA21X1 U101 ( .IN1(n57), .IN2(n10), .IN3(n61), .Q(n62) );
  AOI22X1 U102 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n62), .QN(n60) );
  OA22X1 U103 ( .IN1(n67), .IN2(n10), .IN3(n141), .IN4(n58), .Q(n59) );
  NOR2X0 U104 ( .IN1(in2[11]), .IN2(n61), .QN(n65) );
  AO21X1 U105 ( .IN1(in2[11]), .IN2(n61), .IN3(n65), .Q(n66) );
  OA22X1 U106 ( .IN1(n10), .IN2(n130), .IN3(n140), .IN4(n66), .Q(n64) );
  AOI22X1 U107 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n62), .QN(n63) );
  OA21X1 U108 ( .IN1(n65), .IN2(n11), .IN3(n77), .Q(n70) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n70), .QN(n69) );
  OA22X1 U110 ( .IN1(n67), .IN2(n11), .IN3(n141), .IN4(n66), .Q(n68) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n12), .S(n71), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n11), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n13), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n12), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n12), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n14), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n13), .IN4(n85), .IN5(n84), 
        .Q(out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n15), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n14), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n14), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n16), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n15), .IN4(n97), .IN5(n96), 
        .Q(out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n17), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n16), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n16), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n18), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n17), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n19), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n18), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n18), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n20), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n19), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n21), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n20), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n20), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n21), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_43 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n33), .IN2(n7), .QN(n37) );
  NAND2X0 U4 ( .IN1(n41), .IN2(n8), .QN(n45) );
  NAND2X0 U5 ( .IN1(n49), .IN2(n9), .QN(n53) );
  NAND2X0 U6 ( .IN1(n57), .IN2(n10), .QN(n61) );
  NAND2X0 U7 ( .IN1(n25), .IN2(n6), .QN(n30) );
  NAND2X0 U8 ( .IN1(n65), .IN2(n11), .QN(n77) );
  NAND2X0 U9 ( .IN1(n81), .IN2(n13), .QN(n89) );
  NAND2X0 U10 ( .IN1(n93), .IN2(n15), .QN(n101) );
  NAND2X0 U11 ( .IN1(n105), .IN2(n17), .QN(n114) );
  NAND2X0 U12 ( .IN1(n118), .IN2(n19), .QN(n125) );
  NAND2X0 U13 ( .IN1(in1[2]), .IN2(n77), .QN(n71) );
  NAND2X0 U14 ( .IN1(n70), .IN2(n132), .QN(n74) );
  NAND2X0 U15 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U16 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U17 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U18 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U19 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U20 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U21 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U22 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NAND2X0 U23 ( .IN1(n27), .IN2(n132), .QN(n4) );
  NAND2X0 U24 ( .IN1(n32), .IN2(n31), .QN(out1[3]) );
  NAND2X0 U25 ( .IN1(n36), .IN2(n35), .QN(out1[4]) );
  NAND2X0 U26 ( .IN1(n40), .IN2(n39), .QN(out1[5]) );
  NAND2X0 U27 ( .IN1(n44), .IN2(n43), .QN(out1[6]) );
  NAND2X0 U28 ( .IN1(n48), .IN2(n47), .QN(out1[7]) );
  NAND2X0 U29 ( .IN1(n52), .IN2(n51), .QN(out1[8]) );
  NAND2X0 U30 ( .IN1(n56), .IN2(n55), .QN(out1[9]) );
  NAND2X0 U31 ( .IN1(n60), .IN2(n59), .QN(out1[10]) );
  NAND2X0 U32 ( .IN1(n64), .IN2(n63), .QN(out1[11]) );
  NAND2X0 U33 ( .IN1(n69), .IN2(n68), .QN(out1[12]) );
  NAND2X0 U34 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U35 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U36 ( .IN1(n141), .IN2(n130), .QN(n24) );
  NAND2X0 U37 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U38 ( .IN1(n23), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U39 ( .IN1(in1[2]), .IN2(n22), .QN(n23) );
  NOR2X0 U40 ( .IN1(n28), .IN2(n26), .QN(n3) );
  NOR2X0 U41 ( .IN1(n142), .IN2(n111), .QN(n138) );
  NOR2X0 U42 ( .IN1(n142), .IN2(n21), .QN(n1) );
  INVX0 U43 ( .INP(n130), .ZN(n137) );
  INVX0 U44 ( .INP(n132), .ZN(n141) );
  NOR3X0 U45 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  NAND3X0 U46 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  MUX21X1 U47 ( .IN1(n22), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  INVX0 U48 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U49 ( .INP(in2[2]), .ZN(n6) );
  INVX0 U50 ( .INP(in2[4]), .ZN(n7) );
  INVX0 U51 ( .INP(in2[6]), .ZN(n8) );
  INVX0 U52 ( .INP(in2[8]), .ZN(n9) );
  INVX0 U53 ( .INP(in2[10]), .ZN(n10) );
  INVX0 U54 ( .INP(in2[12]), .ZN(n11) );
  INVX0 U55 ( .INP(in2[13]), .ZN(n12) );
  INVX0 U56 ( .INP(in2[14]), .ZN(n13) );
  INVX0 U57 ( .INP(in2[15]), .ZN(n14) );
  INVX0 U58 ( .INP(in2[16]), .ZN(n15) );
  INVX0 U59 ( .INP(in2[17]), .ZN(n16) );
  INVX0 U60 ( .INP(in2[18]), .ZN(n17) );
  INVX0 U61 ( .INP(in2[19]), .ZN(n18) );
  INVX0 U62 ( .INP(in2[20]), .ZN(n19) );
  INVX0 U63 ( .INP(in2[21]), .ZN(n20) );
  INVX0 U64 ( .INP(in2[22]), .ZN(n21) );
  INVX0 U65 ( .INP(in1[1]), .ZN(n22) );
  INVX0 U66 ( .INP(in1[2]), .ZN(n111) );
  INVX0 U67 ( .INP(n138), .ZN(n140) );
  NOR2X0 U68 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n25) );
  AOI21X1 U69 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n25), .QN(n27) );
  NOR2X0 U70 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U71 ( .IN1(n24), .IN2(in2[0]), .IN3(n138), .IN4(n27), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U72 ( .INP(n133), .ZN(n67) );
  NOR2X0 U73 ( .IN1(n67), .IN2(n6), .QN(n28) );
  OA21X1 U74 ( .IN1(n25), .IN2(n6), .IN3(n30), .Q(n29) );
  AO22X1 U75 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n29), .Q(n26) );
  AOI22X1 U76 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n29), .QN(n32) );
  NOR2X0 U77 ( .IN1(in2[3]), .IN2(n30), .QN(n33) );
  AO21X1 U78 ( .IN1(in2[3]), .IN2(n30), .IN3(n33), .Q(n34) );
  OA22X1 U79 ( .IN1(n6), .IN2(n130), .IN3(n140), .IN4(n34), .Q(n31) );
  OA21X1 U80 ( .IN1(n33), .IN2(n7), .IN3(n37), .Q(n38) );
  AOI22X1 U81 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n38), .QN(n36) );
  OA22X1 U82 ( .IN1(n67), .IN2(n7), .IN3(n141), .IN4(n34), .Q(n35) );
  NOR2X0 U83 ( .IN1(in2[5]), .IN2(n37), .QN(n41) );
  AO21X1 U84 ( .IN1(in2[5]), .IN2(n37), .IN3(n41), .Q(n42) );
  OA22X1 U85 ( .IN1(n7), .IN2(n130), .IN3(n140), .IN4(n42), .Q(n40) );
  AOI22X1 U86 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n38), .QN(n39) );
  OA21X1 U87 ( .IN1(n41), .IN2(n8), .IN3(n45), .Q(n46) );
  AOI22X1 U88 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n46), .QN(n44) );
  OA22X1 U89 ( .IN1(n67), .IN2(n8), .IN3(n141), .IN4(n42), .Q(n43) );
  NOR2X0 U90 ( .IN1(in2[7]), .IN2(n45), .QN(n49) );
  AO21X1 U91 ( .IN1(in2[7]), .IN2(n45), .IN3(n49), .Q(n50) );
  OA22X1 U92 ( .IN1(n8), .IN2(n130), .IN3(n140), .IN4(n50), .Q(n48) );
  AOI22X1 U93 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n46), .QN(n47) );
  OA21X1 U94 ( .IN1(n49), .IN2(n9), .IN3(n53), .Q(n54) );
  AOI22X1 U95 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n54), .QN(n52) );
  OA22X1 U96 ( .IN1(n67), .IN2(n9), .IN3(n141), .IN4(n50), .Q(n51) );
  NOR2X0 U97 ( .IN1(in2[9]), .IN2(n53), .QN(n57) );
  AO21X1 U98 ( .IN1(in2[9]), .IN2(n53), .IN3(n57), .Q(n58) );
  OA22X1 U99 ( .IN1(n9), .IN2(n130), .IN3(n140), .IN4(n58), .Q(n56) );
  AOI22X1 U100 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n54), .QN(n55) );
  OA21X1 U101 ( .IN1(n57), .IN2(n10), .IN3(n61), .Q(n62) );
  AOI22X1 U102 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n62), .QN(n60) );
  OA22X1 U103 ( .IN1(n67), .IN2(n10), .IN3(n141), .IN4(n58), .Q(n59) );
  NOR2X0 U104 ( .IN1(in2[11]), .IN2(n61), .QN(n65) );
  AO21X1 U105 ( .IN1(in2[11]), .IN2(n61), .IN3(n65), .Q(n66) );
  OA22X1 U106 ( .IN1(n10), .IN2(n130), .IN3(n140), .IN4(n66), .Q(n64) );
  AOI22X1 U107 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n62), .QN(n63) );
  OA21X1 U108 ( .IN1(n65), .IN2(n11), .IN3(n77), .Q(n70) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n70), .QN(n69) );
  OA22X1 U110 ( .IN1(n67), .IN2(n11), .IN3(n141), .IN4(n66), .Q(n68) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n12), .S(n71), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n11), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n13), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n12), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n12), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n14), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n13), .IN4(n85), .IN5(n84), 
        .Q(out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n15), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n14), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n14), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n16), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n15), .IN4(n97), .IN5(n96), 
        .Q(out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n17), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n16), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n16), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n18), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n17), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n19), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n18), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n18), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n20), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n19), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n21), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n20), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n20), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n21), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_44 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n41), .IN2(n8), .QN(n45) );
  NAND2X0 U4 ( .IN1(n49), .IN2(n9), .QN(n53) );
  NAND2X0 U5 ( .IN1(n57), .IN2(n10), .QN(n61) );
  NAND2X0 U6 ( .IN1(n33), .IN2(n7), .QN(n37) );
  NAND2X0 U7 ( .IN1(n25), .IN2(n6), .QN(n30) );
  NAND2X0 U8 ( .IN1(n65), .IN2(n11), .QN(n77) );
  NAND2X0 U9 ( .IN1(n81), .IN2(n13), .QN(n89) );
  NAND2X0 U10 ( .IN1(n93), .IN2(n15), .QN(n101) );
  NAND2X0 U11 ( .IN1(in1[2]), .IN2(n77), .QN(n71) );
  NAND2X0 U12 ( .IN1(n70), .IN2(n132), .QN(n74) );
  NAND2X0 U13 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U14 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U15 ( .IN1(n105), .IN2(n17), .QN(n114) );
  NAND2X0 U16 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U17 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U18 ( .IN1(n27), .IN2(n132), .QN(n4) );
  NAND2X0 U19 ( .IN1(n141), .IN2(n130), .QN(n24) );
  NAND2X0 U20 ( .IN1(n40), .IN2(n39), .QN(out1[5]) );
  NAND2X0 U21 ( .IN1(n44), .IN2(n43), .QN(out1[6]) );
  NAND2X0 U22 ( .IN1(n48), .IN2(n47), .QN(out1[7]) );
  NAND2X0 U23 ( .IN1(n52), .IN2(n51), .QN(out1[8]) );
  NAND2X0 U24 ( .IN1(n56), .IN2(n55), .QN(out1[9]) );
  NAND2X0 U25 ( .IN1(n60), .IN2(n59), .QN(out1[10]) );
  NAND2X0 U26 ( .IN1(n64), .IN2(n63), .QN(out1[11]) );
  NAND2X0 U27 ( .IN1(n69), .IN2(n68), .QN(out1[12]) );
  NAND2X0 U28 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U29 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U30 ( .IN1(n118), .IN2(n19), .QN(n125) );
  NAND2X0 U31 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U32 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U33 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U34 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U35 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NAND2X0 U36 ( .IN1(n32), .IN2(n31), .QN(out1[3]) );
  NAND2X0 U37 ( .IN1(n36), .IN2(n35), .QN(out1[4]) );
  NAND2X0 U38 ( .IN1(n23), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U39 ( .IN1(in1[2]), .IN2(n22), .QN(n23) );
  INVX0 U40 ( .INP(in1[2]), .ZN(n111) );
  NOR2X0 U41 ( .IN1(n28), .IN2(n26), .QN(n3) );
  NOR2X0 U42 ( .IN1(n142), .IN2(n21), .QN(n1) );
  INVX0 U43 ( .INP(n132), .ZN(n141) );
  INVX0 U44 ( .INP(n130), .ZN(n137) );
  NOR2X0 U45 ( .IN1(n142), .IN2(n111), .QN(n138) );
  MUX21X1 U46 ( .IN1(n22), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  NAND3X0 U47 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  NOR3X0 U48 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  INVX0 U49 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U50 ( .INP(in2[2]), .ZN(n6) );
  INVX0 U51 ( .INP(in2[4]), .ZN(n7) );
  INVX0 U52 ( .INP(in2[6]), .ZN(n8) );
  INVX0 U53 ( .INP(in2[8]), .ZN(n9) );
  INVX0 U54 ( .INP(in2[10]), .ZN(n10) );
  INVX0 U55 ( .INP(in2[12]), .ZN(n11) );
  INVX0 U56 ( .INP(in2[13]), .ZN(n12) );
  INVX0 U57 ( .INP(in2[14]), .ZN(n13) );
  INVX0 U58 ( .INP(in2[15]), .ZN(n14) );
  INVX0 U59 ( .INP(in2[16]), .ZN(n15) );
  INVX0 U60 ( .INP(in2[17]), .ZN(n16) );
  INVX0 U61 ( .INP(in2[18]), .ZN(n17) );
  INVX0 U62 ( .INP(in2[19]), .ZN(n18) );
  INVX0 U63 ( .INP(in2[20]), .ZN(n19) );
  INVX0 U64 ( .INP(in2[21]), .ZN(n20) );
  INVX0 U65 ( .INP(in2[22]), .ZN(n21) );
  INVX0 U66 ( .INP(in1[1]), .ZN(n22) );
  INVX0 U67 ( .INP(n138), .ZN(n140) );
  NOR2X0 U68 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n25) );
  AOI21X1 U69 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n25), .QN(n27) );
  NOR2X0 U70 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U71 ( .IN1(n24), .IN2(in2[0]), .IN3(n138), .IN4(n27), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U72 ( .INP(n133), .ZN(n67) );
  NOR2X0 U73 ( .IN1(n67), .IN2(n6), .QN(n28) );
  OA21X1 U74 ( .IN1(n25), .IN2(n6), .IN3(n30), .Q(n29) );
  AO22X1 U75 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n29), .Q(n26) );
  AOI22X1 U76 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n29), .QN(n32) );
  NOR2X0 U77 ( .IN1(in2[3]), .IN2(n30), .QN(n33) );
  AO21X1 U78 ( .IN1(in2[3]), .IN2(n30), .IN3(n33), .Q(n34) );
  OA22X1 U79 ( .IN1(n6), .IN2(n130), .IN3(n140), .IN4(n34), .Q(n31) );
  OA21X1 U80 ( .IN1(n33), .IN2(n7), .IN3(n37), .Q(n38) );
  AOI22X1 U81 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n38), .QN(n36) );
  OA22X1 U82 ( .IN1(n67), .IN2(n7), .IN3(n141), .IN4(n34), .Q(n35) );
  NOR2X0 U83 ( .IN1(in2[5]), .IN2(n37), .QN(n41) );
  AO21X1 U84 ( .IN1(in2[5]), .IN2(n37), .IN3(n41), .Q(n42) );
  OA22X1 U85 ( .IN1(n7), .IN2(n130), .IN3(n140), .IN4(n42), .Q(n40) );
  AOI22X1 U86 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n38), .QN(n39) );
  OA21X1 U87 ( .IN1(n41), .IN2(n8), .IN3(n45), .Q(n46) );
  AOI22X1 U88 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n46), .QN(n44) );
  OA22X1 U89 ( .IN1(n67), .IN2(n8), .IN3(n141), .IN4(n42), .Q(n43) );
  NOR2X0 U90 ( .IN1(in2[7]), .IN2(n45), .QN(n49) );
  AO21X1 U91 ( .IN1(in2[7]), .IN2(n45), .IN3(n49), .Q(n50) );
  OA22X1 U92 ( .IN1(n8), .IN2(n130), .IN3(n140), .IN4(n50), .Q(n48) );
  AOI22X1 U93 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n46), .QN(n47) );
  OA21X1 U94 ( .IN1(n49), .IN2(n9), .IN3(n53), .Q(n54) );
  AOI22X1 U95 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n54), .QN(n52) );
  OA22X1 U96 ( .IN1(n67), .IN2(n9), .IN3(n141), .IN4(n50), .Q(n51) );
  NOR2X0 U97 ( .IN1(in2[9]), .IN2(n53), .QN(n57) );
  AO21X1 U98 ( .IN1(in2[9]), .IN2(n53), .IN3(n57), .Q(n58) );
  OA22X1 U99 ( .IN1(n9), .IN2(n130), .IN3(n140), .IN4(n58), .Q(n56) );
  AOI22X1 U100 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n54), .QN(n55) );
  OA21X1 U101 ( .IN1(n57), .IN2(n10), .IN3(n61), .Q(n62) );
  AOI22X1 U102 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n62), .QN(n60) );
  OA22X1 U103 ( .IN1(n67), .IN2(n10), .IN3(n141), .IN4(n58), .Q(n59) );
  NOR2X0 U104 ( .IN1(in2[11]), .IN2(n61), .QN(n65) );
  AO21X1 U105 ( .IN1(in2[11]), .IN2(n61), .IN3(n65), .Q(n66) );
  OA22X1 U106 ( .IN1(n10), .IN2(n130), .IN3(n140), .IN4(n66), .Q(n64) );
  AOI22X1 U107 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n62), .QN(n63) );
  OA21X1 U108 ( .IN1(n65), .IN2(n11), .IN3(n77), .Q(n70) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n70), .QN(n69) );
  OA22X1 U110 ( .IN1(n67), .IN2(n11), .IN3(n141), .IN4(n66), .Q(n68) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n12), .S(n71), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n11), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n13), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n12), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n12), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n14), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n13), .IN4(n85), .IN5(n84), 
        .Q(out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n15), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n14), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n14), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n16), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n15), .IN4(n97), .IN5(n96), 
        .Q(out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n17), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n16), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n16), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n18), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n17), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n19), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n18), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n18), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n20), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n19), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n21), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n20), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n20), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n21), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_45 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n49), .IN2(n9), .QN(n53) );
  NAND2X0 U4 ( .IN1(n57), .IN2(n10), .QN(n61) );
  NAND2X0 U5 ( .IN1(n25), .IN2(n6), .QN(n30) );
  NAND2X0 U6 ( .IN1(n41), .IN2(n8), .QN(n45) );
  NAND2X0 U7 ( .IN1(n33), .IN2(n7), .QN(n37) );
  NAND2X0 U8 ( .IN1(n65), .IN2(n11), .QN(n77) );
  NAND2X0 U9 ( .IN1(n81), .IN2(n13), .QN(n89) );
  NAND2X0 U10 ( .IN1(n93), .IN2(n15), .QN(n101) );
  NAND2X0 U11 ( .IN1(n105), .IN2(n17), .QN(n114) );
  NAND2X0 U12 ( .IN1(in1[2]), .IN2(n77), .QN(n71) );
  NAND2X0 U13 ( .IN1(n70), .IN2(n132), .QN(n74) );
  NAND2X0 U14 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U15 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U16 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U17 ( .IN1(n118), .IN2(n19), .QN(n125) );
  NAND2X0 U18 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U19 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U20 ( .IN1(n27), .IN2(n132), .QN(n4) );
  NAND2X0 U21 ( .IN1(n48), .IN2(n47), .QN(out1[7]) );
  NAND2X0 U22 ( .IN1(n52), .IN2(n51), .QN(out1[8]) );
  NAND2X0 U23 ( .IN1(n56), .IN2(n55), .QN(out1[9]) );
  NAND2X0 U24 ( .IN1(n60), .IN2(n59), .QN(out1[10]) );
  NAND2X0 U25 ( .IN1(n64), .IN2(n63), .QN(out1[11]) );
  NAND2X0 U26 ( .IN1(n69), .IN2(n68), .QN(out1[12]) );
  NAND2X0 U27 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U28 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U29 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U30 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U31 ( .IN1(n141), .IN2(n130), .QN(n24) );
  NAND2X0 U32 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NAND2X0 U33 ( .IN1(n36), .IN2(n35), .QN(out1[4]) );
  NAND2X0 U34 ( .IN1(n32), .IN2(n31), .QN(out1[3]) );
  NAND2X0 U35 ( .IN1(n40), .IN2(n39), .QN(out1[5]) );
  NAND2X0 U36 ( .IN1(n44), .IN2(n43), .QN(out1[6]) );
  NAND2X0 U37 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U38 ( .IN1(n23), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U39 ( .IN1(in1[2]), .IN2(n22), .QN(n23) );
  NOR2X0 U40 ( .IN1(n28), .IN2(n26), .QN(n3) );
  INVX0 U41 ( .INP(n130), .ZN(n137) );
  NAND3X0 U42 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  NOR2X0 U43 ( .IN1(n142), .IN2(n21), .QN(n1) );
  NOR2X0 U44 ( .IN1(n142), .IN2(n111), .QN(n138) );
  MUX21X1 U45 ( .IN1(n22), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  INVX0 U46 ( .INP(n132), .ZN(n141) );
  NOR3X0 U47 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  INVX0 U48 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U49 ( .INP(in2[2]), .ZN(n6) );
  INVX0 U50 ( .INP(in2[4]), .ZN(n7) );
  INVX0 U51 ( .INP(in2[6]), .ZN(n8) );
  INVX0 U52 ( .INP(in2[8]), .ZN(n9) );
  INVX0 U53 ( .INP(in2[10]), .ZN(n10) );
  INVX0 U54 ( .INP(in2[12]), .ZN(n11) );
  INVX0 U55 ( .INP(in2[13]), .ZN(n12) );
  INVX0 U56 ( .INP(in2[14]), .ZN(n13) );
  INVX0 U57 ( .INP(in2[15]), .ZN(n14) );
  INVX0 U58 ( .INP(in2[16]), .ZN(n15) );
  INVX0 U59 ( .INP(in2[17]), .ZN(n16) );
  INVX0 U60 ( .INP(in2[18]), .ZN(n17) );
  INVX0 U61 ( .INP(in2[19]), .ZN(n18) );
  INVX0 U62 ( .INP(in2[20]), .ZN(n19) );
  INVX0 U63 ( .INP(in2[21]), .ZN(n20) );
  INVX0 U64 ( .INP(in2[22]), .ZN(n21) );
  INVX0 U65 ( .INP(in1[1]), .ZN(n22) );
  INVX0 U66 ( .INP(in1[2]), .ZN(n111) );
  INVX0 U67 ( .INP(n138), .ZN(n140) );
  NOR2X0 U68 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n25) );
  AOI21X1 U69 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n25), .QN(n27) );
  NOR2X0 U70 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U71 ( .IN1(n24), .IN2(in2[0]), .IN3(n138), .IN4(n27), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U72 ( .INP(n133), .ZN(n67) );
  NOR2X0 U73 ( .IN1(n67), .IN2(n6), .QN(n28) );
  OA21X1 U74 ( .IN1(n25), .IN2(n6), .IN3(n30), .Q(n29) );
  AO22X1 U75 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n29), .Q(n26) );
  AOI22X1 U76 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n29), .QN(n32) );
  NOR2X0 U77 ( .IN1(in2[3]), .IN2(n30), .QN(n33) );
  AO21X1 U78 ( .IN1(in2[3]), .IN2(n30), .IN3(n33), .Q(n34) );
  OA22X1 U79 ( .IN1(n6), .IN2(n130), .IN3(n140), .IN4(n34), .Q(n31) );
  OA21X1 U80 ( .IN1(n33), .IN2(n7), .IN3(n37), .Q(n38) );
  AOI22X1 U81 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n38), .QN(n36) );
  OA22X1 U82 ( .IN1(n67), .IN2(n7), .IN3(n141), .IN4(n34), .Q(n35) );
  NOR2X0 U83 ( .IN1(in2[5]), .IN2(n37), .QN(n41) );
  AO21X1 U84 ( .IN1(in2[5]), .IN2(n37), .IN3(n41), .Q(n42) );
  OA22X1 U85 ( .IN1(n7), .IN2(n130), .IN3(n140), .IN4(n42), .Q(n40) );
  AOI22X1 U86 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n38), .QN(n39) );
  OA21X1 U87 ( .IN1(n41), .IN2(n8), .IN3(n45), .Q(n46) );
  AOI22X1 U88 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n46), .QN(n44) );
  OA22X1 U89 ( .IN1(n67), .IN2(n8), .IN3(n141), .IN4(n42), .Q(n43) );
  NOR2X0 U90 ( .IN1(in2[7]), .IN2(n45), .QN(n49) );
  AO21X1 U91 ( .IN1(in2[7]), .IN2(n45), .IN3(n49), .Q(n50) );
  OA22X1 U92 ( .IN1(n8), .IN2(n130), .IN3(n140), .IN4(n50), .Q(n48) );
  AOI22X1 U93 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n46), .QN(n47) );
  OA21X1 U94 ( .IN1(n49), .IN2(n9), .IN3(n53), .Q(n54) );
  AOI22X1 U95 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n54), .QN(n52) );
  OA22X1 U96 ( .IN1(n67), .IN2(n9), .IN3(n141), .IN4(n50), .Q(n51) );
  NOR2X0 U97 ( .IN1(in2[9]), .IN2(n53), .QN(n57) );
  AO21X1 U98 ( .IN1(in2[9]), .IN2(n53), .IN3(n57), .Q(n58) );
  OA22X1 U99 ( .IN1(n9), .IN2(n130), .IN3(n140), .IN4(n58), .Q(n56) );
  AOI22X1 U100 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n54), .QN(n55) );
  OA21X1 U101 ( .IN1(n57), .IN2(n10), .IN3(n61), .Q(n62) );
  AOI22X1 U102 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n62), .QN(n60) );
  OA22X1 U103 ( .IN1(n67), .IN2(n10), .IN3(n141), .IN4(n58), .Q(n59) );
  NOR2X0 U104 ( .IN1(in2[11]), .IN2(n61), .QN(n65) );
  AO21X1 U105 ( .IN1(in2[11]), .IN2(n61), .IN3(n65), .Q(n66) );
  OA22X1 U106 ( .IN1(n10), .IN2(n130), .IN3(n140), .IN4(n66), .Q(n64) );
  AOI22X1 U107 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n62), .QN(n63) );
  OA21X1 U108 ( .IN1(n65), .IN2(n11), .IN3(n77), .Q(n70) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n70), .QN(n69) );
  OA22X1 U110 ( .IN1(n67), .IN2(n11), .IN3(n141), .IN4(n66), .Q(n68) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n12), .S(n71), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n11), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n13), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n12), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n12), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n14), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n13), .IN4(n85), .IN5(n84), 
        .Q(out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n15), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n14), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n14), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n16), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n15), .IN4(n97), .IN5(n96), 
        .Q(out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n17), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n16), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n16), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n18), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n17), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n19), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n18), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n18), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n20), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n19), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n21), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n20), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n20), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n21), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_46 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n57), .IN2(n10), .QN(n61) );
  NAND2X0 U4 ( .IN1(n33), .IN2(n7), .QN(n37) );
  NAND2X0 U5 ( .IN1(n49), .IN2(n9), .QN(n53) );
  NAND2X0 U6 ( .IN1(n41), .IN2(n8), .QN(n45) );
  NAND2X0 U7 ( .IN1(n65), .IN2(n11), .QN(n77) );
  NAND2X0 U8 ( .IN1(n81), .IN2(n13), .QN(n89) );
  NAND2X0 U9 ( .IN1(n93), .IN2(n15), .QN(n101) );
  NAND2X0 U10 ( .IN1(n105), .IN2(n17), .QN(n114) );
  NAND2X0 U11 ( .IN1(n118), .IN2(n19), .QN(n125) );
  NAND2X0 U12 ( .IN1(n25), .IN2(n6), .QN(n30) );
  NAND2X0 U13 ( .IN1(in1[2]), .IN2(n77), .QN(n71) );
  NAND2X0 U14 ( .IN1(n70), .IN2(n132), .QN(n74) );
  NAND2X0 U15 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U16 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U17 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U18 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U19 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U20 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U21 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U22 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U23 ( .IN1(n56), .IN2(n55), .QN(out1[9]) );
  NAND2X0 U24 ( .IN1(n60), .IN2(n59), .QN(out1[10]) );
  NAND2X0 U25 ( .IN1(n64), .IN2(n63), .QN(out1[11]) );
  NAND2X0 U26 ( .IN1(n69), .IN2(n68), .QN(out1[12]) );
  NAND2X0 U27 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U28 ( .IN1(n23), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U29 ( .IN1(in1[2]), .IN2(n22), .QN(n23) );
  NAND2X0 U30 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NAND2X0 U31 ( .IN1(n27), .IN2(n132), .QN(n4) );
  NAND2X0 U32 ( .IN1(n32), .IN2(n31), .QN(out1[3]) );
  NAND2X0 U33 ( .IN1(n36), .IN2(n35), .QN(out1[4]) );
  NAND2X0 U34 ( .IN1(n44), .IN2(n43), .QN(out1[6]) );
  NAND2X0 U35 ( .IN1(n40), .IN2(n39), .QN(out1[5]) );
  NAND2X0 U36 ( .IN1(n48), .IN2(n47), .QN(out1[7]) );
  NAND2X0 U37 ( .IN1(n52), .IN2(n51), .QN(out1[8]) );
  NAND2X0 U38 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U39 ( .IN1(n141), .IN2(n130), .QN(n24) );
  NOR2X0 U40 ( .IN1(n28), .IN2(n26), .QN(n3) );
  NOR2X0 U41 ( .IN1(n142), .IN2(n21), .QN(n1) );
  INVX0 U42 ( .INP(n132), .ZN(n141) );
  INVX0 U43 ( .INP(n130), .ZN(n137) );
  NAND3X0 U44 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  NOR3X0 U45 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  NOR2X0 U46 ( .IN1(n142), .IN2(n111), .QN(n138) );
  MUX21X1 U47 ( .IN1(n22), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  INVX0 U48 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U49 ( .INP(in2[2]), .ZN(n6) );
  INVX0 U50 ( .INP(in2[4]), .ZN(n7) );
  INVX0 U51 ( .INP(in2[6]), .ZN(n8) );
  INVX0 U52 ( .INP(in2[8]), .ZN(n9) );
  INVX0 U53 ( .INP(in2[10]), .ZN(n10) );
  INVX0 U54 ( .INP(in2[12]), .ZN(n11) );
  INVX0 U55 ( .INP(in2[13]), .ZN(n12) );
  INVX0 U56 ( .INP(in2[14]), .ZN(n13) );
  INVX0 U57 ( .INP(in2[15]), .ZN(n14) );
  INVX0 U58 ( .INP(in2[16]), .ZN(n15) );
  INVX0 U59 ( .INP(in2[17]), .ZN(n16) );
  INVX0 U60 ( .INP(in2[18]), .ZN(n17) );
  INVX0 U61 ( .INP(in2[19]), .ZN(n18) );
  INVX0 U62 ( .INP(in2[20]), .ZN(n19) );
  INVX0 U63 ( .INP(in2[21]), .ZN(n20) );
  INVX0 U64 ( .INP(in2[22]), .ZN(n21) );
  INVX0 U65 ( .INP(in1[1]), .ZN(n22) );
  INVX0 U66 ( .INP(in1[2]), .ZN(n111) );
  INVX0 U67 ( .INP(n138), .ZN(n140) );
  NOR2X0 U68 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n25) );
  AOI21X1 U69 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n25), .QN(n27) );
  NOR2X0 U70 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U71 ( .IN1(n24), .IN2(in2[0]), .IN3(n138), .IN4(n27), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U72 ( .INP(n133), .ZN(n67) );
  NOR2X0 U73 ( .IN1(n67), .IN2(n6), .QN(n28) );
  OA21X1 U74 ( .IN1(n25), .IN2(n6), .IN3(n30), .Q(n29) );
  AO22X1 U75 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n29), .Q(n26) );
  AOI22X1 U76 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n29), .QN(n32) );
  NOR2X0 U77 ( .IN1(in2[3]), .IN2(n30), .QN(n33) );
  AO21X1 U78 ( .IN1(in2[3]), .IN2(n30), .IN3(n33), .Q(n34) );
  OA22X1 U79 ( .IN1(n6), .IN2(n130), .IN3(n140), .IN4(n34), .Q(n31) );
  OA21X1 U80 ( .IN1(n33), .IN2(n7), .IN3(n37), .Q(n38) );
  AOI22X1 U81 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n38), .QN(n36) );
  OA22X1 U82 ( .IN1(n67), .IN2(n7), .IN3(n141), .IN4(n34), .Q(n35) );
  NOR2X0 U83 ( .IN1(in2[5]), .IN2(n37), .QN(n41) );
  AO21X1 U84 ( .IN1(in2[5]), .IN2(n37), .IN3(n41), .Q(n42) );
  OA22X1 U85 ( .IN1(n7), .IN2(n130), .IN3(n140), .IN4(n42), .Q(n40) );
  AOI22X1 U86 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n38), .QN(n39) );
  OA21X1 U87 ( .IN1(n41), .IN2(n8), .IN3(n45), .Q(n46) );
  AOI22X1 U88 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n46), .QN(n44) );
  OA22X1 U89 ( .IN1(n67), .IN2(n8), .IN3(n141), .IN4(n42), .Q(n43) );
  NOR2X0 U90 ( .IN1(in2[7]), .IN2(n45), .QN(n49) );
  AO21X1 U91 ( .IN1(in2[7]), .IN2(n45), .IN3(n49), .Q(n50) );
  OA22X1 U92 ( .IN1(n8), .IN2(n130), .IN3(n140), .IN4(n50), .Q(n48) );
  AOI22X1 U93 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n46), .QN(n47) );
  OA21X1 U94 ( .IN1(n49), .IN2(n9), .IN3(n53), .Q(n54) );
  AOI22X1 U95 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n54), .QN(n52) );
  OA22X1 U96 ( .IN1(n67), .IN2(n9), .IN3(n141), .IN4(n50), .Q(n51) );
  NOR2X0 U97 ( .IN1(in2[9]), .IN2(n53), .QN(n57) );
  AO21X1 U98 ( .IN1(in2[9]), .IN2(n53), .IN3(n57), .Q(n58) );
  OA22X1 U99 ( .IN1(n9), .IN2(n130), .IN3(n140), .IN4(n58), .Q(n56) );
  AOI22X1 U100 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n54), .QN(n55) );
  OA21X1 U101 ( .IN1(n57), .IN2(n10), .IN3(n61), .Q(n62) );
  AOI22X1 U102 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n62), .QN(n60) );
  OA22X1 U103 ( .IN1(n67), .IN2(n10), .IN3(n141), .IN4(n58), .Q(n59) );
  NOR2X0 U104 ( .IN1(in2[11]), .IN2(n61), .QN(n65) );
  AO21X1 U105 ( .IN1(in2[11]), .IN2(n61), .IN3(n65), .Q(n66) );
  OA22X1 U106 ( .IN1(n10), .IN2(n130), .IN3(n140), .IN4(n66), .Q(n64) );
  AOI22X1 U107 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n62), .QN(n63) );
  OA21X1 U108 ( .IN1(n65), .IN2(n11), .IN3(n77), .Q(n70) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n70), .QN(n69) );
  OA22X1 U110 ( .IN1(n67), .IN2(n11), .IN3(n141), .IN4(n66), .Q(n68) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n12), .S(n71), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n11), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n13), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n12), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n12), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n14), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n13), .IN4(n85), .IN5(n84), 
        .Q(out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n15), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n14), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n14), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n16), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n15), .IN4(n97), .IN5(n96), 
        .Q(out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n17), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n16), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n16), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n18), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n17), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n19), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n18), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n18), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n20), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n19), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n21), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n20), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n20), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n21), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_47 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n57), .IN2(n10), .QN(n61) );
  NAND2X0 U4 ( .IN1(n25), .IN2(n6), .QN(n30) );
  NAND2X0 U5 ( .IN1(n33), .IN2(n7), .QN(n37) );
  NAND2X0 U6 ( .IN1(n49), .IN2(n9), .QN(n53) );
  NAND2X0 U7 ( .IN1(n41), .IN2(n8), .QN(n45) );
  NAND2X0 U8 ( .IN1(n65), .IN2(n11), .QN(n77) );
  NAND2X0 U9 ( .IN1(n81), .IN2(n13), .QN(n89) );
  NAND2X0 U10 ( .IN1(n93), .IN2(n15), .QN(n101) );
  NAND2X0 U11 ( .IN1(n105), .IN2(n17), .QN(n114) );
  NAND2X0 U12 ( .IN1(in1[2]), .IN2(n77), .QN(n71) );
  NAND2X0 U13 ( .IN1(n70), .IN2(n132), .QN(n74) );
  NAND2X0 U14 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U15 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U16 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U17 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U18 ( .IN1(n118), .IN2(n19), .QN(n125) );
  NAND2X0 U19 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U20 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U21 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U22 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U23 ( .IN1(n141), .IN2(n130), .QN(n24) );
  NAND2X0 U24 ( .IN1(n27), .IN2(n132), .QN(n4) );
  NAND2X0 U25 ( .IN1(n56), .IN2(n55), .QN(out1[9]) );
  NAND2X0 U26 ( .IN1(n60), .IN2(n59), .QN(out1[10]) );
  NAND2X0 U27 ( .IN1(n64), .IN2(n63), .QN(out1[11]) );
  NAND2X0 U28 ( .IN1(n69), .IN2(n68), .QN(out1[12]) );
  NAND2X0 U29 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U30 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U31 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NAND2X0 U32 ( .IN1(n32), .IN2(n31), .QN(out1[3]) );
  NAND2X0 U33 ( .IN1(n36), .IN2(n35), .QN(out1[4]) );
  NAND2X0 U34 ( .IN1(n40), .IN2(n39), .QN(out1[5]) );
  NAND2X0 U35 ( .IN1(n44), .IN2(n43), .QN(out1[6]) );
  NAND2X0 U36 ( .IN1(n48), .IN2(n47), .QN(out1[7]) );
  NAND2X0 U37 ( .IN1(n52), .IN2(n51), .QN(out1[8]) );
  NAND2X0 U38 ( .IN1(n23), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U39 ( .IN1(in1[2]), .IN2(n22), .QN(n23) );
  NOR2X0 U40 ( .IN1(n28), .IN2(n26), .QN(n3) );
  INVX0 U41 ( .INP(n130), .ZN(n137) );
  NAND3X0 U42 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  NOR2X0 U43 ( .IN1(n142), .IN2(n21), .QN(n1) );
  INVX0 U44 ( .INP(n132), .ZN(n141) );
  NOR3X0 U45 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  NOR2X0 U46 ( .IN1(n142), .IN2(n111), .QN(n138) );
  MUX21X1 U47 ( .IN1(n22), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  INVX0 U48 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U49 ( .INP(in2[2]), .ZN(n6) );
  INVX0 U50 ( .INP(in2[4]), .ZN(n7) );
  INVX0 U51 ( .INP(in2[6]), .ZN(n8) );
  INVX0 U52 ( .INP(in2[8]), .ZN(n9) );
  INVX0 U53 ( .INP(in2[10]), .ZN(n10) );
  INVX0 U54 ( .INP(in2[12]), .ZN(n11) );
  INVX0 U55 ( .INP(in2[13]), .ZN(n12) );
  INVX0 U56 ( .INP(in2[14]), .ZN(n13) );
  INVX0 U57 ( .INP(in2[15]), .ZN(n14) );
  INVX0 U58 ( .INP(in2[16]), .ZN(n15) );
  INVX0 U59 ( .INP(in2[17]), .ZN(n16) );
  INVX0 U60 ( .INP(in2[18]), .ZN(n17) );
  INVX0 U61 ( .INP(in2[19]), .ZN(n18) );
  INVX0 U62 ( .INP(in2[20]), .ZN(n19) );
  INVX0 U63 ( .INP(in2[21]), .ZN(n20) );
  INVX0 U64 ( .INP(in2[22]), .ZN(n21) );
  INVX0 U65 ( .INP(in1[1]), .ZN(n22) );
  INVX0 U66 ( .INP(in1[2]), .ZN(n111) );
  INVX0 U67 ( .INP(n138), .ZN(n140) );
  NOR2X0 U68 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n25) );
  AOI21X1 U69 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n25), .QN(n27) );
  NOR2X0 U70 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U71 ( .IN1(n24), .IN2(in2[0]), .IN3(n138), .IN4(n27), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U72 ( .INP(n133), .ZN(n67) );
  NOR2X0 U73 ( .IN1(n67), .IN2(n6), .QN(n28) );
  OA21X1 U74 ( .IN1(n25), .IN2(n6), .IN3(n30), .Q(n29) );
  AO22X1 U75 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n29), .Q(n26) );
  AOI22X1 U76 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n29), .QN(n32) );
  NOR2X0 U77 ( .IN1(in2[3]), .IN2(n30), .QN(n33) );
  AO21X1 U78 ( .IN1(in2[3]), .IN2(n30), .IN3(n33), .Q(n34) );
  OA22X1 U79 ( .IN1(n6), .IN2(n130), .IN3(n140), .IN4(n34), .Q(n31) );
  OA21X1 U80 ( .IN1(n33), .IN2(n7), .IN3(n37), .Q(n38) );
  AOI22X1 U81 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n38), .QN(n36) );
  OA22X1 U82 ( .IN1(n67), .IN2(n7), .IN3(n141), .IN4(n34), .Q(n35) );
  NOR2X0 U83 ( .IN1(in2[5]), .IN2(n37), .QN(n41) );
  AO21X1 U84 ( .IN1(in2[5]), .IN2(n37), .IN3(n41), .Q(n42) );
  OA22X1 U85 ( .IN1(n7), .IN2(n130), .IN3(n140), .IN4(n42), .Q(n40) );
  AOI22X1 U86 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n38), .QN(n39) );
  OA21X1 U87 ( .IN1(n41), .IN2(n8), .IN3(n45), .Q(n46) );
  AOI22X1 U88 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n46), .QN(n44) );
  OA22X1 U89 ( .IN1(n67), .IN2(n8), .IN3(n141), .IN4(n42), .Q(n43) );
  NOR2X0 U90 ( .IN1(in2[7]), .IN2(n45), .QN(n49) );
  AO21X1 U91 ( .IN1(in2[7]), .IN2(n45), .IN3(n49), .Q(n50) );
  OA22X1 U92 ( .IN1(n8), .IN2(n130), .IN3(n140), .IN4(n50), .Q(n48) );
  AOI22X1 U93 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n46), .QN(n47) );
  OA21X1 U94 ( .IN1(n49), .IN2(n9), .IN3(n53), .Q(n54) );
  AOI22X1 U95 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n54), .QN(n52) );
  OA22X1 U96 ( .IN1(n67), .IN2(n9), .IN3(n141), .IN4(n50), .Q(n51) );
  NOR2X0 U97 ( .IN1(in2[9]), .IN2(n53), .QN(n57) );
  AO21X1 U98 ( .IN1(in2[9]), .IN2(n53), .IN3(n57), .Q(n58) );
  OA22X1 U99 ( .IN1(n9), .IN2(n130), .IN3(n140), .IN4(n58), .Q(n56) );
  AOI22X1 U100 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n54), .QN(n55) );
  OA21X1 U101 ( .IN1(n57), .IN2(n10), .IN3(n61), .Q(n62) );
  AOI22X1 U102 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n62), .QN(n60) );
  OA22X1 U103 ( .IN1(n67), .IN2(n10), .IN3(n141), .IN4(n58), .Q(n59) );
  NOR2X0 U104 ( .IN1(in2[11]), .IN2(n61), .QN(n65) );
  AO21X1 U105 ( .IN1(in2[11]), .IN2(n61), .IN3(n65), .Q(n66) );
  OA22X1 U106 ( .IN1(n10), .IN2(n130), .IN3(n140), .IN4(n66), .Q(n64) );
  AOI22X1 U107 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n62), .QN(n63) );
  OA21X1 U108 ( .IN1(n65), .IN2(n11), .IN3(n77), .Q(n70) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n70), .QN(n69) );
  OA22X1 U110 ( .IN1(n67), .IN2(n11), .IN3(n141), .IN4(n66), .Q(n68) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n12), .S(n71), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n11), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n13), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n12), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n12), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n14), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n13), .IN4(n85), .IN5(n84), 
        .Q(out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n15), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n14), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n14), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n16), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n15), .IN4(n97), .IN5(n96), 
        .Q(out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n17), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n16), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n16), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n18), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n17), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n19), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n18), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n18), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n20), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n19), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n21), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n20), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n20), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n21), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_48 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n25), .IN2(n6), .QN(n30) );
  NAND2X0 U4 ( .IN1(n33), .IN2(n7), .QN(n37) );
  NAND2X0 U5 ( .IN1(n41), .IN2(n8), .QN(n45) );
  NAND2X0 U6 ( .IN1(n57), .IN2(n10), .QN(n61) );
  NAND2X0 U7 ( .IN1(n49), .IN2(n9), .QN(n53) );
  NAND2X0 U8 ( .IN1(n65), .IN2(n11), .QN(n77) );
  NAND2X0 U9 ( .IN1(n81), .IN2(n13), .QN(n89) );
  NAND2X0 U10 ( .IN1(n93), .IN2(n15), .QN(n101) );
  NAND2X0 U11 ( .IN1(n105), .IN2(n17), .QN(n114) );
  NAND2X0 U12 ( .IN1(n118), .IN2(n19), .QN(n125) );
  NAND2X0 U13 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U14 ( .IN1(in1[2]), .IN2(n77), .QN(n71) );
  NAND2X0 U15 ( .IN1(n70), .IN2(n132), .QN(n74) );
  NAND2X0 U16 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U17 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U18 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U19 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U20 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U21 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U22 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U23 ( .IN1(n141), .IN2(n130), .QN(n24) );
  NAND2X0 U24 ( .IN1(n27), .IN2(n132), .QN(n4) );
  NAND2X0 U25 ( .IN1(n64), .IN2(n63), .QN(out1[11]) );
  NAND2X0 U26 ( .IN1(n69), .IN2(n68), .QN(out1[12]) );
  NAND2X0 U27 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U28 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U29 ( .IN1(n23), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U30 ( .IN1(in1[2]), .IN2(n22), .QN(n23) );
  NAND2X0 U31 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NAND2X0 U32 ( .IN1(n32), .IN2(n31), .QN(out1[3]) );
  NAND2X0 U33 ( .IN1(n36), .IN2(n35), .QN(out1[4]) );
  NAND2X0 U34 ( .IN1(n40), .IN2(n39), .QN(out1[5]) );
  NAND2X0 U35 ( .IN1(n44), .IN2(n43), .QN(out1[6]) );
  NAND2X0 U36 ( .IN1(n48), .IN2(n47), .QN(out1[7]) );
  NAND2X0 U37 ( .IN1(n52), .IN2(n51), .QN(out1[8]) );
  NAND2X0 U38 ( .IN1(n56), .IN2(n55), .QN(out1[9]) );
  NAND2X0 U39 ( .IN1(n60), .IN2(n59), .QN(out1[10]) );
  NOR2X0 U40 ( .IN1(n28), .IN2(n26), .QN(n3) );
  NOR2X0 U41 ( .IN1(n142), .IN2(n21), .QN(n1) );
  INVX0 U42 ( .INP(n132), .ZN(n141) );
  INVX0 U43 ( .INP(n130), .ZN(n137) );
  NAND3X0 U44 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  NOR3X0 U45 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  NOR2X0 U46 ( .IN1(n142), .IN2(n111), .QN(n138) );
  MUX21X1 U47 ( .IN1(n22), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  INVX0 U48 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U49 ( .INP(in2[2]), .ZN(n6) );
  INVX0 U50 ( .INP(in2[4]), .ZN(n7) );
  INVX0 U51 ( .INP(in2[6]), .ZN(n8) );
  INVX0 U52 ( .INP(in2[8]), .ZN(n9) );
  INVX0 U53 ( .INP(in2[10]), .ZN(n10) );
  INVX0 U54 ( .INP(in2[12]), .ZN(n11) );
  INVX0 U55 ( .INP(in2[13]), .ZN(n12) );
  INVX0 U56 ( .INP(in2[14]), .ZN(n13) );
  INVX0 U57 ( .INP(in2[15]), .ZN(n14) );
  INVX0 U58 ( .INP(in2[16]), .ZN(n15) );
  INVX0 U59 ( .INP(in2[17]), .ZN(n16) );
  INVX0 U60 ( .INP(in2[18]), .ZN(n17) );
  INVX0 U61 ( .INP(in2[19]), .ZN(n18) );
  INVX0 U62 ( .INP(in2[20]), .ZN(n19) );
  INVX0 U63 ( .INP(in2[21]), .ZN(n20) );
  INVX0 U64 ( .INP(in2[22]), .ZN(n21) );
  INVX0 U65 ( .INP(in1[1]), .ZN(n22) );
  INVX0 U66 ( .INP(in1[2]), .ZN(n111) );
  INVX0 U67 ( .INP(n138), .ZN(n140) );
  NOR2X0 U68 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n25) );
  AOI21X1 U69 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n25), .QN(n27) );
  NOR2X0 U70 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U71 ( .IN1(n24), .IN2(in2[0]), .IN3(n138), .IN4(n27), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U72 ( .INP(n133), .ZN(n67) );
  NOR2X0 U73 ( .IN1(n67), .IN2(n6), .QN(n28) );
  OA21X1 U74 ( .IN1(n25), .IN2(n6), .IN3(n30), .Q(n29) );
  AO22X1 U75 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n29), .Q(n26) );
  AOI22X1 U76 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n29), .QN(n32) );
  NOR2X0 U77 ( .IN1(in2[3]), .IN2(n30), .QN(n33) );
  AO21X1 U78 ( .IN1(in2[3]), .IN2(n30), .IN3(n33), .Q(n34) );
  OA22X1 U79 ( .IN1(n6), .IN2(n130), .IN3(n140), .IN4(n34), .Q(n31) );
  OA21X1 U80 ( .IN1(n33), .IN2(n7), .IN3(n37), .Q(n38) );
  AOI22X1 U81 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n38), .QN(n36) );
  OA22X1 U82 ( .IN1(n67), .IN2(n7), .IN3(n141), .IN4(n34), .Q(n35) );
  NOR2X0 U83 ( .IN1(in2[5]), .IN2(n37), .QN(n41) );
  AO21X1 U84 ( .IN1(in2[5]), .IN2(n37), .IN3(n41), .Q(n42) );
  OA22X1 U85 ( .IN1(n7), .IN2(n130), .IN3(n140), .IN4(n42), .Q(n40) );
  AOI22X1 U86 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n38), .QN(n39) );
  OA21X1 U87 ( .IN1(n41), .IN2(n8), .IN3(n45), .Q(n46) );
  AOI22X1 U88 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n46), .QN(n44) );
  OA22X1 U89 ( .IN1(n67), .IN2(n8), .IN3(n141), .IN4(n42), .Q(n43) );
  NOR2X0 U90 ( .IN1(in2[7]), .IN2(n45), .QN(n49) );
  AO21X1 U91 ( .IN1(in2[7]), .IN2(n45), .IN3(n49), .Q(n50) );
  OA22X1 U92 ( .IN1(n8), .IN2(n130), .IN3(n140), .IN4(n50), .Q(n48) );
  AOI22X1 U93 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n46), .QN(n47) );
  OA21X1 U94 ( .IN1(n49), .IN2(n9), .IN3(n53), .Q(n54) );
  AOI22X1 U95 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n54), .QN(n52) );
  OA22X1 U96 ( .IN1(n67), .IN2(n9), .IN3(n141), .IN4(n50), .Q(n51) );
  NOR2X0 U97 ( .IN1(in2[9]), .IN2(n53), .QN(n57) );
  AO21X1 U98 ( .IN1(in2[9]), .IN2(n53), .IN3(n57), .Q(n58) );
  OA22X1 U99 ( .IN1(n9), .IN2(n130), .IN3(n140), .IN4(n58), .Q(n56) );
  AOI22X1 U100 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n54), .QN(n55) );
  OA21X1 U101 ( .IN1(n57), .IN2(n10), .IN3(n61), .Q(n62) );
  AOI22X1 U102 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n62), .QN(n60) );
  OA22X1 U103 ( .IN1(n67), .IN2(n10), .IN3(n141), .IN4(n58), .Q(n59) );
  NOR2X0 U104 ( .IN1(in2[11]), .IN2(n61), .QN(n65) );
  AO21X1 U105 ( .IN1(in2[11]), .IN2(n61), .IN3(n65), .Q(n66) );
  OA22X1 U106 ( .IN1(n10), .IN2(n130), .IN3(n140), .IN4(n66), .Q(n64) );
  AOI22X1 U107 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n62), .QN(n63) );
  OA21X1 U108 ( .IN1(n65), .IN2(n11), .IN3(n77), .Q(n70) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n70), .QN(n69) );
  OA22X1 U110 ( .IN1(n67), .IN2(n11), .IN3(n141), .IN4(n66), .Q(n68) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n12), .S(n71), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n11), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n13), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n12), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n12), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n14), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n13), .IN4(n85), .IN5(n84), 
        .Q(out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n15), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n14), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n14), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n16), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n15), .IN4(n97), .IN5(n96), 
        .Q(out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n17), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n16), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n16), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n18), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n17), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n19), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n18), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n18), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n20), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n19), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n21), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n20), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n20), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n21), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_49 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n25), .IN2(n6), .QN(n30) );
  NAND2X0 U4 ( .IN1(n33), .IN2(n7), .QN(n37) );
  NAND2X0 U5 ( .IN1(n41), .IN2(n8), .QN(n45) );
  NAND2X0 U6 ( .IN1(n49), .IN2(n9), .QN(n53) );
  NAND2X0 U7 ( .IN1(n57), .IN2(n10), .QN(n61) );
  NAND2X0 U8 ( .IN1(n65), .IN2(n11), .QN(n77) );
  NAND2X0 U9 ( .IN1(n81), .IN2(n13), .QN(n89) );
  NAND2X0 U10 ( .IN1(n93), .IN2(n15), .QN(n101) );
  NAND2X0 U11 ( .IN1(n105), .IN2(n17), .QN(n114) );
  NAND2X0 U12 ( .IN1(n118), .IN2(n19), .QN(n125) );
  NAND2X0 U13 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U14 ( .IN1(in1[2]), .IN2(n77), .QN(n71) );
  NAND2X0 U15 ( .IN1(n70), .IN2(n132), .QN(n74) );
  NAND2X0 U16 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U17 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U18 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U19 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U20 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U21 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U22 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U23 ( .IN1(n23), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U24 ( .IN1(in1[2]), .IN2(n22), .QN(n23) );
  NAND2X0 U25 ( .IN1(n32), .IN2(n31), .QN(out1[3]) );
  NAND2X0 U26 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U27 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U28 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NAND2X0 U29 ( .IN1(n27), .IN2(n132), .QN(n4) );
  NAND2X0 U30 ( .IN1(n36), .IN2(n35), .QN(out1[4]) );
  NAND2X0 U31 ( .IN1(n40), .IN2(n39), .QN(out1[5]) );
  NAND2X0 U32 ( .IN1(n44), .IN2(n43), .QN(out1[6]) );
  NAND2X0 U33 ( .IN1(n48), .IN2(n47), .QN(out1[7]) );
  NAND2X0 U34 ( .IN1(n52), .IN2(n51), .QN(out1[8]) );
  NAND2X0 U35 ( .IN1(n56), .IN2(n55), .QN(out1[9]) );
  NAND2X0 U36 ( .IN1(n60), .IN2(n59), .QN(out1[10]) );
  NAND2X0 U37 ( .IN1(n64), .IN2(n63), .QN(out1[11]) );
  NAND2X0 U38 ( .IN1(n69), .IN2(n68), .QN(out1[12]) );
  NAND2X0 U39 ( .IN1(n141), .IN2(n130), .QN(n24) );
  NOR2X0 U40 ( .IN1(n28), .IN2(n26), .QN(n3) );
  NOR2X0 U41 ( .IN1(n142), .IN2(n21), .QN(n1) );
  INVX0 U42 ( .INP(n132), .ZN(n141) );
  INVX0 U43 ( .INP(n130), .ZN(n137) );
  NAND3X0 U44 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  NOR3X0 U45 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  NOR2X0 U46 ( .IN1(n142), .IN2(n111), .QN(n138) );
  MUX21X1 U47 ( .IN1(n22), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  INVX0 U48 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U49 ( .INP(in2[2]), .ZN(n6) );
  INVX0 U50 ( .INP(in2[4]), .ZN(n7) );
  INVX0 U51 ( .INP(in2[6]), .ZN(n8) );
  INVX0 U52 ( .INP(in2[8]), .ZN(n9) );
  INVX0 U53 ( .INP(in2[10]), .ZN(n10) );
  INVX0 U54 ( .INP(in2[12]), .ZN(n11) );
  INVX0 U55 ( .INP(in2[13]), .ZN(n12) );
  INVX0 U56 ( .INP(in2[14]), .ZN(n13) );
  INVX0 U57 ( .INP(in2[15]), .ZN(n14) );
  INVX0 U58 ( .INP(in2[16]), .ZN(n15) );
  INVX0 U59 ( .INP(in2[17]), .ZN(n16) );
  INVX0 U60 ( .INP(in2[18]), .ZN(n17) );
  INVX0 U61 ( .INP(in2[19]), .ZN(n18) );
  INVX0 U62 ( .INP(in2[20]), .ZN(n19) );
  INVX0 U63 ( .INP(in2[21]), .ZN(n20) );
  INVX0 U64 ( .INP(in2[22]), .ZN(n21) );
  INVX0 U65 ( .INP(in1[1]), .ZN(n22) );
  INVX0 U66 ( .INP(in1[2]), .ZN(n111) );
  INVX0 U67 ( .INP(n138), .ZN(n140) );
  NOR2X0 U68 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n25) );
  AOI21X1 U69 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n25), .QN(n27) );
  NOR2X0 U70 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U71 ( .IN1(n24), .IN2(in2[0]), .IN3(n138), .IN4(n27), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U72 ( .INP(n133), .ZN(n67) );
  NOR2X0 U73 ( .IN1(n67), .IN2(n6), .QN(n28) );
  OA21X1 U74 ( .IN1(n25), .IN2(n6), .IN3(n30), .Q(n29) );
  AO22X1 U75 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n29), .Q(n26) );
  AOI22X1 U76 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n29), .QN(n32) );
  NOR2X0 U77 ( .IN1(in2[3]), .IN2(n30), .QN(n33) );
  AO21X1 U78 ( .IN1(in2[3]), .IN2(n30), .IN3(n33), .Q(n34) );
  OA22X1 U79 ( .IN1(n6), .IN2(n130), .IN3(n140), .IN4(n34), .Q(n31) );
  OA21X1 U80 ( .IN1(n33), .IN2(n7), .IN3(n37), .Q(n38) );
  AOI22X1 U81 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n38), .QN(n36) );
  OA22X1 U82 ( .IN1(n67), .IN2(n7), .IN3(n141), .IN4(n34), .Q(n35) );
  NOR2X0 U83 ( .IN1(in2[5]), .IN2(n37), .QN(n41) );
  AO21X1 U84 ( .IN1(in2[5]), .IN2(n37), .IN3(n41), .Q(n42) );
  OA22X1 U85 ( .IN1(n7), .IN2(n130), .IN3(n140), .IN4(n42), .Q(n40) );
  AOI22X1 U86 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n38), .QN(n39) );
  OA21X1 U87 ( .IN1(n41), .IN2(n8), .IN3(n45), .Q(n46) );
  AOI22X1 U88 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n46), .QN(n44) );
  OA22X1 U89 ( .IN1(n67), .IN2(n8), .IN3(n141), .IN4(n42), .Q(n43) );
  NOR2X0 U90 ( .IN1(in2[7]), .IN2(n45), .QN(n49) );
  AO21X1 U91 ( .IN1(in2[7]), .IN2(n45), .IN3(n49), .Q(n50) );
  OA22X1 U92 ( .IN1(n8), .IN2(n130), .IN3(n140), .IN4(n50), .Q(n48) );
  AOI22X1 U93 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n46), .QN(n47) );
  OA21X1 U94 ( .IN1(n49), .IN2(n9), .IN3(n53), .Q(n54) );
  AOI22X1 U95 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n54), .QN(n52) );
  OA22X1 U96 ( .IN1(n67), .IN2(n9), .IN3(n141), .IN4(n50), .Q(n51) );
  NOR2X0 U97 ( .IN1(in2[9]), .IN2(n53), .QN(n57) );
  AO21X1 U98 ( .IN1(in2[9]), .IN2(n53), .IN3(n57), .Q(n58) );
  OA22X1 U99 ( .IN1(n9), .IN2(n130), .IN3(n140), .IN4(n58), .Q(n56) );
  AOI22X1 U100 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n54), .QN(n55) );
  OA21X1 U101 ( .IN1(n57), .IN2(n10), .IN3(n61), .Q(n62) );
  AOI22X1 U102 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n62), .QN(n60) );
  OA22X1 U103 ( .IN1(n67), .IN2(n10), .IN3(n141), .IN4(n58), .Q(n59) );
  NOR2X0 U104 ( .IN1(in2[11]), .IN2(n61), .QN(n65) );
  AO21X1 U105 ( .IN1(in2[11]), .IN2(n61), .IN3(n65), .Q(n66) );
  OA22X1 U106 ( .IN1(n10), .IN2(n130), .IN3(n140), .IN4(n66), .Q(n64) );
  AOI22X1 U107 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n62), .QN(n63) );
  OA21X1 U108 ( .IN1(n65), .IN2(n11), .IN3(n77), .Q(n70) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n70), .QN(n69) );
  OA22X1 U110 ( .IN1(n67), .IN2(n11), .IN3(n141), .IN4(n66), .Q(n68) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n12), .S(n71), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n11), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n13), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n12), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n12), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n14), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n13), .IN4(n85), .IN5(n84), 
        .Q(out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n15), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n14), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n14), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n16), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n15), .IN4(n97), .IN5(n96), 
        .Q(out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n17), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n16), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n16), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n18), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n17), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n19), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n18), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n18), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n20), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n19), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n21), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n20), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n20), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n21), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_50 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n25), .IN2(n6), .QN(n30) );
  NAND2X0 U4 ( .IN1(n33), .IN2(n7), .QN(n37) );
  NAND2X0 U5 ( .IN1(n41), .IN2(n8), .QN(n45) );
  NAND2X0 U6 ( .IN1(n49), .IN2(n9), .QN(n53) );
  NAND2X0 U7 ( .IN1(n57), .IN2(n10), .QN(n61) );
  NAND2X0 U8 ( .IN1(n65), .IN2(n11), .QN(n77) );
  NAND2X0 U9 ( .IN1(n81), .IN2(n13), .QN(n89) );
  NAND2X0 U10 ( .IN1(n105), .IN2(n17), .QN(n114) );
  NAND2X0 U11 ( .IN1(n93), .IN2(n15), .QN(n101) );
  NAND2X0 U12 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U13 ( .IN1(n118), .IN2(n19), .QN(n125) );
  NAND2X0 U14 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U15 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U16 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U17 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U18 ( .IN1(n27), .IN2(n132), .QN(n4) );
  NAND2X0 U19 ( .IN1(n141), .IN2(n130), .QN(n24) );
  NAND2X0 U20 ( .IN1(n32), .IN2(n31), .QN(out1[3]) );
  NAND2X0 U21 ( .IN1(n36), .IN2(n35), .QN(out1[4]) );
  NAND2X0 U22 ( .IN1(in1[2]), .IN2(n77), .QN(n71) );
  NAND2X0 U23 ( .IN1(n70), .IN2(n132), .QN(n74) );
  NAND2X0 U24 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U25 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U26 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U27 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U28 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NAND2X0 U29 ( .IN1(n40), .IN2(n39), .QN(out1[5]) );
  NAND2X0 U30 ( .IN1(n44), .IN2(n43), .QN(out1[6]) );
  NAND2X0 U31 ( .IN1(n48), .IN2(n47), .QN(out1[7]) );
  NAND2X0 U32 ( .IN1(n52), .IN2(n51), .QN(out1[8]) );
  NAND2X0 U33 ( .IN1(n56), .IN2(n55), .QN(out1[9]) );
  NAND2X0 U34 ( .IN1(n60), .IN2(n59), .QN(out1[10]) );
  NAND2X0 U35 ( .IN1(n64), .IN2(n63), .QN(out1[11]) );
  NAND2X0 U36 ( .IN1(n69), .IN2(n68), .QN(out1[12]) );
  NAND2X0 U37 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U38 ( .IN1(n23), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U39 ( .IN1(in1[2]), .IN2(n22), .QN(n23) );
  INVX0 U40 ( .INP(in1[2]), .ZN(n111) );
  NOR2X0 U41 ( .IN1(n28), .IN2(n26), .QN(n3) );
  NOR2X0 U42 ( .IN1(n142), .IN2(n21), .QN(n1) );
  INVX0 U43 ( .INP(n132), .ZN(n141) );
  INVX0 U44 ( .INP(n130), .ZN(n137) );
  NAND3X0 U45 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  NOR3X0 U46 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  NOR2X0 U47 ( .IN1(n142), .IN2(n111), .QN(n138) );
  MUX21X1 U48 ( .IN1(n22), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  INVX0 U49 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U50 ( .INP(in2[2]), .ZN(n6) );
  INVX0 U51 ( .INP(in2[4]), .ZN(n7) );
  INVX0 U52 ( .INP(in2[6]), .ZN(n8) );
  INVX0 U53 ( .INP(in2[8]), .ZN(n9) );
  INVX0 U54 ( .INP(in2[10]), .ZN(n10) );
  INVX0 U55 ( .INP(in2[12]), .ZN(n11) );
  INVX0 U56 ( .INP(in2[13]), .ZN(n12) );
  INVX0 U57 ( .INP(in2[14]), .ZN(n13) );
  INVX0 U58 ( .INP(in2[15]), .ZN(n14) );
  INVX0 U59 ( .INP(in2[16]), .ZN(n15) );
  INVX0 U60 ( .INP(in2[17]), .ZN(n16) );
  INVX0 U61 ( .INP(in2[18]), .ZN(n17) );
  INVX0 U62 ( .INP(in2[19]), .ZN(n18) );
  INVX0 U63 ( .INP(in2[20]), .ZN(n19) );
  INVX0 U64 ( .INP(in2[21]), .ZN(n20) );
  INVX0 U65 ( .INP(in2[22]), .ZN(n21) );
  INVX0 U66 ( .INP(in1[1]), .ZN(n22) );
  INVX0 U67 ( .INP(n138), .ZN(n140) );
  NOR2X0 U68 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n25) );
  AOI21X1 U69 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n25), .QN(n27) );
  NOR2X0 U70 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U71 ( .IN1(n24), .IN2(in2[0]), .IN3(n138), .IN4(n27), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U72 ( .INP(n133), .ZN(n67) );
  NOR2X0 U73 ( .IN1(n67), .IN2(n6), .QN(n28) );
  OA21X1 U74 ( .IN1(n25), .IN2(n6), .IN3(n30), .Q(n29) );
  AO22X1 U75 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n29), .Q(n26) );
  AOI22X1 U76 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n29), .QN(n32) );
  NOR2X0 U77 ( .IN1(in2[3]), .IN2(n30), .QN(n33) );
  AO21X1 U78 ( .IN1(in2[3]), .IN2(n30), .IN3(n33), .Q(n34) );
  OA22X1 U79 ( .IN1(n6), .IN2(n130), .IN3(n140), .IN4(n34), .Q(n31) );
  OA21X1 U80 ( .IN1(n33), .IN2(n7), .IN3(n37), .Q(n38) );
  AOI22X1 U81 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n38), .QN(n36) );
  OA22X1 U82 ( .IN1(n67), .IN2(n7), .IN3(n141), .IN4(n34), .Q(n35) );
  NOR2X0 U83 ( .IN1(in2[5]), .IN2(n37), .QN(n41) );
  AO21X1 U84 ( .IN1(in2[5]), .IN2(n37), .IN3(n41), .Q(n42) );
  OA22X1 U85 ( .IN1(n7), .IN2(n130), .IN3(n140), .IN4(n42), .Q(n40) );
  AOI22X1 U86 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n38), .QN(n39) );
  OA21X1 U87 ( .IN1(n41), .IN2(n8), .IN3(n45), .Q(n46) );
  AOI22X1 U88 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n46), .QN(n44) );
  OA22X1 U89 ( .IN1(n67), .IN2(n8), .IN3(n141), .IN4(n42), .Q(n43) );
  NOR2X0 U90 ( .IN1(in2[7]), .IN2(n45), .QN(n49) );
  AO21X1 U91 ( .IN1(in2[7]), .IN2(n45), .IN3(n49), .Q(n50) );
  OA22X1 U92 ( .IN1(n8), .IN2(n130), .IN3(n140), .IN4(n50), .Q(n48) );
  AOI22X1 U93 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n46), .QN(n47) );
  OA21X1 U94 ( .IN1(n49), .IN2(n9), .IN3(n53), .Q(n54) );
  AOI22X1 U95 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n54), .QN(n52) );
  OA22X1 U96 ( .IN1(n67), .IN2(n9), .IN3(n141), .IN4(n50), .Q(n51) );
  NOR2X0 U97 ( .IN1(in2[9]), .IN2(n53), .QN(n57) );
  AO21X1 U98 ( .IN1(in2[9]), .IN2(n53), .IN3(n57), .Q(n58) );
  OA22X1 U99 ( .IN1(n9), .IN2(n130), .IN3(n140), .IN4(n58), .Q(n56) );
  AOI22X1 U100 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n54), .QN(n55) );
  OA21X1 U101 ( .IN1(n57), .IN2(n10), .IN3(n61), .Q(n62) );
  AOI22X1 U102 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n62), .QN(n60) );
  OA22X1 U103 ( .IN1(n67), .IN2(n10), .IN3(n141), .IN4(n58), .Q(n59) );
  NOR2X0 U104 ( .IN1(in2[11]), .IN2(n61), .QN(n65) );
  AO21X1 U105 ( .IN1(in2[11]), .IN2(n61), .IN3(n65), .Q(n66) );
  OA22X1 U106 ( .IN1(n10), .IN2(n130), .IN3(n140), .IN4(n66), .Q(n64) );
  AOI22X1 U107 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n62), .QN(n63) );
  OA21X1 U108 ( .IN1(n65), .IN2(n11), .IN3(n77), .Q(n70) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n70), .QN(n69) );
  OA22X1 U110 ( .IN1(n67), .IN2(n11), .IN3(n141), .IN4(n66), .Q(n68) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n12), .S(n71), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n11), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n13), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n12), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n12), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n14), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n13), .IN4(n85), .IN5(n84), 
        .Q(out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n15), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n14), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n14), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n16), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n15), .IN4(n97), .IN5(n96), 
        .Q(out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n17), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n16), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n16), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n18), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n17), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n19), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n18), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n18), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n20), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n19), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n21), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n20), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n20), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n21), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_51 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n33), .IN2(n7), .QN(n37) );
  NAND2X0 U4 ( .IN1(n41), .IN2(n8), .QN(n45) );
  NAND2X0 U5 ( .IN1(n49), .IN2(n9), .QN(n53) );
  NAND2X0 U6 ( .IN1(n57), .IN2(n10), .QN(n61) );
  NAND2X0 U7 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U8 ( .IN1(n25), .IN2(n6), .QN(n30) );
  NAND2X0 U9 ( .IN1(n65), .IN2(n11), .QN(n77) );
  NAND2X0 U10 ( .IN1(n81), .IN2(n13), .QN(n89) );
  NAND2X0 U11 ( .IN1(n93), .IN2(n15), .QN(n101) );
  NAND2X0 U12 ( .IN1(n118), .IN2(n19), .QN(n125) );
  NAND2X0 U13 ( .IN1(n105), .IN2(n17), .QN(n114) );
  NAND2X0 U14 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U15 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U16 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U17 ( .IN1(n40), .IN2(n39), .QN(out1[5]) );
  NAND2X0 U18 ( .IN1(n44), .IN2(n43), .QN(out1[6]) );
  NAND2X0 U19 ( .IN1(in1[2]), .IN2(n77), .QN(n71) );
  NAND2X0 U20 ( .IN1(n70), .IN2(n132), .QN(n74) );
  NAND2X0 U21 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U22 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U23 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U24 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U25 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U26 ( .IN1(n23), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U27 ( .IN1(in1[2]), .IN2(n22), .QN(n23) );
  NAND2X0 U28 ( .IN1(n36), .IN2(n35), .QN(out1[4]) );
  NAND2X0 U29 ( .IN1(n32), .IN2(n31), .QN(out1[3]) );
  NAND2X0 U30 ( .IN1(n27), .IN2(n132), .QN(n4) );
  NAND2X0 U31 ( .IN1(n48), .IN2(n47), .QN(out1[7]) );
  NAND2X0 U32 ( .IN1(n52), .IN2(n51), .QN(out1[8]) );
  NAND2X0 U33 ( .IN1(n56), .IN2(n55), .QN(out1[9]) );
  NAND2X0 U34 ( .IN1(n60), .IN2(n59), .QN(out1[10]) );
  NAND2X0 U35 ( .IN1(n64), .IN2(n63), .QN(out1[11]) );
  NAND2X0 U36 ( .IN1(n69), .IN2(n68), .QN(out1[12]) );
  NAND2X0 U37 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U38 ( .IN1(n141), .IN2(n130), .QN(n24) );
  NAND2X0 U39 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NOR2X0 U40 ( .IN1(n28), .IN2(n26), .QN(n3) );
  NOR2X0 U41 ( .IN1(n142), .IN2(n21), .QN(n1) );
  INVX0 U42 ( .INP(n132), .ZN(n141) );
  INVX0 U43 ( .INP(n130), .ZN(n137) );
  NAND3X0 U44 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  NOR3X0 U45 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  NOR2X0 U46 ( .IN1(n142), .IN2(n111), .QN(n138) );
  MUX21X1 U47 ( .IN1(n22), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  INVX0 U48 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U49 ( .INP(in2[2]), .ZN(n6) );
  INVX0 U50 ( .INP(in2[4]), .ZN(n7) );
  INVX0 U51 ( .INP(in2[6]), .ZN(n8) );
  INVX0 U52 ( .INP(in2[8]), .ZN(n9) );
  INVX0 U53 ( .INP(in2[10]), .ZN(n10) );
  INVX0 U54 ( .INP(in2[12]), .ZN(n11) );
  INVX0 U55 ( .INP(in2[13]), .ZN(n12) );
  INVX0 U56 ( .INP(in2[14]), .ZN(n13) );
  INVX0 U57 ( .INP(in2[15]), .ZN(n14) );
  INVX0 U58 ( .INP(in2[16]), .ZN(n15) );
  INVX0 U59 ( .INP(in2[17]), .ZN(n16) );
  INVX0 U60 ( .INP(in2[18]), .ZN(n17) );
  INVX0 U61 ( .INP(in2[19]), .ZN(n18) );
  INVX0 U62 ( .INP(in2[20]), .ZN(n19) );
  INVX0 U63 ( .INP(in2[21]), .ZN(n20) );
  INVX0 U64 ( .INP(in2[22]), .ZN(n21) );
  INVX0 U65 ( .INP(in1[1]), .ZN(n22) );
  INVX0 U66 ( .INP(in1[2]), .ZN(n111) );
  INVX0 U67 ( .INP(n138), .ZN(n140) );
  NOR2X0 U68 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n25) );
  AOI21X1 U69 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n25), .QN(n27) );
  NOR2X0 U70 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U71 ( .IN1(n24), .IN2(in2[0]), .IN3(n138), .IN4(n27), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U72 ( .INP(n133), .ZN(n67) );
  NOR2X0 U73 ( .IN1(n67), .IN2(n6), .QN(n28) );
  OA21X1 U74 ( .IN1(n25), .IN2(n6), .IN3(n30), .Q(n29) );
  AO22X1 U75 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n29), .Q(n26) );
  AOI22X1 U76 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n29), .QN(n32) );
  NOR2X0 U77 ( .IN1(in2[3]), .IN2(n30), .QN(n33) );
  AO21X1 U78 ( .IN1(in2[3]), .IN2(n30), .IN3(n33), .Q(n34) );
  OA22X1 U79 ( .IN1(n6), .IN2(n130), .IN3(n140), .IN4(n34), .Q(n31) );
  OA21X1 U80 ( .IN1(n33), .IN2(n7), .IN3(n37), .Q(n38) );
  AOI22X1 U81 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n38), .QN(n36) );
  OA22X1 U82 ( .IN1(n67), .IN2(n7), .IN3(n141), .IN4(n34), .Q(n35) );
  NOR2X0 U83 ( .IN1(in2[5]), .IN2(n37), .QN(n41) );
  AO21X1 U84 ( .IN1(in2[5]), .IN2(n37), .IN3(n41), .Q(n42) );
  OA22X1 U85 ( .IN1(n7), .IN2(n130), .IN3(n140), .IN4(n42), .Q(n40) );
  AOI22X1 U86 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n38), .QN(n39) );
  OA21X1 U87 ( .IN1(n41), .IN2(n8), .IN3(n45), .Q(n46) );
  AOI22X1 U88 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n46), .QN(n44) );
  OA22X1 U89 ( .IN1(n67), .IN2(n8), .IN3(n141), .IN4(n42), .Q(n43) );
  NOR2X0 U90 ( .IN1(in2[7]), .IN2(n45), .QN(n49) );
  AO21X1 U91 ( .IN1(in2[7]), .IN2(n45), .IN3(n49), .Q(n50) );
  OA22X1 U92 ( .IN1(n8), .IN2(n130), .IN3(n140), .IN4(n50), .Q(n48) );
  AOI22X1 U93 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n46), .QN(n47) );
  OA21X1 U94 ( .IN1(n49), .IN2(n9), .IN3(n53), .Q(n54) );
  AOI22X1 U95 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n54), .QN(n52) );
  OA22X1 U96 ( .IN1(n67), .IN2(n9), .IN3(n141), .IN4(n50), .Q(n51) );
  NOR2X0 U97 ( .IN1(in2[9]), .IN2(n53), .QN(n57) );
  AO21X1 U98 ( .IN1(in2[9]), .IN2(n53), .IN3(n57), .Q(n58) );
  OA22X1 U99 ( .IN1(n9), .IN2(n130), .IN3(n140), .IN4(n58), .Q(n56) );
  AOI22X1 U100 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n54), .QN(n55) );
  OA21X1 U101 ( .IN1(n57), .IN2(n10), .IN3(n61), .Q(n62) );
  AOI22X1 U102 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n62), .QN(n60) );
  OA22X1 U103 ( .IN1(n67), .IN2(n10), .IN3(n141), .IN4(n58), .Q(n59) );
  NOR2X0 U104 ( .IN1(in2[11]), .IN2(n61), .QN(n65) );
  AO21X1 U105 ( .IN1(in2[11]), .IN2(n61), .IN3(n65), .Q(n66) );
  OA22X1 U106 ( .IN1(n10), .IN2(n130), .IN3(n140), .IN4(n66), .Q(n64) );
  AOI22X1 U107 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n62), .QN(n63) );
  OA21X1 U108 ( .IN1(n65), .IN2(n11), .IN3(n77), .Q(n70) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n70), .QN(n69) );
  OA22X1 U110 ( .IN1(n67), .IN2(n11), .IN3(n141), .IN4(n66), .Q(n68) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n12), .S(n71), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n11), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n13), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n12), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n12), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n14), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n13), .IN4(n85), .IN5(n84), 
        .Q(out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n15), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n14), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n14), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n16), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n15), .IN4(n97), .IN5(n96), 
        .Q(out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n17), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n16), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n16), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n18), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n17), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n19), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n18), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n18), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n20), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n19), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n21), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n20), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n20), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n21), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_52 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93;

  NAND2X0 U3 ( .IN1(n30), .IN2(n7), .QN(n32) );
  NAND2X0 U4 ( .IN1(n34), .IN2(n8), .QN(n36) );
  NAND2X0 U5 ( .IN1(n38), .IN2(n9), .QN(n40) );
  NAND2X0 U6 ( .IN1(n42), .IN2(n10), .QN(n47) );
  NAND2X0 U7 ( .IN1(n78), .IN2(n18), .QN(n82) );
  NAND2X0 U8 ( .IN1(n26), .IN2(n6), .QN(n28) );
  NAND2X0 U9 ( .IN1(in1[2]), .IN2(n47), .QN(n44) );
  NAND2X0 U10 ( .IN1(n52), .IN2(n12), .QN(n55) );
  NAND2X0 U11 ( .IN1(in1[2]), .IN2(n55), .QN(n51) );
  NAND2X0 U12 ( .IN1(n60), .IN2(n14), .QN(n63) );
  NAND2X0 U13 ( .IN1(in1[2]), .IN2(n63), .QN(n59) );
  NAND2X0 U14 ( .IN1(n68), .IN2(n16), .QN(n71) );
  NAND2X0 U15 ( .IN1(in1[2]), .IN2(n71), .QN(n67) );
  NAND2X0 U16 ( .IN1(in1[2]), .IN2(n82), .QN(n77) );
  NAND2X0 U17 ( .IN1(in2[21]), .IN2(n82), .QN(n83) );
  NAND2X0 U18 ( .IN1(n75), .IN2(in1[2]), .QN(n86) );
  NAND2X0 U19 ( .IN1(n3), .IN2(n4), .QN(n22) );
  NAND2X0 U20 ( .IN1(in2[1]), .IN2(in2[0]), .QN(n4) );
  NAND2X0 U21 ( .IN1(n23), .IN2(n22), .QN(out1[2]) );
  INVX0 U22 ( .INP(n86), .ZN(n89) );
  NOR2X0 U23 ( .IN1(n21), .IN2(n86), .QN(n3) );
  NOR2X0 U24 ( .IN1(in1[2]), .IN2(n75), .QN(n90) );
  NOR2X0 U25 ( .IN1(n75), .IN2(n72), .QN(n92) );
  NBUFFX2 U26 ( .INP(in1[2]), .Z(out1[26]) );
  NBUFFX2 U27 ( .INP(in1[2]), .Z(out1[25]) );
  INVX0 U28 ( .INP(in2[2]), .ZN(n5) );
  INVX0 U29 ( .INP(in2[4]), .ZN(n6) );
  INVX0 U30 ( .INP(in2[6]), .ZN(n7) );
  INVX0 U31 ( .INP(in2[8]), .ZN(n8) );
  INVX0 U32 ( .INP(in2[10]), .ZN(n9) );
  INVX0 U33 ( .INP(in2[12]), .ZN(n10) );
  INVX0 U34 ( .INP(in2[13]), .ZN(n11) );
  INVX0 U35 ( .INP(in2[14]), .ZN(n12) );
  INVX0 U36 ( .INP(in2[15]), .ZN(n13) );
  INVX0 U37 ( .INP(in2[16]), .ZN(n14) );
  INVX0 U38 ( .INP(in2[17]), .ZN(n15) );
  INVX0 U39 ( .INP(in2[18]), .ZN(n16) );
  INVX0 U40 ( .INP(in2[19]), .ZN(n17) );
  INVX0 U41 ( .INP(in2[20]), .ZN(n18) );
  INVX0 U42 ( .INP(in2[21]), .ZN(n19) );
  INVX0 U43 ( .INP(in2[22]), .ZN(n20) );
  INVX0 U44 ( .INP(in1[1]), .ZN(n75) );
  INVX0 U45 ( .INP(in1[2]), .ZN(n72) );
  NOR2X0 U46 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n21) );
  OR3X1 U47 ( .IN1(in2[2]), .IN2(in2[0]), .IN3(in2[1]), .Q(n24) );
  OA21X1 U48 ( .IN1(n21), .IN2(n5), .IN3(n24), .Q(n25) );
  AOI22X1 U49 ( .IN1(in2[2]), .IN2(n90), .IN3(n92), .IN4(n25), .QN(n23) );
  NOR2X0 U50 ( .IN1(in2[3]), .IN2(n24), .QN(n26) );
  AOI21X1 U51 ( .IN1(in2[3]), .IN2(n24), .IN3(n26), .QN(n27) );
  AO222X1 U52 ( .IN1(in2[3]), .IN2(n90), .IN3(n92), .IN4(n27), .IN5(n89), 
        .IN6(n25), .Q(out1[3]) );
  OA21X1 U53 ( .IN1(n26), .IN2(n6), .IN3(n28), .Q(n29) );
  AO222X1 U54 ( .IN1(in2[4]), .IN2(n90), .IN3(n92), .IN4(n29), .IN5(n89), 
        .IN6(n27), .Q(out1[4]) );
  NOR2X0 U55 ( .IN1(in2[5]), .IN2(n28), .QN(n30) );
  AOI21X1 U56 ( .IN1(in2[5]), .IN2(n28), .IN3(n30), .QN(n31) );
  AO222X1 U57 ( .IN1(in2[5]), .IN2(n90), .IN3(n92), .IN4(n31), .IN5(n89), 
        .IN6(n29), .Q(out1[5]) );
  OA21X1 U58 ( .IN1(n30), .IN2(n7), .IN3(n32), .Q(n33) );
  AO222X1 U59 ( .IN1(in2[6]), .IN2(n90), .IN3(n92), .IN4(n33), .IN5(n89), 
        .IN6(n31), .Q(out1[6]) );
  NOR2X0 U60 ( .IN1(in2[7]), .IN2(n32), .QN(n34) );
  AOI21X1 U61 ( .IN1(in2[7]), .IN2(n32), .IN3(n34), .QN(n35) );
  AO222X1 U62 ( .IN1(in2[7]), .IN2(n90), .IN3(n92), .IN4(n35), .IN5(n89), 
        .IN6(n33), .Q(out1[7]) );
  OA21X1 U63 ( .IN1(n34), .IN2(n8), .IN3(n36), .Q(n37) );
  AO222X1 U64 ( .IN1(in2[8]), .IN2(n90), .IN3(n92), .IN4(n37), .IN5(n89), 
        .IN6(n35), .Q(out1[8]) );
  NOR2X0 U65 ( .IN1(in2[9]), .IN2(n36), .QN(n38) );
  AOI21X1 U66 ( .IN1(in2[9]), .IN2(n36), .IN3(n38), .QN(n39) );
  AO222X1 U67 ( .IN1(in2[9]), .IN2(n90), .IN3(n92), .IN4(n39), .IN5(n89), 
        .IN6(n37), .Q(out1[9]) );
  OA21X1 U68 ( .IN1(n38), .IN2(n9), .IN3(n40), .Q(n41) );
  AO222X1 U69 ( .IN1(in2[10]), .IN2(n90), .IN3(n92), .IN4(n41), .IN5(n89), 
        .IN6(n39), .Q(out1[10]) );
  NOR2X0 U70 ( .IN1(in2[11]), .IN2(n40), .QN(n42) );
  AOI21X1 U71 ( .IN1(in2[11]), .IN2(n40), .IN3(n42), .QN(n43) );
  AO222X1 U72 ( .IN1(in2[11]), .IN2(n90), .IN3(n92), .IN4(n43), .IN5(n89), 
        .IN6(n41), .Q(out1[11]) );
  OA21X1 U73 ( .IN1(n42), .IN2(n10), .IN3(n47), .Q(n45) );
  AO222X1 U74 ( .IN1(in2[12]), .IN2(n90), .IN3(n92), .IN4(n45), .IN5(n89), 
        .IN6(n43), .Q(out1[12]) );
  MUX21X1 U75 ( .IN1(n11), .IN2(in2[13]), .S(n44), .Q(n46) );
  AO22X1 U76 ( .IN1(in1[1]), .IN2(n46), .IN3(n89), .IN4(n45), .Q(out1[13]) );
  NOR2X0 U77 ( .IN1(in2[13]), .IN2(n47), .QN(n52) );
  AO21X1 U78 ( .IN1(in2[13]), .IN2(n47), .IN3(n86), .Q(n50) );
  NOR2X0 U79 ( .IN1(n52), .IN2(n72), .QN(n48) );
  MUX21X1 U80 ( .IN1(n12), .IN2(in2[14]), .S(n48), .Q(n49) );
  OAI22X1 U81 ( .IN1(n52), .IN2(n50), .IN3(n75), .IN4(n49), .QN(out1[14]) );
  MUX21X1 U82 ( .IN1(n13), .IN2(in2[15]), .S(n51), .Q(n54) );
  OA21X1 U83 ( .IN1(n52), .IN2(n12), .IN3(n89), .Q(n53) );
  AO22X1 U84 ( .IN1(in1[1]), .IN2(n54), .IN3(n53), .IN4(n55), .Q(out1[15]) );
  NOR2X0 U85 ( .IN1(in2[15]), .IN2(n55), .QN(n60) );
  AO21X1 U86 ( .IN1(in2[15]), .IN2(n55), .IN3(n86), .Q(n58) );
  NOR2X0 U87 ( .IN1(n60), .IN2(n72), .QN(n56) );
  MUX21X1 U88 ( .IN1(n14), .IN2(in2[16]), .S(n56), .Q(n57) );
  OAI22X1 U89 ( .IN1(n60), .IN2(n58), .IN3(n75), .IN4(n57), .QN(out1[16]) );
  MUX21X1 U90 ( .IN1(n15), .IN2(in2[17]), .S(n59), .Q(n62) );
  OA21X1 U91 ( .IN1(n60), .IN2(n14), .IN3(n89), .Q(n61) );
  AO22X1 U92 ( .IN1(in1[1]), .IN2(n62), .IN3(n61), .IN4(n63), .Q(out1[17]) );
  NOR2X0 U93 ( .IN1(in2[17]), .IN2(n63), .QN(n68) );
  AO21X1 U94 ( .IN1(in2[17]), .IN2(n63), .IN3(n86), .Q(n66) );
  NOR2X0 U95 ( .IN1(n68), .IN2(n72), .QN(n64) );
  MUX21X1 U96 ( .IN1(n16), .IN2(in2[18]), .S(n64), .Q(n65) );
  OAI22X1 U97 ( .IN1(n68), .IN2(n66), .IN3(n75), .IN4(n65), .QN(out1[18]) );
  MUX21X1 U98 ( .IN1(n17), .IN2(in2[19]), .S(n67), .Q(n70) );
  OA21X1 U99 ( .IN1(n68), .IN2(n16), .IN3(n89), .Q(n69) );
  AO22X1 U100 ( .IN1(in1[1]), .IN2(n70), .IN3(n69), .IN4(n71), .Q(out1[19]) );
  NOR2X0 U101 ( .IN1(in2[19]), .IN2(n71), .QN(n78) );
  AO21X1 U102 ( .IN1(in2[19]), .IN2(n71), .IN3(n86), .Q(n76) );
  NOR2X0 U103 ( .IN1(n78), .IN2(n72), .QN(n73) );
  MUX21X1 U104 ( .IN1(n18), .IN2(in2[20]), .S(n73), .Q(n74) );
  OAI22X1 U105 ( .IN1(n78), .IN2(n76), .IN3(n75), .IN4(n74), .QN(out1[20]) );
  MUX21X1 U106 ( .IN1(n19), .IN2(in2[21]), .S(n77), .Q(n80) );
  MUX21X1 U107 ( .IN1(n18), .IN2(in2[20]), .S(n78), .Q(n79) );
  AO22X1 U108 ( .IN1(in1[1]), .IN2(n80), .IN3(n89), .IN4(n79), .Q(out1[21]) );
  INVX0 U109 ( .INP(n92), .ZN(n81) );
  OR2X1 U110 ( .IN1(n82), .IN2(in2[21]), .Q(n88) );
  NOR2X0 U111 ( .IN1(n81), .IN2(n88), .QN(n87) );
  NOR2X0 U112 ( .IN1(in2[22]), .IN2(n81), .QN(n84) );
  OA221X1 U113 ( .IN1(n84), .IN2(n89), .IN3(n84), .IN4(n83), .IN5(n88), .Q(n85) );
  AO221X1 U114 ( .IN1(in2[22]), .IN2(n87), .IN3(in2[22]), .IN4(n90), .IN5(n85), 
        .Q(out1[22]) );
  NOR2X0 U115 ( .IN1(n86), .IN2(n88), .QN(n93) );
  AO21X1 U116 ( .IN1(n89), .IN2(n88), .IN3(n87), .Q(n91) );
  AO221X1 U117 ( .IN1(in2[22]), .IN2(n93), .IN3(n20), .IN4(n91), .IN5(n90), 
        .Q(out1[23]) );
  AO21X1 U118 ( .IN1(n93), .IN2(n20), .IN3(n92), .Q(out1[24]) );
endmodule


module mul26_4 ( clk, rst_n, in1, in2, en, mulout );
  input [25:0] in1;
  input [25:0] in2;
  output [50:0] mulout;
  input clk, rst_n, en;
  wire   N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24,
         N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38,
         N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N62, N63,
         N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77,
         N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91,
         N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n131, n132, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22,
         SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24,
         SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26,
         SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28,
         SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30,
         SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32,
         SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34,
         SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36,
         SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38,
         SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40,
         SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42,
         SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44,
         SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46,
         SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48,
         SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50,
         SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52,
         SYNOPSYS_UNCONNECTED_53, SYNOPSYS_UNCONNECTED_54,
         SYNOPSYS_UNCONNECTED_55, SYNOPSYS_UNCONNECTED_56,
         SYNOPSYS_UNCONNECTED_57, SYNOPSYS_UNCONNECTED_58,
         SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_60,
         SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_62,
         SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_64,
         SYNOPSYS_UNCONNECTED_65, SYNOPSYS_UNCONNECTED_66,
         SYNOPSYS_UNCONNECTED_67, SYNOPSYS_UNCONNECTED_68,
         SYNOPSYS_UNCONNECTED_69, SYNOPSYS_UNCONNECTED_70,
         SYNOPSYS_UNCONNECTED_71, SYNOPSYS_UNCONNECTED_72,
         SYNOPSYS_UNCONNECTED_73, SYNOPSYS_UNCONNECTED_74,
         SYNOPSYS_UNCONNECTED_75, SYNOPSYS_UNCONNECTED_76,
         SYNOPSYS_UNCONNECTED_77, SYNOPSYS_UNCONNECTED_78,
         SYNOPSYS_UNCONNECTED_79, SYNOPSYS_UNCONNECTED_80,
         SYNOPSYS_UNCONNECTED_81, SYNOPSYS_UNCONNECTED_82,
         SYNOPSYS_UNCONNECTED_83, SYNOPSYS_UNCONNECTED_84,
         SYNOPSYS_UNCONNECTED_85, SYNOPSYS_UNCONNECTED_86,
         SYNOPSYS_UNCONNECTED_87, SYNOPSYS_UNCONNECTED_88,
         SYNOPSYS_UNCONNECTED_89, SYNOPSYS_UNCONNECTED_90,
         SYNOPSYS_UNCONNECTED_91, SYNOPSYS_UNCONNECTED_92,
         SYNOPSYS_UNCONNECTED_93, SYNOPSYS_UNCONNECTED_94,
         SYNOPSYS_UNCONNECTED_95, SYNOPSYS_UNCONNECTED_96,
         SYNOPSYS_UNCONNECTED_97, SYNOPSYS_UNCONNECTED_98,
         SYNOPSYS_UNCONNECTED_99, SYNOPSYS_UNCONNECTED_100,
         SYNOPSYS_UNCONNECTED_101, SYNOPSYS_UNCONNECTED_102,
         SYNOPSYS_UNCONNECTED_103, SYNOPSYS_UNCONNECTED_104,
         SYNOPSYS_UNCONNECTED_105, SYNOPSYS_UNCONNECTED_106,
         SYNOPSYS_UNCONNECTED_107, SYNOPSYS_UNCONNECTED_108,
         SYNOPSYS_UNCONNECTED_109, SYNOPSYS_UNCONNECTED_110,
         SYNOPSYS_UNCONNECTED_111, SYNOPSYS_UNCONNECTED_112,
         SYNOPSYS_UNCONNECTED_113, SYNOPSYS_UNCONNECTED_114,
         SYNOPSYS_UNCONNECTED_115, SYNOPSYS_UNCONNECTED_116,
         SYNOPSYS_UNCONNECTED_117, SYNOPSYS_UNCONNECTED_118,
         SYNOPSYS_UNCONNECTED_119, SYNOPSYS_UNCONNECTED_120,
         SYNOPSYS_UNCONNECTED_121, SYNOPSYS_UNCONNECTED_122,
         SYNOPSYS_UNCONNECTED_123, SYNOPSYS_UNCONNECTED_124,
         SYNOPSYS_UNCONNECTED_125, SYNOPSYS_UNCONNECTED_126,
         SYNOPSYS_UNCONNECTED_127, SYNOPSYS_UNCONNECTED_128,
         SYNOPSYS_UNCONNECTED_129, SYNOPSYS_UNCONNECTED_130,
         SYNOPSYS_UNCONNECTED_131, SYNOPSYS_UNCONNECTED_132,
         SYNOPSYS_UNCONNECTED_133, SYNOPSYS_UNCONNECTED_134,
         SYNOPSYS_UNCONNECTED_135, SYNOPSYS_UNCONNECTED_136,
         SYNOPSYS_UNCONNECTED_137, SYNOPSYS_UNCONNECTED_138,
         SYNOPSYS_UNCONNECTED_139, SYNOPSYS_UNCONNECTED_140,
         SYNOPSYS_UNCONNECTED_141, SYNOPSYS_UNCONNECTED_142,
         SYNOPSYS_UNCONNECTED_143, SYNOPSYS_UNCONNECTED_144,
         SYNOPSYS_UNCONNECTED_145, SYNOPSYS_UNCONNECTED_146,
         SYNOPSYS_UNCONNECTED_147, SYNOPSYS_UNCONNECTED_148,
         SYNOPSYS_UNCONNECTED_149, SYNOPSYS_UNCONNECTED_150,
         SYNOPSYS_UNCONNECTED_151, SYNOPSYS_UNCONNECTED_152,
         SYNOPSYS_UNCONNECTED_153, SYNOPSYS_UNCONNECTED_154,
         SYNOPSYS_UNCONNECTED_155, SYNOPSYS_UNCONNECTED_156,
         SYNOPSYS_UNCONNECTED_157, SYNOPSYS_UNCONNECTED_158,
         SYNOPSYS_UNCONNECTED_159, SYNOPSYS_UNCONNECTED_160,
         SYNOPSYS_UNCONNECTED_161, SYNOPSYS_UNCONNECTED_162,
         SYNOPSYS_UNCONNECTED_163, SYNOPSYS_UNCONNECTED_164,
         SYNOPSYS_UNCONNECTED_165, SYNOPSYS_UNCONNECTED_166,
         SYNOPSYS_UNCONNECTED_167, SYNOPSYS_UNCONNECTED_168,
         SYNOPSYS_UNCONNECTED_169, SYNOPSYS_UNCONNECTED_170,
         SYNOPSYS_UNCONNECTED_171, SYNOPSYS_UNCONNECTED_172,
         SYNOPSYS_UNCONNECTED_173, SYNOPSYS_UNCONNECTED_174,
         SYNOPSYS_UNCONNECTED_175, SYNOPSYS_UNCONNECTED_176,
         SYNOPSYS_UNCONNECTED_177, SYNOPSYS_UNCONNECTED_178,
         SYNOPSYS_UNCONNECTED_179, SYNOPSYS_UNCONNECTED_180,
         SYNOPSYS_UNCONNECTED_181, SYNOPSYS_UNCONNECTED_182,
         SYNOPSYS_UNCONNECTED_183, SYNOPSYS_UNCONNECTED_184,
         SYNOPSYS_UNCONNECTED_185, SYNOPSYS_UNCONNECTED_186,
         SYNOPSYS_UNCONNECTED_187, SYNOPSYS_UNCONNECTED_188,
         SYNOPSYS_UNCONNECTED_189, SYNOPSYS_UNCONNECTED_190,
         SYNOPSYS_UNCONNECTED_191, SYNOPSYS_UNCONNECTED_192,
         SYNOPSYS_UNCONNECTED_193, SYNOPSYS_UNCONNECTED_194,
         SYNOPSYS_UNCONNECTED_195, SYNOPSYS_UNCONNECTED_196,
         SYNOPSYS_UNCONNECTED_197, SYNOPSYS_UNCONNECTED_198,
         SYNOPSYS_UNCONNECTED_199, SYNOPSYS_UNCONNECTED_200,
         SYNOPSYS_UNCONNECTED_201, SYNOPSYS_UNCONNECTED_202,
         SYNOPSYS_UNCONNECTED_203, SYNOPSYS_UNCONNECTED_204,
         SYNOPSYS_UNCONNECTED_205, SYNOPSYS_UNCONNECTED_206,
         SYNOPSYS_UNCONNECTED_207, SYNOPSYS_UNCONNECTED_208,
         SYNOPSYS_UNCONNECTED_209, SYNOPSYS_UNCONNECTED_210,
         SYNOPSYS_UNCONNECTED_211, SYNOPSYS_UNCONNECTED_212,
         SYNOPSYS_UNCONNECTED_213, SYNOPSYS_UNCONNECTED_214,
         SYNOPSYS_UNCONNECTED_215, SYNOPSYS_UNCONNECTED_216,
         SYNOPSYS_UNCONNECTED_217, SYNOPSYS_UNCONNECTED_218,
         SYNOPSYS_UNCONNECTED_219, SYNOPSYS_UNCONNECTED_220,
         SYNOPSYS_UNCONNECTED_221, SYNOPSYS_UNCONNECTED_222,
         SYNOPSYS_UNCONNECTED_223, SYNOPSYS_UNCONNECTED_224,
         SYNOPSYS_UNCONNECTED_225, SYNOPSYS_UNCONNECTED_226,
         SYNOPSYS_UNCONNECTED_227, SYNOPSYS_UNCONNECTED_228,
         SYNOPSYS_UNCONNECTED_229, SYNOPSYS_UNCONNECTED_230,
         SYNOPSYS_UNCONNECTED_231, SYNOPSYS_UNCONNECTED_232,
         SYNOPSYS_UNCONNECTED_233, SYNOPSYS_UNCONNECTED_234,
         SYNOPSYS_UNCONNECTED_235, SYNOPSYS_UNCONNECTED_236,
         SYNOPSYS_UNCONNECTED_237, SYNOPSYS_UNCONNECTED_238,
         SYNOPSYS_UNCONNECTED_239, SYNOPSYS_UNCONNECTED_240,
         SYNOPSYS_UNCONNECTED_241, SYNOPSYS_UNCONNECTED_242,
         SYNOPSYS_UNCONNECTED_243, SYNOPSYS_UNCONNECTED_244,
         SYNOPSYS_UNCONNECTED_245, SYNOPSYS_UNCONNECTED_246,
         SYNOPSYS_UNCONNECTED_247, SYNOPSYS_UNCONNECTED_248,
         SYNOPSYS_UNCONNECTED_249, SYNOPSYS_UNCONNECTED_250,
         SYNOPSYS_UNCONNECTED_251, SYNOPSYS_UNCONNECTED_252,
         SYNOPSYS_UNCONNECTED_253, SYNOPSYS_UNCONNECTED_254,
         SYNOPSYS_UNCONNECTED_255, SYNOPSYS_UNCONNECTED_256,
         SYNOPSYS_UNCONNECTED_257, SYNOPSYS_UNCONNECTED_258,
         SYNOPSYS_UNCONNECTED_259, SYNOPSYS_UNCONNECTED_260,
         SYNOPSYS_UNCONNECTED_261, SYNOPSYS_UNCONNECTED_262,
         SYNOPSYS_UNCONNECTED_263, SYNOPSYS_UNCONNECTED_264,
         SYNOPSYS_UNCONNECTED_265, SYNOPSYS_UNCONNECTED_266,
         SYNOPSYS_UNCONNECTED_267, SYNOPSYS_UNCONNECTED_268,
         SYNOPSYS_UNCONNECTED_269, SYNOPSYS_UNCONNECTED_270,
         SYNOPSYS_UNCONNECTED_271, SYNOPSYS_UNCONNECTED_272,
         SYNOPSYS_UNCONNECTED_273, SYNOPSYS_UNCONNECTED_274,
         SYNOPSYS_UNCONNECTED_275, SYNOPSYS_UNCONNECTED_276,
         SYNOPSYS_UNCONNECTED_277, SYNOPSYS_UNCONNECTED_278,
         SYNOPSYS_UNCONNECTED_279, SYNOPSYS_UNCONNECTED_280,
         SYNOPSYS_UNCONNECTED_281, SYNOPSYS_UNCONNECTED_282,
         SYNOPSYS_UNCONNECTED_283, SYNOPSYS_UNCONNECTED_284,
         SYNOPSYS_UNCONNECTED_285, SYNOPSYS_UNCONNECTED_286,
         SYNOPSYS_UNCONNECTED_287, SYNOPSYS_UNCONNECTED_288,
         SYNOPSYS_UNCONNECTED_289, SYNOPSYS_UNCONNECTED_290,
         SYNOPSYS_UNCONNECTED_291, SYNOPSYS_UNCONNECTED_292,
         SYNOPSYS_UNCONNECTED_293, SYNOPSYS_UNCONNECTED_294,
         SYNOPSYS_UNCONNECTED_295, SYNOPSYS_UNCONNECTED_296,
         SYNOPSYS_UNCONNECTED_297, SYNOPSYS_UNCONNECTED_298,
         SYNOPSYS_UNCONNECTED_299, SYNOPSYS_UNCONNECTED_300,
         SYNOPSYS_UNCONNECTED_301, SYNOPSYS_UNCONNECTED_302,
         SYNOPSYS_UNCONNECTED_303, SYNOPSYS_UNCONNECTED_304,
         SYNOPSYS_UNCONNECTED_305, SYNOPSYS_UNCONNECTED_306,
         SYNOPSYS_UNCONNECTED_307, SYNOPSYS_UNCONNECTED_308,
         SYNOPSYS_UNCONNECTED_309, SYNOPSYS_UNCONNECTED_310,
         SYNOPSYS_UNCONNECTED_311, SYNOPSYS_UNCONNECTED_312,
         SYNOPSYS_UNCONNECTED_313, SYNOPSYS_UNCONNECTED_314,
         SYNOPSYS_UNCONNECTED_315, SYNOPSYS_UNCONNECTED_316,
         SYNOPSYS_UNCONNECTED_317, SYNOPSYS_UNCONNECTED_318,
         SYNOPSYS_UNCONNECTED_319, SYNOPSYS_UNCONNECTED_320,
         SYNOPSYS_UNCONNECTED_321, SYNOPSYS_UNCONNECTED_322,
         SYNOPSYS_UNCONNECTED_323, SYNOPSYS_UNCONNECTED_324,
         SYNOPSYS_UNCONNECTED_325, SYNOPSYS_UNCONNECTED_326,
         SYNOPSYS_UNCONNECTED_327, SYNOPSYS_UNCONNECTED_328,
         SYNOPSYS_UNCONNECTED_329, SYNOPSYS_UNCONNECTED_330,
         SYNOPSYS_UNCONNECTED_331, SYNOPSYS_UNCONNECTED_332,
         SYNOPSYS_UNCONNECTED_333, SYNOPSYS_UNCONNECTED_334,
         SYNOPSYS_UNCONNECTED_335, SYNOPSYS_UNCONNECTED_336,
         SYNOPSYS_UNCONNECTED_337, SYNOPSYS_UNCONNECTED_338,
         SYNOPSYS_UNCONNECTED_339, SYNOPSYS_UNCONNECTED_340,
         SYNOPSYS_UNCONNECTED_341, SYNOPSYS_UNCONNECTED_342,
         SYNOPSYS_UNCONNECTED_343, SYNOPSYS_UNCONNECTED_344,
         SYNOPSYS_UNCONNECTED_345, SYNOPSYS_UNCONNECTED_346,
         SYNOPSYS_UNCONNECTED_347, SYNOPSYS_UNCONNECTED_348,
         SYNOPSYS_UNCONNECTED_349, SYNOPSYS_UNCONNECTED_350,
         SYNOPSYS_UNCONNECTED_351, SYNOPSYS_UNCONNECTED_352,
         SYNOPSYS_UNCONNECTED_353, SYNOPSYS_UNCONNECTED_354,
         SYNOPSYS_UNCONNECTED_355, SYNOPSYS_UNCONNECTED_356,
         SYNOPSYS_UNCONNECTED_357, SYNOPSYS_UNCONNECTED_358,
         SYNOPSYS_UNCONNECTED_359, SYNOPSYS_UNCONNECTED_360,
         SYNOPSYS_UNCONNECTED_361, SYNOPSYS_UNCONNECTED_362,
         SYNOPSYS_UNCONNECTED_363, SYNOPSYS_UNCONNECTED_364,
         SYNOPSYS_UNCONNECTED_365, SYNOPSYS_UNCONNECTED_366,
         SYNOPSYS_UNCONNECTED_367, SYNOPSYS_UNCONNECTED_368,
         SYNOPSYS_UNCONNECTED_369, SYNOPSYS_UNCONNECTED_370,
         SYNOPSYS_UNCONNECTED_371, SYNOPSYS_UNCONNECTED_372,
         SYNOPSYS_UNCONNECTED_373, SYNOPSYS_UNCONNECTED_374,
         SYNOPSYS_UNCONNECTED_375, SYNOPSYS_UNCONNECTED_376,
         SYNOPSYS_UNCONNECTED_377, SYNOPSYS_UNCONNECTED_378,
         SYNOPSYS_UNCONNECTED_379, SYNOPSYS_UNCONNECTED_380,
         SYNOPSYS_UNCONNECTED_381, SYNOPSYS_UNCONNECTED_382,
         SYNOPSYS_UNCONNECTED_383, SYNOPSYS_UNCONNECTED_384,
         SYNOPSYS_UNCONNECTED_385, SYNOPSYS_UNCONNECTED_386,
         SYNOPSYS_UNCONNECTED_387, SYNOPSYS_UNCONNECTED_388,
         SYNOPSYS_UNCONNECTED_389, SYNOPSYS_UNCONNECTED_390,
         SYNOPSYS_UNCONNECTED_391, SYNOPSYS_UNCONNECTED_392,
         SYNOPSYS_UNCONNECTED_393, SYNOPSYS_UNCONNECTED_394,
         SYNOPSYS_UNCONNECTED_395, SYNOPSYS_UNCONNECTED_396,
         SYNOPSYS_UNCONNECTED_397, SYNOPSYS_UNCONNECTED_398,
         SYNOPSYS_UNCONNECTED_399, SYNOPSYS_UNCONNECTED_400,
         SYNOPSYS_UNCONNECTED_401, SYNOPSYS_UNCONNECTED_402,
         SYNOPSYS_UNCONNECTED_403, SYNOPSYS_UNCONNECTED_404,
         SYNOPSYS_UNCONNECTED_405, SYNOPSYS_UNCONNECTED_406,
         SYNOPSYS_UNCONNECTED_407, SYNOPSYS_UNCONNECTED_408,
         SYNOPSYS_UNCONNECTED_409, SYNOPSYS_UNCONNECTED_410,
         SYNOPSYS_UNCONNECTED_411, SYNOPSYS_UNCONNECTED_412;
  wire   [26:2] boothout1;
  wire   [26:0] boothout2;
  wire   [26:0] boothout3;
  wire   [26:0] boothout4;
  wire   [26:0] boothout5;
  wire   [26:0] boothout6;
  wire   [26:0] boothout7;
  wire   [26:0] boothout8;
  wire   [26:0] boothout9;
  wire   [26:0] boothout10;
  wire   [26:0] boothout11;
  wire   [25:0] boothout12;
  wire   [22:0] boothout13;
  wire   [29:2] cout1;
  wire   [31:3] mulout1;
  wire   [35:8] cout2;
  wire   [37:6] mulout2;
  wire   [41:14] cout3;
  wire   [42:12] mulout3;
  wire   [46:20] cout4;
  wire   [47:18] mulout4;
  wire   [31:3] cout5;
  wire   [46:4] mulout5;
  wire   [37:9] cout6;
  wire   [42:6] mulout6;
  wire   [46:18] cout7;
  wire   [47:12] mulout7;
  wire   [38:4] cout8;
  wire   [46:5] mulout8;
  wire   [46:12] cout9;
  wire   [47:6] mulout9;
  wire   [46:5] cout10;
  wire   [47:6] mulout10;
  wire   [46:6] cout11;
  wire   [47:7] mulout11;
  wire   [47:0] a;
  wire   [47:8] b;

  booth27_52 booth1 ( .out1({boothout1, SYNOPSYS_UNCONNECTED_1, 
        SYNOPSYS_UNCONNECTED_2}), .in1({in1[1:0], 1'b0}), .in2({1'b0, 1'b0, 
        1'b1, n34, n33, n32, n31, n30, n29, n28, n27, n26, n25, in2[12], n24, 
        in2[10], n23, in2[8], n21, in2[6], n20, in2[4], n19, in2[2], n18, n17}) );
  booth27_51 booth2 ( .out1(boothout2), .in1(in1[3:1]), .in2({1'b0, 1'b0, 1'b1, 
        n34, n33, n32, n31, n30, n29, n28, n27, n26, n25, in2[12], n24, 
        in2[10], n23, in2[8], n21, in2[6], n20, in2[4], n19, in2[2], n18, n17}) );
  booth27_50 booth3 ( .out1(boothout3), .in1(in1[5:3]), .in2({1'b0, 1'b0, 1'b1, 
        n34, n33, n32, n31, n30, n29, n28, n27, n26, n25, in2[12], n24, 
        in2[10], n23, in2[8], n21, in2[6], n20, in2[4], n19, in2[2], n18, n17}) );
  booth27_49 booth4 ( .out1(boothout4), .in1(in1[7:5]), .in2({1'b0, 1'b0, 1'b1, 
        n34, n33, n32, n31, n30, n29, n28, n27, n26, n25, in2[12], n24, 
        in2[10], n23, in2[8], n21, in2[6], n20, in2[4], n19, in2[2], n18, n17}) );
  booth27_48 booth5 ( .out1(boothout5), .in1(in1[9:7]), .in2({1'b0, 1'b0, 1'b1, 
        n34, n33, n32, n31, n30, n29, n28, n27, n26, n25, in2[12], n24, 
        in2[10], n23, in2[8], n21, in2[6], n20, in2[4], n19, in2[2], n18, n17}) );
  booth27_47 booth6 ( .out1(boothout6), .in1(in1[11:9]), .in2({1'b0, 1'b0, 
        1'b1, n34, n33, n32, n31, n30, n29, n28, n27, n26, n25, in2[12], n24, 
        in2[10], n23, in2[8], n21, in2[6], n20, in2[4], n19, in2[2], n18, n17}) );
  booth27_46 booth7 ( .out1(boothout7), .in1(in1[13:11]), .in2({1'b0, 1'b0, 
        1'b1, n34, n33, n32, n31, n30, n29, n28, n27, n26, n25, in2[12], n24, 
        in2[10], n23, in2[8], n21, in2[6], n20, in2[4], n19, in2[2], n18, n17}) );
  booth27_45 booth8 ( .out1(boothout8), .in1(in1[15:13]), .in2({1'b0, 1'b0, 
        1'b1, n34, n33, n32, n31, n30, n29, n28, n27, n26, n25, in2[12], n24, 
        in2[10], n23, in2[8], n21, in2[6], n20, in2[4], n19, in2[2], n18, n17}) );
  booth27_44 booth9 ( .out1(boothout9), .in1(in1[17:15]), .in2({1'b0, 1'b0, 
        1'b1, n34, n33, n32, n31, n30, n29, n28, n27, n26, n25, in2[12], n24, 
        in2[10], n23, in2[8], n21, in2[6], n20, in2[4], n19, in2[2], n18, n17}) );
  booth27_43 booth10 ( .out1(boothout10), .in1(in1[19:17]), .in2({1'b0, 1'b0, 
        1'b1, n34, n33, n32, n31, n30, n29, n28, n27, n26, n25, in2[12], n24, 
        in2[10], n23, in2[8], n21, in2[6], n20, in2[4], n19, in2[2], n18, n17}) );
  booth27_42 booth11 ( .out1(boothout11), .in1(in1[21:19]), .in2({1'b0, 1'b0, 
        1'b1, n34, n33, n32, n31, n30, n29, n28, n27, n26, n25, in2[12], n24, 
        in2[10], n23, in2[8], n21, in2[6], n20, in2[4], n19, in2[2], n18, n17}) );
  booth27_41 booth12 ( .out1({SYNOPSYS_UNCONNECTED_3, boothout12}), .in1({1'b1, 
        in1[22:21]}), .in2({1'b0, 1'b0, 1'b1, n34, n33, n32, n31, n30, n29, 
        n28, n27, n26, n25, in2[12], n24, in2[10], n23, in2[8], n21, in2[6], 
        n20, in2[4], n19, in2[2], n18, n17}) );
  booth27_40 booth13 ( .out1({SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, 
        SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, boothout13}), .in1({
        1'b0, 1'b0, 1'b1}), .in2({1'b0, 1'b0, 1'b1, n34, n33, n32, n31, n30, 
        n29, n28, n27, n26, n25, in2[12], n24, in2[10], n23, in2[8], n21, 
        in2[6], n20, in2[4], n19, in2[2], n18, n17}) );
  csa51squ_48 csa51squ1 ( .cout({SYNOPSYS_UNCONNECTED_8, 
        SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10, 
        SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12, 
        SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14, 
        SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16, 
        SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18, 
        SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20, 
        SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22, 
        SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24, 
        SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26, 
        SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28, cout1, 
        SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30}), .sumout({
        SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32, 
        SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34, 
        SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36, 
        SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38, 
        SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40, 
        SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42, 
        SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44, 
        SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46, 
        SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48, 
        SYNOPSYS_UNCONNECTED_49, mulout1[31], SYNOPSYS_UNCONNECTED_50, 
        mulout1[29:3], SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52, 
        SYNOPSYS_UNCONNECTED_53}), .in1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, boothout1, 1'b0, 1'b0}), .in2({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, boothout2, 
        1'b0, 1'b0}), .in3({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n132, 
        1'b0, boothout3[25:0], 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_47 csa51squ2 ( .cout({SYNOPSYS_UNCONNECTED_54, 
        SYNOPSYS_UNCONNECTED_55, SYNOPSYS_UNCONNECTED_56, 
        SYNOPSYS_UNCONNECTED_57, SYNOPSYS_UNCONNECTED_58, 
        SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_60, 
        SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_62, 
        SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_64, 
        SYNOPSYS_UNCONNECTED_65, SYNOPSYS_UNCONNECTED_66, 
        SYNOPSYS_UNCONNECTED_67, SYNOPSYS_UNCONNECTED_68, cout2, 
        SYNOPSYS_UNCONNECTED_69, SYNOPSYS_UNCONNECTED_70, 
        SYNOPSYS_UNCONNECTED_71, SYNOPSYS_UNCONNECTED_72, 
        SYNOPSYS_UNCONNECTED_73, SYNOPSYS_UNCONNECTED_74, 
        SYNOPSYS_UNCONNECTED_75, SYNOPSYS_UNCONNECTED_76}), .sumout({
        SYNOPSYS_UNCONNECTED_77, SYNOPSYS_UNCONNECTED_78, 
        SYNOPSYS_UNCONNECTED_79, SYNOPSYS_UNCONNECTED_80, 
        SYNOPSYS_UNCONNECTED_81, SYNOPSYS_UNCONNECTED_82, 
        SYNOPSYS_UNCONNECTED_83, SYNOPSYS_UNCONNECTED_84, 
        SYNOPSYS_UNCONNECTED_85, SYNOPSYS_UNCONNECTED_86, 
        SYNOPSYS_UNCONNECTED_87, SYNOPSYS_UNCONNECTED_88, 
        SYNOPSYS_UNCONNECTED_89, mulout2[37], SYNOPSYS_UNCONNECTED_90, 
        mulout2[35:6], SYNOPSYS_UNCONNECTED_91, SYNOPSYS_UNCONNECTED_92, 
        SYNOPSYS_UNCONNECTED_93, SYNOPSYS_UNCONNECTED_94, 
        SYNOPSYS_UNCONNECTED_95, SYNOPSYS_UNCONNECTED_96}), .in1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, boothout4, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, boothout5, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .in3({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n131, 1'b0, boothout6[25:0], 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_46 csa51squ3 ( .cout({SYNOPSYS_UNCONNECTED_97, 
        SYNOPSYS_UNCONNECTED_98, SYNOPSYS_UNCONNECTED_99, 
        SYNOPSYS_UNCONNECTED_100, SYNOPSYS_UNCONNECTED_101, 
        SYNOPSYS_UNCONNECTED_102, SYNOPSYS_UNCONNECTED_103, 
        SYNOPSYS_UNCONNECTED_104, SYNOPSYS_UNCONNECTED_105, cout3, 
        SYNOPSYS_UNCONNECTED_106, SYNOPSYS_UNCONNECTED_107, 
        SYNOPSYS_UNCONNECTED_108, SYNOPSYS_UNCONNECTED_109, 
        SYNOPSYS_UNCONNECTED_110, SYNOPSYS_UNCONNECTED_111, 
        SYNOPSYS_UNCONNECTED_112, SYNOPSYS_UNCONNECTED_113, 
        SYNOPSYS_UNCONNECTED_114, SYNOPSYS_UNCONNECTED_115, 
        SYNOPSYS_UNCONNECTED_116, SYNOPSYS_UNCONNECTED_117, 
        SYNOPSYS_UNCONNECTED_118, SYNOPSYS_UNCONNECTED_119}), .sumout({
        SYNOPSYS_UNCONNECTED_120, SYNOPSYS_UNCONNECTED_121, 
        SYNOPSYS_UNCONNECTED_122, SYNOPSYS_UNCONNECTED_123, 
        SYNOPSYS_UNCONNECTED_124, SYNOPSYS_UNCONNECTED_125, 
        SYNOPSYS_UNCONNECTED_126, SYNOPSYS_UNCONNECTED_127, mulout3, 
        SYNOPSYS_UNCONNECTED_128, SYNOPSYS_UNCONNECTED_129, 
        SYNOPSYS_UNCONNECTED_130, SYNOPSYS_UNCONNECTED_131, 
        SYNOPSYS_UNCONNECTED_132, SYNOPSYS_UNCONNECTED_133, 
        SYNOPSYS_UNCONNECTED_134, SYNOPSYS_UNCONNECTED_135, 
        SYNOPSYS_UNCONNECTED_136, SYNOPSYS_UNCONNECTED_137, 
        SYNOPSYS_UNCONNECTED_138, SYNOPSYS_UNCONNECTED_139}), .in1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, boothout7, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, boothout8, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .in3({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        boothout9, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_45 csa51squ4 ( .cout({SYNOPSYS_UNCONNECTED_140, 
        SYNOPSYS_UNCONNECTED_141, SYNOPSYS_UNCONNECTED_142, 
        SYNOPSYS_UNCONNECTED_143, cout4, SYNOPSYS_UNCONNECTED_144, 
        SYNOPSYS_UNCONNECTED_145, SYNOPSYS_UNCONNECTED_146, 
        SYNOPSYS_UNCONNECTED_147, SYNOPSYS_UNCONNECTED_148, 
        SYNOPSYS_UNCONNECTED_149, SYNOPSYS_UNCONNECTED_150, 
        SYNOPSYS_UNCONNECTED_151, SYNOPSYS_UNCONNECTED_152, 
        SYNOPSYS_UNCONNECTED_153, SYNOPSYS_UNCONNECTED_154, 
        SYNOPSYS_UNCONNECTED_155, SYNOPSYS_UNCONNECTED_156, 
        SYNOPSYS_UNCONNECTED_157, SYNOPSYS_UNCONNECTED_158, 
        SYNOPSYS_UNCONNECTED_159, SYNOPSYS_UNCONNECTED_160, 
        SYNOPSYS_UNCONNECTED_161, SYNOPSYS_UNCONNECTED_162, 
        SYNOPSYS_UNCONNECTED_163}), .sumout({SYNOPSYS_UNCONNECTED_164, 
        SYNOPSYS_UNCONNECTED_165, SYNOPSYS_UNCONNECTED_166, mulout4, 
        SYNOPSYS_UNCONNECTED_167, SYNOPSYS_UNCONNECTED_168, 
        SYNOPSYS_UNCONNECTED_169, SYNOPSYS_UNCONNECTED_170, 
        SYNOPSYS_UNCONNECTED_171, SYNOPSYS_UNCONNECTED_172, 
        SYNOPSYS_UNCONNECTED_173, SYNOPSYS_UNCONNECTED_174, 
        SYNOPSYS_UNCONNECTED_175, SYNOPSYS_UNCONNECTED_176, 
        SYNOPSYS_UNCONNECTED_177, SYNOPSYS_UNCONNECTED_178, 
        SYNOPSYS_UNCONNECTED_179, SYNOPSYS_UNCONNECTED_180, 
        SYNOPSYS_UNCONNECTED_181, SYNOPSYS_UNCONNECTED_182, 
        SYNOPSYS_UNCONNECTED_183, SYNOPSYS_UNCONNECTED_184}), .in1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, boothout10, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 1'b0, 1'b0, 1'b0, boothout11, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .in3({1'b0, 1'b0, 1'b0, boothout12, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_44 csa51squ5 ( .cout({SYNOPSYS_UNCONNECTED_185, 
        SYNOPSYS_UNCONNECTED_186, SYNOPSYS_UNCONNECTED_187, 
        SYNOPSYS_UNCONNECTED_188, SYNOPSYS_UNCONNECTED_189, 
        SYNOPSYS_UNCONNECTED_190, SYNOPSYS_UNCONNECTED_191, 
        SYNOPSYS_UNCONNECTED_192, SYNOPSYS_UNCONNECTED_193, 
        SYNOPSYS_UNCONNECTED_194, SYNOPSYS_UNCONNECTED_195, 
        SYNOPSYS_UNCONNECTED_196, SYNOPSYS_UNCONNECTED_197, 
        SYNOPSYS_UNCONNECTED_198, SYNOPSYS_UNCONNECTED_199, 
        SYNOPSYS_UNCONNECTED_200, SYNOPSYS_UNCONNECTED_201, 
        SYNOPSYS_UNCONNECTED_202, SYNOPSYS_UNCONNECTED_203, cout5, 
        SYNOPSYS_UNCONNECTED_204, SYNOPSYS_UNCONNECTED_205, 
        SYNOPSYS_UNCONNECTED_206}), .sumout({SYNOPSYS_UNCONNECTED_207, 
        SYNOPSYS_UNCONNECTED_208, SYNOPSYS_UNCONNECTED_209, 
        SYNOPSYS_UNCONNECTED_210, mulout5, SYNOPSYS_UNCONNECTED_211, 
        SYNOPSYS_UNCONNECTED_212, SYNOPSYS_UNCONNECTED_213, 
        SYNOPSYS_UNCONNECTED_214}), .in1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, cout1, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, mulout1[31], 1'b0, mulout1[29:3], 1'b0, 1'b0, 1'b0}), 
        .in3({1'b0, 1'b0, 1'b0, 1'b1, boothout13, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_43 csa51squ6 ( .cout({SYNOPSYS_UNCONNECTED_215, 
        SYNOPSYS_UNCONNECTED_216, SYNOPSYS_UNCONNECTED_217, 
        SYNOPSYS_UNCONNECTED_218, SYNOPSYS_UNCONNECTED_219, 
        SYNOPSYS_UNCONNECTED_220, SYNOPSYS_UNCONNECTED_221, 
        SYNOPSYS_UNCONNECTED_222, SYNOPSYS_UNCONNECTED_223, 
        SYNOPSYS_UNCONNECTED_224, SYNOPSYS_UNCONNECTED_225, 
        SYNOPSYS_UNCONNECTED_226, SYNOPSYS_UNCONNECTED_227, cout6, 
        SYNOPSYS_UNCONNECTED_228, SYNOPSYS_UNCONNECTED_229, 
        SYNOPSYS_UNCONNECTED_230, SYNOPSYS_UNCONNECTED_231, 
        SYNOPSYS_UNCONNECTED_232, SYNOPSYS_UNCONNECTED_233, 
        SYNOPSYS_UNCONNECTED_234, SYNOPSYS_UNCONNECTED_235, 
        SYNOPSYS_UNCONNECTED_236}), .sumout({SYNOPSYS_UNCONNECTED_237, 
        SYNOPSYS_UNCONNECTED_238, SYNOPSYS_UNCONNECTED_239, 
        SYNOPSYS_UNCONNECTED_240, SYNOPSYS_UNCONNECTED_241, 
        SYNOPSYS_UNCONNECTED_242, SYNOPSYS_UNCONNECTED_243, 
        SYNOPSYS_UNCONNECTED_244, mulout6, SYNOPSYS_UNCONNECTED_245, 
        SYNOPSYS_UNCONNECTED_246, SYNOPSYS_UNCONNECTED_247, 
        SYNOPSYS_UNCONNECTED_248, SYNOPSYS_UNCONNECTED_249, 
        SYNOPSYS_UNCONNECTED_250}), .in1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, cout2, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        mulout2[37], 1'b0, mulout2[35:6], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .in3({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, cout3, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  csa51squ_42 csa51squ7 ( .cout({SYNOPSYS_UNCONNECTED_251, 
        SYNOPSYS_UNCONNECTED_252, SYNOPSYS_UNCONNECTED_253, 
        SYNOPSYS_UNCONNECTED_254, cout7, SYNOPSYS_UNCONNECTED_255, 
        SYNOPSYS_UNCONNECTED_256, SYNOPSYS_UNCONNECTED_257, 
        SYNOPSYS_UNCONNECTED_258, SYNOPSYS_UNCONNECTED_259, 
        SYNOPSYS_UNCONNECTED_260, SYNOPSYS_UNCONNECTED_261, 
        SYNOPSYS_UNCONNECTED_262, SYNOPSYS_UNCONNECTED_263, 
        SYNOPSYS_UNCONNECTED_264, SYNOPSYS_UNCONNECTED_265, 
        SYNOPSYS_UNCONNECTED_266, SYNOPSYS_UNCONNECTED_267, 
        SYNOPSYS_UNCONNECTED_268, SYNOPSYS_UNCONNECTED_269, 
        SYNOPSYS_UNCONNECTED_270, SYNOPSYS_UNCONNECTED_271, 
        SYNOPSYS_UNCONNECTED_272}), .sumout({SYNOPSYS_UNCONNECTED_273, 
        SYNOPSYS_UNCONNECTED_274, SYNOPSYS_UNCONNECTED_275, mulout7, 
        SYNOPSYS_UNCONNECTED_276, SYNOPSYS_UNCONNECTED_277, 
        SYNOPSYS_UNCONNECTED_278, SYNOPSYS_UNCONNECTED_279, 
        SYNOPSYS_UNCONNECTED_280, SYNOPSYS_UNCONNECTED_281, 
        SYNOPSYS_UNCONNECTED_282, SYNOPSYS_UNCONNECTED_283, 
        SYNOPSYS_UNCONNECTED_284, SYNOPSYS_UNCONNECTED_285, 
        SYNOPSYS_UNCONNECTED_286, SYNOPSYS_UNCONNECTED_287}), .in1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mulout3, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 1'b0, 
        1'b0, cout4, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in3({1'b0, 1'b0, 1'b0, mulout4, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_41 csa51squ8 ( .cout({SYNOPSYS_UNCONNECTED_288, 
        SYNOPSYS_UNCONNECTED_289, SYNOPSYS_UNCONNECTED_290, 
        SYNOPSYS_UNCONNECTED_291, SYNOPSYS_UNCONNECTED_292, 
        SYNOPSYS_UNCONNECTED_293, SYNOPSYS_UNCONNECTED_294, 
        SYNOPSYS_UNCONNECTED_295, SYNOPSYS_UNCONNECTED_296, 
        SYNOPSYS_UNCONNECTED_297, SYNOPSYS_UNCONNECTED_298, 
        SYNOPSYS_UNCONNECTED_299, cout8, SYNOPSYS_UNCONNECTED_300, 
        SYNOPSYS_UNCONNECTED_301, SYNOPSYS_UNCONNECTED_302, 
        SYNOPSYS_UNCONNECTED_303}), .sumout({SYNOPSYS_UNCONNECTED_304, 
        SYNOPSYS_UNCONNECTED_305, SYNOPSYS_UNCONNECTED_306, 
        SYNOPSYS_UNCONNECTED_307, mulout8, SYNOPSYS_UNCONNECTED_308, 
        SYNOPSYS_UNCONNECTED_309, SYNOPSYS_UNCONNECTED_310, 
        SYNOPSYS_UNCONNECTED_311, SYNOPSYS_UNCONNECTED_312}), .in1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, cout5, 1'b0, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 
        1'b0, 1'b0, 1'b1, mulout5, 1'b0, 1'b0, 1'b0, 1'b0}), .in3({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, cout6, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_40 csa51squ9 ( .cout({SYNOPSYS_UNCONNECTED_313, 
        SYNOPSYS_UNCONNECTED_314, SYNOPSYS_UNCONNECTED_315, 
        SYNOPSYS_UNCONNECTED_316, cout9, SYNOPSYS_UNCONNECTED_317, 
        SYNOPSYS_UNCONNECTED_318, SYNOPSYS_UNCONNECTED_319, 
        SYNOPSYS_UNCONNECTED_320, SYNOPSYS_UNCONNECTED_321, 
        SYNOPSYS_UNCONNECTED_322, SYNOPSYS_UNCONNECTED_323, 
        SYNOPSYS_UNCONNECTED_324, SYNOPSYS_UNCONNECTED_325, 
        SYNOPSYS_UNCONNECTED_326, SYNOPSYS_UNCONNECTED_327, 
        SYNOPSYS_UNCONNECTED_328}), .sumout({SYNOPSYS_UNCONNECTED_329, 
        SYNOPSYS_UNCONNECTED_330, SYNOPSYS_UNCONNECTED_331, mulout9, 
        SYNOPSYS_UNCONNECTED_332, SYNOPSYS_UNCONNECTED_333, 
        SYNOPSYS_UNCONNECTED_334, SYNOPSYS_UNCONNECTED_335, 
        SYNOPSYS_UNCONNECTED_336, SYNOPSYS_UNCONNECTED_337}), .in1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mulout6, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .in2({1'b0, 1'b0, 1'b0, cout7, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .in3({1'b0, 1'b0, 1'b0, mulout7, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_39 csa51squ10 ( .cout({SYNOPSYS_UNCONNECTED_338, 
        SYNOPSYS_UNCONNECTED_339, SYNOPSYS_UNCONNECTED_340, 
        SYNOPSYS_UNCONNECTED_341, cout10, SYNOPSYS_UNCONNECTED_342, 
        SYNOPSYS_UNCONNECTED_343, SYNOPSYS_UNCONNECTED_344, 
        SYNOPSYS_UNCONNECTED_345, SYNOPSYS_UNCONNECTED_346}), .sumout({
        SYNOPSYS_UNCONNECTED_347, SYNOPSYS_UNCONNECTED_348, 
        SYNOPSYS_UNCONNECTED_349, mulout10, SYNOPSYS_UNCONNECTED_350, 
        SYNOPSYS_UNCONNECTED_351, SYNOPSYS_UNCONNECTED_352, 
        SYNOPSYS_UNCONNECTED_353, SYNOPSYS_UNCONNECTED_354, 
        SYNOPSYS_UNCONNECTED_355}), .in1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, cout8, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .in2({1'b0, 1'b0, 1'b0, 1'b1, mulout8, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .in3({1'b0, 1'b0, 1'b0, cout9, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_38 csa51squ11 ( .cout({SYNOPSYS_UNCONNECTED_356, 
        SYNOPSYS_UNCONNECTED_357, SYNOPSYS_UNCONNECTED_358, 
        SYNOPSYS_UNCONNECTED_359, cout11, SYNOPSYS_UNCONNECTED_360, 
        SYNOPSYS_UNCONNECTED_361, SYNOPSYS_UNCONNECTED_362, 
        SYNOPSYS_UNCONNECTED_363, SYNOPSYS_UNCONNECTED_364, 
        SYNOPSYS_UNCONNECTED_365}), .sumout({SYNOPSYS_UNCONNECTED_366, 
        SYNOPSYS_UNCONNECTED_367, SYNOPSYS_UNCONNECTED_368, mulout11, 
        SYNOPSYS_UNCONNECTED_369, SYNOPSYS_UNCONNECTED_370, 
        SYNOPSYS_UNCONNECTED_371, SYNOPSYS_UNCONNECTED_372, 
        SYNOPSYS_UNCONNECTED_373, SYNOPSYS_UNCONNECTED_374, 
        SYNOPSYS_UNCONNECTED_375}), .in1({1'b0, 1'b0, 1'b0, mulout9, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 1'b0, 1'b0, cout10, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in3({1'b0, 1'b0, 1'b0, mulout10, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_37 csa51squ12 ( .sumout({SYNOPSYS_UNCONNECTED_376, 
        SYNOPSYS_UNCONNECTED_377, SYNOPSYS_UNCONNECTED_378, N101, N100, N99, 
        N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, 
        N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, 
        N70, N69, N68, N67, N66, N65, N64, N63, N62, SYNOPSYS_UNCONNECTED_379, 
        SYNOPSYS_UNCONNECTED_380, SYNOPSYS_UNCONNECTED_381, 
        SYNOPSYS_UNCONNECTED_382, SYNOPSYS_UNCONNECTED_383, 
        SYNOPSYS_UNCONNECTED_384, SYNOPSYS_UNCONNECTED_385, 
        SYNOPSYS_UNCONNECTED_386}), .in1({1'b0, 1'b0, 1'b0, mulout11, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 1'b0, 1'b0, cout11, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in3({1'b1, 1'b0, 1'b1, 
        1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 
        1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .cout_46_(N50), .cout_44_(N48), .cout_42_(N46), .cout_40_(N44), .cout_38_(
        N42), .cout_36_(N40), .cout_34_(N38), .cout_32_(N36), .cout_30_(N34), 
        .cout_28_(N32), .cout_27_(N31), .cout_7__BAR(N11), .cout_8__BAR(N12), 
        .cout_9__BAR(N13), .cout_10__BAR(N14), .cout_11__BAR(N15), 
        .cout_12__BAR(N16), .cout_13__BAR(N17), .cout_14__BAR(N18), 
        .cout_15__BAR(N19), .cout_16__BAR(N20), .cout_17__BAR(N21), 
        .cout_18__BAR(N22), .cout_19__BAR(N23), .cout_20__BAR(N24), 
        .cout_21__BAR(N25), .cout_22__BAR(N26), .cout_23__BAR(N27), 
        .cout_24__BAR(N28), .cout_25__BAR(N29), .cout_26__BAR(N30), 
        .cout_29__BAR(N33), .cout_31__BAR(N35), .cout_33__BAR(N37), 
        .cout_35__BAR(N39), .cout_37__BAR(N41), .cout_39__BAR(N43), 
        .cout_41__BAR(N45), .cout_43__BAR(N47), .cout_45__BAR(N49) );
  cla51squ_4 cla51squ ( .out({SYNOPSYS_UNCONNECTED_387, 
        SYNOPSYS_UNCONNECTED_388, SYNOPSYS_UNCONNECTED_389, mulout[47:23], 
        SYNOPSYS_UNCONNECTED_390, SYNOPSYS_UNCONNECTED_391, 
        SYNOPSYS_UNCONNECTED_392, SYNOPSYS_UNCONNECTED_393, 
        SYNOPSYS_UNCONNECTED_394, SYNOPSYS_UNCONNECTED_395, 
        SYNOPSYS_UNCONNECTED_396, SYNOPSYS_UNCONNECTED_397, 
        SYNOPSYS_UNCONNECTED_398, SYNOPSYS_UNCONNECTED_399, 
        SYNOPSYS_UNCONNECTED_400, SYNOPSYS_UNCONNECTED_401, 
        SYNOPSYS_UNCONNECTED_402, SYNOPSYS_UNCONNECTED_403, 
        SYNOPSYS_UNCONNECTED_404, SYNOPSYS_UNCONNECTED_405, 
        SYNOPSYS_UNCONNECTED_406, SYNOPSYS_UNCONNECTED_407, 
        SYNOPSYS_UNCONNECTED_408, SYNOPSYS_UNCONNECTED_409, 
        SYNOPSYS_UNCONNECTED_410, SYNOPSYS_UNCONNECTED_411, 
        SYNOPSYS_UNCONNECTED_412}), .a({1'b0, 1'b0, 1'b0, a[47:8], 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({1'b0, 1'b0, 1'b0, b, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  DFFARX1 b_reg_47_ ( .D(N101), .CLK(clk), .RSTB(rst_n), .Q(b[47]) );
  DFFARX1 b_reg_46_ ( .D(N100), .CLK(clk), .RSTB(rst_n), .Q(b[46]) );
  DFFARX1 b_reg_45_ ( .D(N99), .CLK(clk), .RSTB(rst_n), .Q(b[45]) );
  DFFARX1 b_reg_44_ ( .D(N98), .CLK(clk), .RSTB(rst_n), .Q(b[44]) );
  DFFARX1 b_reg_43_ ( .D(N97), .CLK(clk), .RSTB(rst_n), .Q(b[43]) );
  DFFARX1 b_reg_42_ ( .D(N96), .CLK(clk), .RSTB(rst_n), .Q(b[42]) );
  DFFARX1 b_reg_41_ ( .D(N95), .CLK(clk), .RSTB(rst_n), .Q(b[41]) );
  DFFARX1 b_reg_40_ ( .D(N94), .CLK(clk), .RSTB(rst_n), .Q(b[40]) );
  DFFARX1 b_reg_39_ ( .D(N93), .CLK(clk), .RSTB(rst_n), .Q(b[39]) );
  DFFARX1 b_reg_38_ ( .D(N92), .CLK(clk), .RSTB(rst_n), .Q(b[38]) );
  DFFARX1 b_reg_37_ ( .D(N91), .CLK(clk), .RSTB(rst_n), .Q(b[37]) );
  DFFARX1 b_reg_36_ ( .D(N90), .CLK(clk), .RSTB(rst_n), .Q(b[36]) );
  DFFARX1 b_reg_35_ ( .D(N89), .CLK(clk), .RSTB(rst_n), .Q(b[35]) );
  DFFARX1 b_reg_34_ ( .D(N88), .CLK(clk), .RSTB(rst_n), .Q(b[34]) );
  DFFARX1 b_reg_33_ ( .D(N87), .CLK(clk), .RSTB(rst_n), .Q(b[33]) );
  DFFARX1 b_reg_32_ ( .D(N86), .CLK(clk), .RSTB(rst_n), .Q(b[32]) );
  DFFARX1 b_reg_31_ ( .D(N85), .CLK(clk), .RSTB(rst_n), .Q(b[31]) );
  DFFARX1 b_reg_30_ ( .D(N84), .CLK(clk), .RSTB(rst_n), .Q(b[30]) );
  DFFARX1 b_reg_29_ ( .D(N83), .CLK(clk), .RSTB(rst_n), .Q(b[29]) );
  DFFARX1 b_reg_28_ ( .D(N82), .CLK(clk), .RSTB(rst_n), .Q(b[28]) );
  DFFARX1 b_reg_27_ ( .D(N81), .CLK(clk), .RSTB(rst_n), .Q(b[27]) );
  DFFARX1 b_reg_26_ ( .D(N80), .CLK(clk), .RSTB(rst_n), .Q(b[26]) );
  DFFARX1 b_reg_25_ ( .D(N79), .CLK(clk), .RSTB(rst_n), .Q(b[25]) );
  DFFARX1 b_reg_24_ ( .D(N78), .CLK(clk), .RSTB(rst_n), .Q(b[24]) );
  DFFARX1 b_reg_23_ ( .D(N77), .CLK(clk), .RSTB(rst_n), .Q(b[23]) );
  DFFARX1 b_reg_22_ ( .D(N76), .CLK(clk), .RSTB(rst_n), .Q(b[22]) );
  DFFARX1 b_reg_21_ ( .D(N75), .CLK(clk), .RSTB(rst_n), .Q(b[21]) );
  DFFARX1 b_reg_20_ ( .D(N74), .CLK(clk), .RSTB(rst_n), .Q(b[20]) );
  DFFARX1 b_reg_19_ ( .D(N73), .CLK(clk), .RSTB(rst_n), .Q(b[19]) );
  DFFARX1 b_reg_18_ ( .D(N72), .CLK(clk), .RSTB(rst_n), .Q(b[18]) );
  DFFARX1 b_reg_17_ ( .D(N71), .CLK(clk), .RSTB(rst_n), .Q(b[17]) );
  DFFARX1 b_reg_16_ ( .D(N70), .CLK(clk), .RSTB(rst_n), .Q(b[16]) );
  DFFARX1 b_reg_15_ ( .D(N69), .CLK(clk), .RSTB(rst_n), .Q(b[15]) );
  DFFARX1 b_reg_14_ ( .D(N68), .CLK(clk), .RSTB(rst_n), .Q(b[14]) );
  DFFARX1 b_reg_13_ ( .D(N67), .CLK(clk), .RSTB(rst_n), .Q(b[13]) );
  DFFARX1 b_reg_12_ ( .D(N66), .CLK(clk), .RSTB(rst_n), .Q(b[12]) );
  DFFARX1 b_reg_11_ ( .D(N65), .CLK(clk), .RSTB(rst_n), .Q(b[11]) );
  DFFARX1 b_reg_10_ ( .D(N64), .CLK(clk), .RSTB(rst_n), .Q(b[10]) );
  DFFARX1 b_reg_9_ ( .D(N63), .CLK(clk), .RSTB(rst_n), .Q(b[9]) );
  DFFARX1 b_reg_8_ ( .D(N62), .CLK(clk), .RSTB(rst_n), .Q(b[8]) );
  DFFARX1 a_reg_47_ ( .D(N50), .CLK(clk), .RSTB(rst_n), .Q(a[47]) );
  DFFARX1 a_reg_46_ ( .D(n63), .CLK(clk), .RSTB(rst_n), .Q(a[46]) );
  DFFARX1 a_reg_45_ ( .D(N48), .CLK(clk), .RSTB(rst_n), .Q(a[45]) );
  DFFARX1 a_reg_44_ ( .D(n64), .CLK(clk), .RSTB(rst_n), .Q(a[44]) );
  DFFARX1 a_reg_43_ ( .D(N46), .CLK(clk), .RSTB(rst_n), .Q(a[43]) );
  DFFARX1 a_reg_42_ ( .D(n65), .CLK(clk), .RSTB(rst_n), .Q(a[42]) );
  DFFARX1 a_reg_41_ ( .D(N44), .CLK(clk), .RSTB(rst_n), .Q(a[41]) );
  DFFARX1 a_reg_40_ ( .D(n66), .CLK(clk), .RSTB(rst_n), .Q(a[40]) );
  DFFARX1 a_reg_39_ ( .D(N42), .CLK(clk), .RSTB(rst_n), .Q(a[39]) );
  DFFARX1 a_reg_38_ ( .D(n67), .CLK(clk), .RSTB(rst_n), .Q(a[38]) );
  DFFARX1 a_reg_37_ ( .D(N40), .CLK(clk), .RSTB(rst_n), .Q(a[37]) );
  DFFARX1 a_reg_36_ ( .D(n68), .CLK(clk), .RSTB(rst_n), .Q(a[36]) );
  DFFARX1 a_reg_35_ ( .D(N38), .CLK(clk), .RSTB(rst_n), .Q(a[35]) );
  DFFARX1 a_reg_34_ ( .D(n69), .CLK(clk), .RSTB(rst_n), .Q(a[34]) );
  DFFARX1 a_reg_33_ ( .D(N36), .CLK(clk), .RSTB(rst_n), .Q(a[33]) );
  DFFARX1 a_reg_32_ ( .D(n70), .CLK(clk), .RSTB(rst_n), .Q(a[32]) );
  DFFARX1 a_reg_31_ ( .D(N34), .CLK(clk), .RSTB(rst_n), .Q(a[31]) );
  DFFARX1 a_reg_30_ ( .D(n71), .CLK(clk), .RSTB(rst_n), .Q(a[30]) );
  DFFARX1 a_reg_29_ ( .D(N32), .CLK(clk), .RSTB(rst_n), .Q(a[29]) );
  DFFARX1 a_reg_28_ ( .D(N31), .CLK(clk), .RSTB(rst_n), .Q(a[28]) );
  DFFARX1 a_reg_27_ ( .D(n72), .CLK(clk), .RSTB(rst_n), .Q(a[27]) );
  DFFARX1 a_reg_26_ ( .D(n73), .CLK(clk), .RSTB(rst_n), .Q(a[26]) );
  DFFARX1 a_reg_25_ ( .D(n74), .CLK(clk), .RSTB(rst_n), .Q(a[25]) );
  DFFARX1 a_reg_24_ ( .D(n75), .CLK(clk), .RSTB(rst_n), .Q(a[24]) );
  DFFARX1 a_reg_23_ ( .D(n76), .CLK(clk), .RSTB(rst_n), .Q(a[23]) );
  DFFARX1 a_reg_22_ ( .D(n77), .CLK(clk), .RSTB(rst_n), .Q(a[22]) );
  DFFARX1 a_reg_21_ ( .D(n78), .CLK(clk), .RSTB(rst_n), .Q(a[21]) );
  DFFARX1 a_reg_20_ ( .D(n79), .CLK(clk), .RSTB(rst_n), .Q(a[20]) );
  DFFARX1 a_reg_19_ ( .D(n80), .CLK(clk), .RSTB(rst_n), .Q(a[19]) );
  DFFARX1 a_reg_18_ ( .D(n81), .CLK(clk), .RSTB(rst_n), .Q(a[18]) );
  DFFARX1 a_reg_17_ ( .D(n82), .CLK(clk), .RSTB(rst_n), .Q(a[17]) );
  DFFARX1 a_reg_16_ ( .D(n83), .CLK(clk), .RSTB(rst_n), .Q(a[16]) );
  DFFARX1 a_reg_15_ ( .D(n84), .CLK(clk), .RSTB(rst_n), .Q(a[15]) );
  DFFARX1 a_reg_14_ ( .D(n85), .CLK(clk), .RSTB(rst_n), .Q(a[14]) );
  DFFARX1 a_reg_13_ ( .D(n86), .CLK(clk), .RSTB(rst_n), .Q(a[13]) );
  DFFARX1 a_reg_12_ ( .D(n87), .CLK(clk), .RSTB(rst_n), .Q(a[12]) );
  DFFARX1 a_reg_11_ ( .D(n88), .CLK(clk), .RSTB(rst_n), .Q(a[11]) );
  DFFARX1 a_reg_10_ ( .D(n89), .CLK(clk), .RSTB(rst_n), .Q(a[10]) );
  DFFARX1 a_reg_9_ ( .D(n90), .CLK(clk), .RSTB(rst_n), .Q(a[9]) );
  DFFARX1 a_reg_8_ ( .D(n91), .CLK(clk), .RSTB(rst_n), .Q(a[8]) );
  INVX0 U5 ( .INP(boothout3[26]), .ZN(n132) );
  INVX0 U8 ( .INP(boothout6[26]), .ZN(n131) );
  NBUFFX8 U3 ( .INP(in2[18]), .Z(n30) );
  NBUFFX8 U4 ( .INP(in2[16]), .Z(n28) );
  NBUFFX8 U6 ( .INP(in2[14]), .Z(n26) );
  NBUFFX8 U7 ( .INP(in2[20]), .Z(n32) );
  NBUFFX8 U9 ( .INP(in2[19]), .Z(n31) );
  NBUFFX8 U10 ( .INP(in2[15]), .Z(n27) );
  NBUFFX8 U11 ( .INP(in2[17]), .Z(n29) );
  NBUFFX8 U12 ( .INP(in2[13]), .Z(n25) );
  NBUFFX8 U13 ( .INP(in2[21]), .Z(n33) );
  NBUFFX8 U14 ( .INP(in2[22]), .Z(n34) );
  NBUFFX8 U15 ( .INP(in2[3]), .Z(n19) );
  NBUFFX8 U16 ( .INP(in2[5]), .Z(n20) );
  NBUFFX8 U17 ( .INP(in2[9]), .Z(n23) );
  NBUFFX8 U18 ( .INP(in2[11]), .Z(n24) );
  INVX0 U19 ( .INP(n22), .ZN(n21) );
  NBUFFX8 U20 ( .INP(in2[1]), .Z(n18) );
  NBUFFX8 U21 ( .INP(in2[0]), .Z(n17) );
  INVX0 U36 ( .INP(in2[7]), .ZN(n22) );
  INVX0 U72 ( .INP(N49), .ZN(n63) );
  INVX0 U73 ( .INP(N47), .ZN(n64) );
  INVX0 U74 ( .INP(N45), .ZN(n65) );
  INVX0 U75 ( .INP(N43), .ZN(n66) );
  INVX0 U76 ( .INP(N41), .ZN(n67) );
  INVX0 U77 ( .INP(N39), .ZN(n68) );
  INVX0 U78 ( .INP(N37), .ZN(n69) );
  INVX0 U79 ( .INP(N35), .ZN(n70) );
  INVX0 U80 ( .INP(N33), .ZN(n71) );
  INVX0 U81 ( .INP(N30), .ZN(n72) );
  INVX0 U82 ( .INP(N29), .ZN(n73) );
  INVX0 U83 ( .INP(N28), .ZN(n74) );
  INVX0 U84 ( .INP(N27), .ZN(n75) );
  INVX0 U85 ( .INP(N26), .ZN(n76) );
  INVX0 U86 ( .INP(N25), .ZN(n77) );
  INVX0 U87 ( .INP(N24), .ZN(n78) );
  INVX0 U88 ( .INP(N23), .ZN(n79) );
  INVX0 U89 ( .INP(N22), .ZN(n80) );
  INVX0 U90 ( .INP(N21), .ZN(n81) );
  INVX0 U91 ( .INP(N20), .ZN(n82) );
  INVX0 U92 ( .INP(N19), .ZN(n83) );
  INVX0 U93 ( .INP(N18), .ZN(n84) );
  INVX0 U94 ( .INP(N17), .ZN(n85) );
  INVX0 U95 ( .INP(N16), .ZN(n86) );
  INVX0 U96 ( .INP(N15), .ZN(n87) );
  INVX0 U97 ( .INP(N14), .ZN(n88) );
  INVX0 U98 ( .INP(N13), .ZN(n89) );
  INVX0 U99 ( .INP(N12), .ZN(n90) );
  INVX0 U100 ( .INP(N11), .ZN(n91) );
endmodule


module add_433 ( s, a, b, co, ci_BAR );
  input a, b, ci_BAR;
  output s, co;


  XOR2X1 U1 ( .IN1(a), .IN2(ci_BAR), .Q(s) );
endmodule


module add_434 ( s, a, b, ci, co_BAR );
  input a, b, ci;
  output s, co_BAR;


  NAND2X0 U1 ( .IN1(ci), .IN2(a), .QN(co_BAR) );
  OA21X1 U2 ( .IN1(ci), .IN2(a), .IN3(co_BAR), .Q(s) );
endmodule


module add_435 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_436 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_437 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_438 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_439 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  INVX0 U1 ( .INP(a), .ZN(s) );
  NBUFFX2 U2 ( .INP(a), .Z(co) );
endmodule


module add_440 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  NBUFFX2 U1 ( .INP(a), .Z(s) );
endmodule


module adder8_31 ( out, a, b, cin );
  output [7:0] out;
  input [7:0] a;
  input [7:0] b;
  input cin;

  wire   [6:1] c;

  add_440 add_01 ( .s(out[0]), .a(a[0]), .b(1'b1), .ci(1'b1) );
  add_439 add_02 ( .s(out[1]), .a(a[1]), .b(1'b0), .ci(1'b1), .co(c[1]) );
  add_438 add_03 ( .s(out[2]), .a(a[2]), .b(1'b0), .ci(c[1]), .co(c[2]) );
  add_437 add_04 ( .s(out[3]), .a(a[3]), .b(1'b0), .ci(c[2]), .co(c[3]) );
  add_436 add_05 ( .s(out[4]), .a(a[4]), .b(1'b0), .ci(c[3]), .co(c[4]) );
  add_435 add_06 ( .s(out[5]), .a(a[5]), .b(1'b0), .ci(c[4]), .co(c[5]) );
  add_434 add_07 ( .s(out[6]), .a(a[6]), .b(1'b0), .ci(c[5]), .co_BAR(c[6]) );
  add_433 add_08 ( .s(out[7]), .a(a[7]), .b(1'b1), .ci_BAR(c[6]) );
endmodule


module add_441 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  XOR3X1 U1 ( .IN1(b), .IN2(ci), .IN3(a), .Q(s) );
endmodule


module add_442 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_443 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_444 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_445 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_446 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_447 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_448 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(b), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(b), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module adder8_32 ( out, a, b, cin );
  output [7:0] out;
  input [7:0] a;
  input [7:0] b;
  input cin;

  wire   [6:0] c;

  add_448 add_01 ( .s(out[0]), .a(a[0]), .b(b[0]), .ci(1'b0), .co(c[0]) );
  add_447 add_02 ( .s(out[1]), .a(a[1]), .b(b[1]), .ci(c[0]), .co(c[1]) );
  add_446 add_03 ( .s(out[2]), .a(a[2]), .b(b[2]), .ci(c[1]), .co(c[2]) );
  add_445 add_04 ( .s(out[3]), .a(a[3]), .b(b[3]), .ci(c[2]), .co(c[3]) );
  add_444 add_05 ( .s(out[4]), .a(a[4]), .b(b[4]), .ci(c[3]), .co(c[4]) );
  add_443 add_06 ( .s(out[5]), .a(a[5]), .b(b[5]), .ci(c[4]), .co(c[5]) );
  add_442 add_07 ( .s(out[6]), .a(a[6]), .b(b[6]), .ci(c[5]), .co(c[6]) );
  add_441 add_08 ( .s(out[7]), .a(a[7]), .b(b[7]), .ci(c[6]) );
endmodule


module floating_point_multiple_4 ( clk, rst_n, input_factor_01, 
        input_factor_02, output_multiply );
  input [31:0] input_factor_01;
  input [31:0] input_factor_02;
  output [31:0] output_multiply;
  input clk, rst_n;
  wire   N5, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22,
         N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N48, N49, N50, N51,
         N52, N53, N54, N55, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22,
         SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24,
         SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26;
  wire   [47:23] base_multiply_result;
  wire   [47:23] mulout;
  wire   [7:0] exponent_factor_12;
  wire   [7:0] pre_mul_output_exponent;

  mul26_4 mul26_01 ( .clk(clk), .rst_n(rst_n), .in1({1'b0, 1'b0, 1'b1, 
        input_factor_01[22:0]}), .in2({1'b0, 1'b0, 1'b1, input_factor_02[22:0]}), .en(1'b1), .mulout({SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, 
        SYNOPSYS_UNCONNECTED_3, mulout, SYNOPSYS_UNCONNECTED_4, 
        SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, 
        SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, 
        SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11, 
        SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13, 
        SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, 
        SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17, 
        SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19, 
        SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21, 
        SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_23, 
        SYNOPSYS_UNCONNECTED_24, SYNOPSYS_UNCONNECTED_25, 
        SYNOPSYS_UNCONNECTED_26}) );
  adder8_32 adder8_01 ( .out(exponent_factor_12), .a(input_factor_01[30:23]), 
        .b(input_factor_02[30:23]), .cin(1'b0) );
  adder8_31 adder8_02 ( .out(pre_mul_output_exponent), .a(exponent_factor_12), 
        .b({1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0}), .cin(1'b1) );
  DFFARX1 mul_output_sign_reg ( .D(N5), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[31]) );
  DFFARX1 base_multiply_result_reg_47_ ( .D(mulout[47]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[47]) );
  DFFARX1 base_multiply_result_reg_46_ ( .D(mulout[46]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[46]) );
  DFFARX1 base_multiply_result_reg_45_ ( .D(mulout[45]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[45]) );
  DFFARX1 base_multiply_result_reg_44_ ( .D(mulout[44]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[44]) );
  DFFARX1 base_multiply_result_reg_43_ ( .D(mulout[43]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[43]) );
  DFFARX1 base_multiply_result_reg_42_ ( .D(mulout[42]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[42]) );
  DFFARX1 base_multiply_result_reg_41_ ( .D(mulout[41]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[41]) );
  DFFARX1 base_multiply_result_reg_40_ ( .D(mulout[40]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[40]) );
  DFFARX1 base_multiply_result_reg_39_ ( .D(mulout[39]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[39]) );
  DFFARX1 base_multiply_result_reg_38_ ( .D(mulout[38]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[38]) );
  DFFARX1 base_multiply_result_reg_37_ ( .D(mulout[37]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[37]) );
  DFFARX1 base_multiply_result_reg_36_ ( .D(mulout[36]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[36]) );
  DFFARX1 base_multiply_result_reg_35_ ( .D(mulout[35]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[35]) );
  DFFARX1 base_multiply_result_reg_34_ ( .D(mulout[34]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[34]) );
  DFFARX1 base_multiply_result_reg_33_ ( .D(mulout[33]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[33]) );
  DFFARX1 base_multiply_result_reg_32_ ( .D(mulout[32]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[32]) );
  DFFARX1 base_multiply_result_reg_31_ ( .D(mulout[31]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[31]) );
  DFFARX1 base_multiply_result_reg_30_ ( .D(mulout[30]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[30]) );
  DFFARX1 base_multiply_result_reg_29_ ( .D(mulout[29]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[29]) );
  DFFARX1 base_multiply_result_reg_28_ ( .D(mulout[28]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[28]) );
  DFFARX1 base_multiply_result_reg_27_ ( .D(mulout[27]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[27]) );
  DFFARX1 base_multiply_result_reg_26_ ( .D(mulout[26]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[26]) );
  DFFARX1 base_multiply_result_reg_25_ ( .D(mulout[25]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[25]) );
  DFFARX1 base_multiply_result_reg_24_ ( .D(mulout[24]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[24]) );
  DFFARX1 base_multiply_result_reg_23_ ( .D(mulout[23]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[23]) );
  DFFARX1 mul_output_significand_reg_22_ ( .D(N32), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[22]) );
  DFFARX1 mul_output_significand_reg_21_ ( .D(N31), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[21]) );
  DFFARX1 mul_output_significand_reg_20_ ( .D(N30), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[20]) );
  DFFARX1 mul_output_significand_reg_19_ ( .D(N29), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[19]) );
  DFFARX1 mul_output_significand_reg_18_ ( .D(N28), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[18]) );
  DFFARX1 mul_output_significand_reg_17_ ( .D(N27), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[17]) );
  DFFARX1 mul_output_significand_reg_16_ ( .D(N26), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[16]) );
  DFFARX1 mul_output_significand_reg_15_ ( .D(N25), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[15]) );
  DFFARX1 mul_output_significand_reg_14_ ( .D(N24), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[14]) );
  DFFARX1 mul_output_significand_reg_13_ ( .D(N23), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[13]) );
  DFFARX1 mul_output_significand_reg_12_ ( .D(N22), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[12]) );
  DFFARX1 mul_output_significand_reg_11_ ( .D(N21), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[11]) );
  DFFARX1 mul_output_significand_reg_10_ ( .D(N20), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[10]) );
  DFFARX1 mul_output_significand_reg_9_ ( .D(N19), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[9]) );
  DFFARX1 mul_output_significand_reg_8_ ( .D(N18), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[8]) );
  DFFARX1 mul_output_significand_reg_7_ ( .D(N17), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[7]) );
  DFFARX1 mul_output_significand_reg_6_ ( .D(N16), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[6]) );
  DFFARX1 mul_output_significand_reg_5_ ( .D(N15), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[5]) );
  DFFARX1 mul_output_significand_reg_4_ ( .D(N14), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[4]) );
  DFFARX1 mul_output_significand_reg_3_ ( .D(N13), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[3]) );
  DFFARX1 mul_output_significand_reg_2_ ( .D(N12), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[2]) );
  DFFARX1 mul_output_significand_reg_1_ ( .D(N11), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[1]) );
  DFFARX1 mul_output_significand_reg_0_ ( .D(N10), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[0]) );
  DFFARX1 mul_output_exponent_reg_7_ ( .D(N55), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[30]) );
  DFFARX1 mul_output_exponent_reg_6_ ( .D(N54), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[29]) );
  DFFARX1 mul_output_exponent_reg_5_ ( .D(N53), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[28]) );
  DFFARX1 mul_output_exponent_reg_4_ ( .D(N52), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[27]) );
  DFFARX1 mul_output_exponent_reg_3_ ( .D(N51), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[26]) );
  DFFARX1 mul_output_exponent_reg_2_ ( .D(N50), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[25]) );
  DFFARX1 mul_output_exponent_reg_1_ ( .D(N49), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[24]) );
  DFFARX1 mul_output_exponent_reg_0_ ( .D(N48), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[23]) );
  AND2X1 U3 ( .IN1(base_multiply_result[47]), .IN2(n35), .Q(n32) );
  INVX0 U4 ( .INP(n1), .ZN(n2) );
  OR2X1 U5 ( .IN1(base_multiply_result[47]), .IN2(n24), .Q(n1) );
  INVX0 U6 ( .INP(input_factor_02[31]), .ZN(n3) );
  NOR4X0 U7 ( .IN1(input_factor_01[0]), .IN2(input_factor_01[10]), .IN3(
        input_factor_01[11]), .IN4(input_factor_01[12]), .QN(n7) );
  NOR4X0 U8 ( .IN1(input_factor_01[13]), .IN2(input_factor_01[14]), .IN3(
        input_factor_01[15]), .IN4(input_factor_01[16]), .QN(n6) );
  NOR4X0 U9 ( .IN1(input_factor_01[17]), .IN2(input_factor_01[18]), .IN3(
        input_factor_01[19]), .IN4(input_factor_01[1]), .QN(n5) );
  NOR4X0 U10 ( .IN1(input_factor_01[20]), .IN2(input_factor_01[21]), .IN3(
        input_factor_01[22]), .IN4(input_factor_01[23]), .QN(n4) );
  NAND4X0 U11 ( .IN1(n7), .IN2(n6), .IN3(n5), .IN4(n4), .QN(n23) );
  NOR4X0 U12 ( .IN1(input_factor_01[24]), .IN2(input_factor_01[25]), .IN3(
        input_factor_01[26]), .IN4(input_factor_01[27]), .QN(n11) );
  NOR4X0 U13 ( .IN1(input_factor_01[28]), .IN2(input_factor_01[29]), .IN3(
        input_factor_01[2]), .IN4(input_factor_01[30]), .QN(n10) );
  NOR4X0 U14 ( .IN1(input_factor_01[31]), .IN2(input_factor_01[3]), .IN3(
        input_factor_01[4]), .IN4(input_factor_01[5]), .QN(n9) );
  NOR4X0 U15 ( .IN1(input_factor_01[6]), .IN2(input_factor_01[7]), .IN3(
        input_factor_01[8]), .IN4(input_factor_01[9]), .QN(n8) );
  NAND4X0 U16 ( .IN1(n11), .IN2(n10), .IN3(n9), .IN4(n8), .QN(n22) );
  NOR4X0 U17 ( .IN1(input_factor_02[0]), .IN2(input_factor_02[10]), .IN3(
        input_factor_02[11]), .IN4(input_factor_02[12]), .QN(n15) );
  NOR4X0 U18 ( .IN1(input_factor_02[13]), .IN2(input_factor_02[14]), .IN3(
        input_factor_02[15]), .IN4(input_factor_02[16]), .QN(n14) );
  NOR4X0 U19 ( .IN1(input_factor_02[17]), .IN2(input_factor_02[18]), .IN3(
        input_factor_02[19]), .IN4(input_factor_02[1]), .QN(n13) );
  NOR4X0 U20 ( .IN1(input_factor_02[20]), .IN2(input_factor_02[21]), .IN3(
        input_factor_02[22]), .IN4(input_factor_02[23]), .QN(n12) );
  NAND4X0 U21 ( .IN1(n15), .IN2(n14), .IN3(n13), .IN4(n12), .QN(n21) );
  NOR4X0 U22 ( .IN1(input_factor_02[24]), .IN2(input_factor_02[25]), .IN3(
        input_factor_02[26]), .IN4(input_factor_02[27]), .QN(n19) );
  NOR4X0 U23 ( .IN1(input_factor_02[28]), .IN2(input_factor_02[29]), .IN3(
        input_factor_02[2]), .IN4(input_factor_02[30]), .QN(n18) );
  NOR4X0 U24 ( .IN1(input_factor_02[31]), .IN2(input_factor_02[3]), .IN3(
        input_factor_02[4]), .IN4(input_factor_02[5]), .QN(n17) );
  NOR4X0 U25 ( .IN1(input_factor_02[6]), .IN2(input_factor_02[7]), .IN3(
        input_factor_02[8]), .IN4(input_factor_02[9]), .QN(n16) );
  NAND4X0 U26 ( .IN1(n19), .IN2(n18), .IN3(n17), .IN4(n16), .QN(n20) );
  OA22X1 U27 ( .IN1(n23), .IN2(n22), .IN3(n21), .IN4(n20), .Q(n35) );
  INVX0 U28 ( .INP(n35), .ZN(n24) );
  AO22X1 U29 ( .IN1(n2), .IN2(base_multiply_result[23]), .IN3(n32), .IN4(
        base_multiply_result[24]), .Q(N10) );
  AO22X1 U30 ( .IN1(n2), .IN2(base_multiply_result[24]), .IN3(n32), .IN4(
        base_multiply_result[25]), .Q(N11) );
  AO22X1 U31 ( .IN1(n2), .IN2(base_multiply_result[25]), .IN3(n32), .IN4(
        base_multiply_result[26]), .Q(N12) );
  AO22X1 U32 ( .IN1(n2), .IN2(base_multiply_result[26]), .IN3(n32), .IN4(
        base_multiply_result[27]), .Q(N13) );
  AO22X1 U33 ( .IN1(n2), .IN2(base_multiply_result[27]), .IN3(n32), .IN4(
        base_multiply_result[28]), .Q(N14) );
  AO22X1 U34 ( .IN1(n2), .IN2(base_multiply_result[28]), .IN3(n32), .IN4(
        base_multiply_result[29]), .Q(N15) );
  AO22X1 U35 ( .IN1(n2), .IN2(base_multiply_result[29]), .IN3(n32), .IN4(
        base_multiply_result[30]), .Q(N16) );
  AO22X1 U36 ( .IN1(n2), .IN2(base_multiply_result[30]), .IN3(n32), .IN4(
        base_multiply_result[31]), .Q(N17) );
  AO22X1 U37 ( .IN1(n2), .IN2(base_multiply_result[31]), .IN3(n32), .IN4(
        base_multiply_result[32]), .Q(N18) );
  AO22X1 U38 ( .IN1(n2), .IN2(base_multiply_result[32]), .IN3(n32), .IN4(
        base_multiply_result[33]), .Q(N19) );
  AO22X1 U39 ( .IN1(n2), .IN2(base_multiply_result[33]), .IN3(n32), .IN4(
        base_multiply_result[34]), .Q(N20) );
  AO22X1 U40 ( .IN1(n2), .IN2(base_multiply_result[34]), .IN3(n32), .IN4(
        base_multiply_result[35]), .Q(N21) );
  AO22X1 U41 ( .IN1(n2), .IN2(base_multiply_result[35]), .IN3(n32), .IN4(
        base_multiply_result[36]), .Q(N22) );
  AO22X1 U42 ( .IN1(n2), .IN2(base_multiply_result[36]), .IN3(n32), .IN4(
        base_multiply_result[37]), .Q(N23) );
  AO22X1 U43 ( .IN1(n2), .IN2(base_multiply_result[37]), .IN3(n32), .IN4(
        base_multiply_result[38]), .Q(N24) );
  AO22X1 U44 ( .IN1(n2), .IN2(base_multiply_result[38]), .IN3(n32), .IN4(
        base_multiply_result[39]), .Q(N25) );
  AO22X1 U45 ( .IN1(n2), .IN2(base_multiply_result[39]), .IN3(n32), .IN4(
        base_multiply_result[40]), .Q(N26) );
  AO22X1 U46 ( .IN1(n2), .IN2(base_multiply_result[40]), .IN3(n32), .IN4(
        base_multiply_result[41]), .Q(N27) );
  AO22X1 U47 ( .IN1(n2), .IN2(base_multiply_result[41]), .IN3(n32), .IN4(
        base_multiply_result[42]), .Q(N28) );
  AO22X1 U48 ( .IN1(n2), .IN2(base_multiply_result[42]), .IN3(n32), .IN4(
        base_multiply_result[43]), .Q(N29) );
  AO22X1 U49 ( .IN1(n2), .IN2(base_multiply_result[43]), .IN3(n32), .IN4(
        base_multiply_result[44]), .Q(N30) );
  AO22X1 U50 ( .IN1(n2), .IN2(base_multiply_result[44]), .IN3(n32), .IN4(
        base_multiply_result[45]), .Q(N31) );
  AO22X1 U51 ( .IN1(n2), .IN2(base_multiply_result[45]), .IN3(n32), .IN4(
        base_multiply_result[46]), .Q(N32) );
  MUX21X1 U52 ( .IN1(n2), .IN2(n32), .S(pre_mul_output_exponent[0]), .Q(N48)
         );
  AO21X1 U53 ( .IN1(pre_mul_output_exponent[0]), .IN2(n2), .IN3(n32), .Q(n25)
         );
  NOR3X0 U54 ( .IN1(pre_mul_output_exponent[1]), .IN2(
        pre_mul_output_exponent[0]), .IN3(n1), .QN(n27) );
  AO21X1 U55 ( .IN1(pre_mul_output_exponent[1]), .IN2(n25), .IN3(n27), .Q(N49)
         );
  INVX0 U56 ( .INP(input_factor_01[31]), .ZN(n26) );
  OA221X1 U57 ( .IN1(input_factor_01[31]), .IN2(input_factor_02[31]), .IN3(n26), .IN4(n3), .IN5(n35), .Q(N5) );
  AO221X1 U58 ( .IN1(n2), .IN2(pre_mul_output_exponent[1]), .IN3(n2), .IN4(
        pre_mul_output_exponent[0]), .IN5(n32), .Q(n28) );
  MUX21X1 U59 ( .IN1(n27), .IN2(n28), .S(pre_mul_output_exponent[2]), .Q(N50)
         );
  AND2X1 U60 ( .IN1(n2), .IN2(pre_mul_output_exponent[2]), .Q(n29) );
  OR4X1 U61 ( .IN1(pre_mul_output_exponent[1]), .IN2(
        pre_mul_output_exponent[0]), .IN3(pre_mul_output_exponent[3]), .IN4(
        pre_mul_output_exponent[2]), .Q(n34) );
  NOR2X0 U62 ( .IN1(n1), .IN2(n34), .QN(n31) );
  AO221X1 U63 ( .IN1(pre_mul_output_exponent[3]), .IN2(n29), .IN3(
        pre_mul_output_exponent[3]), .IN4(n28), .IN5(n31), .Q(N51) );
  OA21X1 U64 ( .IN1(base_multiply_result[47]), .IN2(n34), .IN3(n35), .Q(n30)
         );
  MUX21X1 U65 ( .IN1(n31), .IN2(n30), .S(pre_mul_output_exponent[4]), .Q(N52)
         );
  AO221X1 U66 ( .IN1(n2), .IN2(pre_mul_output_exponent[4]), .IN3(n2), .IN4(n34), .IN5(n32), .Q(n33) );
  NOR4X0 U67 ( .IN1(pre_mul_output_exponent[5]), .IN2(
        pre_mul_output_exponent[4]), .IN3(n34), .IN4(n1), .QN(n37) );
  AO21X1 U68 ( .IN1(pre_mul_output_exponent[5]), .IN2(n33), .IN3(n37), .Q(N53)
         );
  OR3X1 U69 ( .IN1(pre_mul_output_exponent[5]), .IN2(
        pre_mul_output_exponent[4]), .IN3(n34), .Q(n36) );
  OA21X1 U70 ( .IN1(base_multiply_result[47]), .IN2(n36), .IN3(n35), .Q(n39)
         );
  INVX0 U71 ( .INP(n37), .ZN(n38) );
  NOR2X0 U72 ( .IN1(pre_mul_output_exponent[6]), .IN2(n38), .QN(n41) );
  AO21X1 U73 ( .IN1(pre_mul_output_exponent[6]), .IN2(n39), .IN3(n41), .Q(N54)
         );
  AO21X1 U74 ( .IN1(n2), .IN2(pre_mul_output_exponent[6]), .IN3(n39), .Q(n40)
         );
  MUX21X1 U75 ( .IN1(n41), .IN2(n40), .S(pre_mul_output_exponent[7]), .Q(N55)
         );
endmodule


module cla51squ_5 ( out, a, b );
  output [50:0] out;
  input [50:0] a;
  input [50:0] b;
  wire   intadd_5_CI, intadd_5_n24, intadd_5_n23, intadd_5_n22, intadd_5_n21,
         intadd_5_n20, intadd_5_n19, intadd_5_n18, intadd_5_n17, intadd_5_n16,
         intadd_5_n15, intadd_5_n14, intadd_5_n13, intadd_5_n12, intadd_5_n11,
         intadd_5_n10, intadd_5_n9, intadd_5_n8, intadd_5_n7, intadd_5_n6,
         intadd_5_n5, intadd_5_n4, intadd_5_n3, intadd_5_n2, intadd_5_n1, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14;

  FADDX1 intadd_5_U25 ( .A(b[23]), .B(a[23]), .CI(intadd_5_CI), .CO(
        intadd_5_n24), .S(out[23]) );
  FADDX1 intadd_5_U24 ( .A(b[24]), .B(a[24]), .CI(intadd_5_n24), .CO(
        intadd_5_n23), .S(out[24]) );
  FADDX1 intadd_5_U23 ( .A(b[25]), .B(a[25]), .CI(intadd_5_n23), .CO(
        intadd_5_n22), .S(out[25]) );
  FADDX1 intadd_5_U22 ( .A(b[26]), .B(a[26]), .CI(intadd_5_n22), .CO(
        intadd_5_n21), .S(out[26]) );
  FADDX1 intadd_5_U21 ( .A(b[27]), .B(a[27]), .CI(intadd_5_n21), .CO(
        intadd_5_n20), .S(out[27]) );
  FADDX1 intadd_5_U20 ( .A(b[28]), .B(a[28]), .CI(intadd_5_n20), .CO(
        intadd_5_n19), .S(out[28]) );
  FADDX1 intadd_5_U19 ( .A(b[29]), .B(a[29]), .CI(intadd_5_n19), .CO(
        intadd_5_n18), .S(out[29]) );
  FADDX1 intadd_5_U18 ( .A(b[30]), .B(a[30]), .CI(intadd_5_n18), .CO(
        intadd_5_n17), .S(out[30]) );
  FADDX1 intadd_5_U17 ( .A(b[31]), .B(a[31]), .CI(intadd_5_n17), .CO(
        intadd_5_n16), .S(out[31]) );
  FADDX1 intadd_5_U16 ( .A(b[32]), .B(a[32]), .CI(intadd_5_n16), .CO(
        intadd_5_n15), .S(out[32]) );
  FADDX1 intadd_5_U15 ( .A(b[33]), .B(a[33]), .CI(intadd_5_n15), .CO(
        intadd_5_n14), .S(out[33]) );
  FADDX1 intadd_5_U14 ( .A(b[34]), .B(a[34]), .CI(intadd_5_n14), .CO(
        intadd_5_n13), .S(out[34]) );
  FADDX1 intadd_5_U13 ( .A(b[35]), .B(a[35]), .CI(intadd_5_n13), .CO(
        intadd_5_n12), .S(out[35]) );
  FADDX1 intadd_5_U12 ( .A(b[36]), .B(a[36]), .CI(intadd_5_n12), .CO(
        intadd_5_n11), .S(out[36]) );
  FADDX1 intadd_5_U11 ( .A(b[37]), .B(a[37]), .CI(intadd_5_n11), .CO(
        intadd_5_n10), .S(out[37]) );
  FADDX1 intadd_5_U10 ( .A(b[38]), .B(a[38]), .CI(intadd_5_n10), .CO(
        intadd_5_n9), .S(out[38]) );
  FADDX1 intadd_5_U9 ( .A(b[39]), .B(a[39]), .CI(intadd_5_n9), .CO(intadd_5_n8), .S(out[39]) );
  FADDX1 intadd_5_U8 ( .A(b[40]), .B(a[40]), .CI(intadd_5_n8), .CO(intadd_5_n7), .S(out[40]) );
  FADDX1 intadd_5_U7 ( .A(b[41]), .B(a[41]), .CI(intadd_5_n7), .CO(intadd_5_n6), .S(out[41]) );
  FADDX1 intadd_5_U6 ( .A(b[42]), .B(a[42]), .CI(intadd_5_n6), .CO(intadd_5_n5), .S(out[42]) );
  FADDX1 intadd_5_U5 ( .A(b[43]), .B(a[43]), .CI(intadd_5_n5), .CO(intadd_5_n4), .S(out[43]) );
  FADDX1 intadd_5_U4 ( .A(b[44]), .B(a[44]), .CI(intadd_5_n4), .CO(intadd_5_n3), .S(out[44]) );
  FADDX1 intadd_5_U3 ( .A(b[45]), .B(a[45]), .CI(intadd_5_n3), .CO(intadd_5_n2), .S(out[45]) );
  FADDX1 intadd_5_U2 ( .A(b[46]), .B(a[46]), .CI(intadd_5_n2), .CO(intadd_5_n1), .S(out[46]) );
  OA21X1 U2 ( .IN1(b[9]), .IN2(a[9]), .IN3(a[8]), .Q(n1) );
  AO22X1 U3 ( .IN1(b[9]), .IN2(a[9]), .IN3(b[8]), .IN4(n1), .Q(n2) );
  AO222X1 U4 ( .IN1(b[10]), .IN2(a[10]), .IN3(b[10]), .IN4(n2), .IN5(a[10]), 
        .IN6(n2), .Q(n3) );
  AO222X1 U5 ( .IN1(b[11]), .IN2(a[11]), .IN3(b[11]), .IN4(n3), .IN5(a[11]), 
        .IN6(n3), .Q(n4) );
  AO222X1 U6 ( .IN1(b[12]), .IN2(a[12]), .IN3(b[12]), .IN4(n4), .IN5(a[12]), 
        .IN6(n4), .Q(n5) );
  AO222X1 U7 ( .IN1(b[13]), .IN2(a[13]), .IN3(b[13]), .IN4(n5), .IN5(a[13]), 
        .IN6(n5), .Q(n6) );
  AO222X1 U8 ( .IN1(b[14]), .IN2(a[14]), .IN3(b[14]), .IN4(n6), .IN5(a[14]), 
        .IN6(n6), .Q(n7) );
  AO222X1 U9 ( .IN1(b[15]), .IN2(a[15]), .IN3(b[15]), .IN4(n7), .IN5(a[15]), 
        .IN6(n7), .Q(n8) );
  AO222X1 U10 ( .IN1(b[16]), .IN2(a[16]), .IN3(b[16]), .IN4(n8), .IN5(a[16]), 
        .IN6(n8), .Q(n9) );
  AO222X1 U11 ( .IN1(b[17]), .IN2(a[17]), .IN3(b[17]), .IN4(n9), .IN5(a[17]), 
        .IN6(n9), .Q(n10) );
  AO222X1 U12 ( .IN1(b[18]), .IN2(a[18]), .IN3(b[18]), .IN4(n10), .IN5(a[18]), 
        .IN6(n10), .Q(n11) );
  AO222X1 U13 ( .IN1(b[19]), .IN2(a[19]), .IN3(b[19]), .IN4(n11), .IN5(a[19]), 
        .IN6(n11), .Q(n12) );
  AO222X1 U14 ( .IN1(b[20]), .IN2(a[20]), .IN3(b[20]), .IN4(n12), .IN5(a[20]), 
        .IN6(n12), .Q(n13) );
  AO222X1 U15 ( .IN1(b[21]), .IN2(a[21]), .IN3(b[21]), .IN4(n13), .IN5(a[21]), 
        .IN6(n13), .Q(n14) );
  AO222X1 U16 ( .IN1(b[22]), .IN2(a[22]), .IN3(b[22]), .IN4(n14), .IN5(a[22]), 
        .IN6(n14), .Q(intadd_5_CI) );
  XOR3X1 U17 ( .IN1(intadd_5_n1), .IN2(a[47]), .IN3(b[47]), .Q(out[47]) );
endmodule


module csa51squ_49 ( sumout, in1, in2, in3, cout_50_, cout_49_, cout_48_, 
        cout_47_, cout_46_, cout_44_, cout_42_, cout_40_, cout_38_, cout_36_, 
        cout_34_, cout_32_, cout_30_, cout_28_, cout_27_, cout_7__BAR, cout_6_, 
        cout_5_, cout_4_, cout_3_, cout_2_, cout_1_, cout_0_, cout_8__BAR, 
        cout_9__BAR, cout_10__BAR, cout_11__BAR, cout_12__BAR, cout_13__BAR, 
        cout_14__BAR, cout_15__BAR, cout_16__BAR, cout_17__BAR, cout_18__BAR, 
        cout_19__BAR, cout_20__BAR, cout_21__BAR, cout_22__BAR, cout_23__BAR, 
        cout_24__BAR, cout_25__BAR, cout_26__BAR, cout_29__BAR, cout_31__BAR, 
        cout_33__BAR, cout_35__BAR, cout_37__BAR, cout_39__BAR, cout_41__BAR, 
        cout_43__BAR, cout_45__BAR );
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  output cout_50_, cout_49_, cout_48_, cout_47_, cout_46_, cout_44_, cout_42_,
         cout_40_, cout_38_, cout_36_, cout_34_, cout_32_, cout_30_, cout_28_,
         cout_27_, cout_7__BAR, cout_6_, cout_5_, cout_4_, cout_3_, cout_2_,
         cout_1_, cout_0_, cout_8__BAR, cout_9__BAR, cout_10__BAR,
         cout_11__BAR, cout_12__BAR, cout_13__BAR, cout_14__BAR, cout_15__BAR,
         cout_16__BAR, cout_17__BAR, cout_18__BAR, cout_19__BAR, cout_20__BAR,
         cout_21__BAR, cout_22__BAR, cout_23__BAR, cout_24__BAR, cout_25__BAR,
         cout_26__BAR, cout_29__BAR, cout_31__BAR, cout_33__BAR, cout_35__BAR,
         cout_37__BAR, cout_39__BAR, cout_41__BAR, cout_43__BAR, cout_45__BAR;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11;

  NAND2X0 U1 ( .IN1(in2[8]), .IN2(in1[8]), .QN(cout_8__BAR) );
  NAND2X0 U2 ( .IN1(in2[9]), .IN2(in1[9]), .QN(cout_9__BAR) );
  NAND2X0 U3 ( .IN1(in2[10]), .IN2(in1[10]), .QN(cout_10__BAR) );
  NAND2X0 U4 ( .IN1(in2[11]), .IN2(in1[11]), .QN(cout_11__BAR) );
  NAND2X0 U5 ( .IN1(in2[12]), .IN2(in1[12]), .QN(cout_12__BAR) );
  NAND2X0 U6 ( .IN1(in2[13]), .IN2(in1[13]), .QN(cout_13__BAR) );
  NAND2X0 U7 ( .IN1(in2[14]), .IN2(in1[14]), .QN(cout_14__BAR) );
  NAND2X0 U8 ( .IN1(in2[15]), .IN2(in1[15]), .QN(cout_15__BAR) );
  NAND2X0 U9 ( .IN1(in2[16]), .IN2(in1[16]), .QN(cout_16__BAR) );
  NAND2X0 U10 ( .IN1(in2[17]), .IN2(in1[17]), .QN(cout_17__BAR) );
  NAND2X0 U11 ( .IN1(in2[18]), .IN2(in1[18]), .QN(cout_18__BAR) );
  NAND2X0 U12 ( .IN1(in2[19]), .IN2(in1[19]), .QN(cout_19__BAR) );
  NAND2X0 U13 ( .IN1(in2[20]), .IN2(in1[20]), .QN(cout_20__BAR) );
  NAND2X0 U14 ( .IN1(in2[21]), .IN2(in1[21]), .QN(cout_21__BAR) );
  NAND2X0 U15 ( .IN1(in2[22]), .IN2(in1[22]), .QN(cout_22__BAR) );
  NAND2X0 U16 ( .IN1(in2[23]), .IN2(in1[23]), .QN(cout_23__BAR) );
  NAND2X0 U17 ( .IN1(in2[24]), .IN2(in1[24]), .QN(cout_24__BAR) );
  NAND2X0 U18 ( .IN1(in2[25]), .IN2(in1[25]), .QN(cout_25__BAR) );
  NAND2X0 U19 ( .IN1(in2[26]), .IN2(in1[26]), .QN(cout_26__BAR) );
  NAND2X0 U20 ( .IN1(in2[29]), .IN2(in1[29]), .QN(cout_29__BAR) );
  NAND2X0 U21 ( .IN1(in2[31]), .IN2(in1[31]), .QN(cout_31__BAR) );
  NAND2X0 U22 ( .IN1(in2[33]), .IN2(in1[33]), .QN(cout_33__BAR) );
  NAND2X0 U23 ( .IN1(in2[35]), .IN2(in1[35]), .QN(cout_35__BAR) );
  NAND2X0 U24 ( .IN1(in2[37]), .IN2(in1[37]), .QN(cout_37__BAR) );
  NAND2X0 U25 ( .IN1(in2[39]), .IN2(in1[39]), .QN(cout_39__BAR) );
  NAND2X0 U26 ( .IN1(in2[41]), .IN2(in1[41]), .QN(cout_41__BAR) );
  NAND2X0 U27 ( .IN1(in2[43]), .IN2(in1[43]), .QN(cout_43__BAR) );
  NAND2X0 U28 ( .IN1(in2[45]), .IN2(in1[45]), .QN(cout_45__BAR) );
  NAND2X0 U29 ( .IN1(in2[7]), .IN2(in1[7]), .QN(cout_7__BAR) );
  NAND2X0 U30 ( .IN1(n1), .IN2(cout_27_), .QN(sumout[27]) );
  NAND2X0 U31 ( .IN1(in1[27]), .IN2(in2[27]), .QN(n1) );
  NAND2X0 U32 ( .IN1(n2), .IN2(cout_28_), .QN(sumout[28]) );
  NAND2X0 U33 ( .IN1(in1[28]), .IN2(in2[28]), .QN(n2) );
  NAND2X0 U34 ( .IN1(n3), .IN2(cout_30_), .QN(sumout[30]) );
  NAND2X0 U35 ( .IN1(in1[30]), .IN2(in2[30]), .QN(n3) );
  NAND2X0 U36 ( .IN1(n4), .IN2(cout_32_), .QN(sumout[32]) );
  NAND2X0 U37 ( .IN1(in1[32]), .IN2(in2[32]), .QN(n4) );
  NAND2X0 U38 ( .IN1(n5), .IN2(cout_34_), .QN(sumout[34]) );
  NAND2X0 U39 ( .IN1(in1[34]), .IN2(in2[34]), .QN(n5) );
  NAND2X0 U40 ( .IN1(n6), .IN2(cout_36_), .QN(sumout[36]) );
  NAND2X0 U41 ( .IN1(in1[36]), .IN2(in2[36]), .QN(n6) );
  NAND2X0 U42 ( .IN1(n7), .IN2(cout_38_), .QN(sumout[38]) );
  NAND2X0 U43 ( .IN1(in1[38]), .IN2(in2[38]), .QN(n7) );
  NAND2X0 U44 ( .IN1(n8), .IN2(cout_40_), .QN(sumout[40]) );
  NAND2X0 U45 ( .IN1(in1[40]), .IN2(in2[40]), .QN(n8) );
  NAND2X0 U46 ( .IN1(n9), .IN2(cout_42_), .QN(sumout[42]) );
  NAND2X0 U47 ( .IN1(in1[42]), .IN2(in2[42]), .QN(n9) );
  NAND2X0 U48 ( .IN1(n10), .IN2(cout_44_), .QN(sumout[44]) );
  NAND2X0 U49 ( .IN1(in1[44]), .IN2(in2[44]), .QN(n10) );
  NAND2X0 U50 ( .IN1(n11), .IN2(cout_46_), .QN(sumout[46]) );
  NAND2X0 U51 ( .IN1(in1[46]), .IN2(in2[46]), .QN(n11) );
  OR2X1 U52 ( .IN1(in2[27]), .IN2(in1[27]), .Q(cout_27_) );
  OR2X1 U53 ( .IN1(in2[28]), .IN2(in1[28]), .Q(cout_28_) );
  OR2X1 U54 ( .IN1(in2[30]), .IN2(in1[30]), .Q(cout_30_) );
  OR2X1 U55 ( .IN1(in2[32]), .IN2(in1[32]), .Q(cout_32_) );
  OR2X1 U56 ( .IN1(in2[34]), .IN2(in1[34]), .Q(cout_34_) );
  OR2X1 U57 ( .IN1(in2[36]), .IN2(in1[36]), .Q(cout_36_) );
  OR2X1 U58 ( .IN1(in2[38]), .IN2(in1[38]), .Q(cout_38_) );
  OR2X1 U59 ( .IN1(in2[40]), .IN2(in1[40]), .Q(cout_40_) );
  OR2X1 U60 ( .IN1(in2[42]), .IN2(in1[42]), .Q(cout_42_) );
  OR2X1 U61 ( .IN1(in2[44]), .IN2(in1[44]), .Q(cout_44_) );
  OR2X1 U62 ( .IN1(in2[46]), .IN2(in1[46]), .Q(cout_46_) );
  OA21X1 U63 ( .IN1(in2[8]), .IN2(in1[8]), .IN3(cout_8__BAR), .Q(sumout[8]) );
  OA21X1 U64 ( .IN1(in2[9]), .IN2(in1[9]), .IN3(cout_9__BAR), .Q(sumout[9]) );
  OA21X1 U65 ( .IN1(in2[10]), .IN2(in1[10]), .IN3(cout_10__BAR), .Q(sumout[10]) );
  OA21X1 U66 ( .IN1(in2[11]), .IN2(in1[11]), .IN3(cout_11__BAR), .Q(sumout[11]) );
  OA21X1 U67 ( .IN1(in2[12]), .IN2(in1[12]), .IN3(cout_12__BAR), .Q(sumout[12]) );
  OA21X1 U68 ( .IN1(in2[13]), .IN2(in1[13]), .IN3(cout_13__BAR), .Q(sumout[13]) );
  OA21X1 U69 ( .IN1(in2[14]), .IN2(in1[14]), .IN3(cout_14__BAR), .Q(sumout[14]) );
  OA21X1 U70 ( .IN1(in2[15]), .IN2(in1[15]), .IN3(cout_15__BAR), .Q(sumout[15]) );
  OA21X1 U71 ( .IN1(in2[16]), .IN2(in1[16]), .IN3(cout_16__BAR), .Q(sumout[16]) );
  OA21X1 U72 ( .IN1(in2[17]), .IN2(in1[17]), .IN3(cout_17__BAR), .Q(sumout[17]) );
  OA21X1 U73 ( .IN1(in2[18]), .IN2(in1[18]), .IN3(cout_18__BAR), .Q(sumout[18]) );
  OA21X1 U74 ( .IN1(in2[19]), .IN2(in1[19]), .IN3(cout_19__BAR), .Q(sumout[19]) );
  OA21X1 U75 ( .IN1(in2[20]), .IN2(in1[20]), .IN3(cout_20__BAR), .Q(sumout[20]) );
  OA21X1 U76 ( .IN1(in2[21]), .IN2(in1[21]), .IN3(cout_21__BAR), .Q(sumout[21]) );
  OA21X1 U77 ( .IN1(in2[22]), .IN2(in1[22]), .IN3(cout_22__BAR), .Q(sumout[22]) );
  OA21X1 U78 ( .IN1(in2[23]), .IN2(in1[23]), .IN3(cout_23__BAR), .Q(sumout[23]) );
  OA21X1 U79 ( .IN1(in2[24]), .IN2(in1[24]), .IN3(cout_24__BAR), .Q(sumout[24]) );
  OA21X1 U80 ( .IN1(in2[25]), .IN2(in1[25]), .IN3(cout_25__BAR), .Q(sumout[25]) );
  OA21X1 U81 ( .IN1(in2[26]), .IN2(in1[26]), .IN3(cout_26__BAR), .Q(sumout[26]) );
  OA21X1 U82 ( .IN1(in2[29]), .IN2(in1[29]), .IN3(cout_29__BAR), .Q(sumout[29]) );
  OA21X1 U83 ( .IN1(in2[31]), .IN2(in1[31]), .IN3(cout_31__BAR), .Q(sumout[31]) );
  OA21X1 U84 ( .IN1(in2[33]), .IN2(in1[33]), .IN3(cout_33__BAR), .Q(sumout[33]) );
  OA21X1 U85 ( .IN1(in2[35]), .IN2(in1[35]), .IN3(cout_35__BAR), .Q(sumout[35]) );
  OA21X1 U86 ( .IN1(in2[37]), .IN2(in1[37]), .IN3(cout_37__BAR), .Q(sumout[37]) );
  OA21X1 U87 ( .IN1(in2[39]), .IN2(in1[39]), .IN3(cout_39__BAR), .Q(sumout[39]) );
  OA21X1 U88 ( .IN1(in2[41]), .IN2(in1[41]), .IN3(cout_41__BAR), .Q(sumout[41]) );
  OA21X1 U89 ( .IN1(in2[43]), .IN2(in1[43]), .IN3(cout_43__BAR), .Q(sumout[43]) );
  OA21X1 U90 ( .IN1(in2[45]), .IN2(in1[45]), .IN3(cout_45__BAR), .Q(sumout[45]) );
  XOR2X1 U91 ( .IN1(in1[47]), .IN2(in2[47]), .Q(sumout[47]) );
endmodule


module csa51squ_50 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;


  AO222X1 U1 ( .IN1(in2[6]), .IN2(in3[6]), .IN3(in2[6]), .IN4(in1[6]), .IN5(
        in3[6]), .IN6(in1[6]), .Q(cout[6]) );
  FADDX1 U2 ( .A(in1[10]), .B(in2[10]), .CI(in3[10]), .CO(cout[10]), .S(
        sumout[10]) );
  FADDX1 U3 ( .A(in1[11]), .B(in2[11]), .CI(in3[11]), .CO(cout[11]), .S(
        sumout[11]) );
  FADDX1 U4 ( .A(in1[12]), .B(in2[12]), .CI(in3[12]), .CO(cout[12]), .S(
        sumout[12]) );
  FADDX1 U5 ( .A(in1[13]), .B(in2[13]), .CI(in3[13]), .CO(cout[13]), .S(
        sumout[13]) );
  FADDX1 U6 ( .A(in1[14]), .B(in2[14]), .CI(in3[14]), .CO(cout[14]), .S(
        sumout[14]) );
  FADDX1 U7 ( .A(in1[15]), .B(in2[15]), .CI(in3[15]), .CO(cout[15]), .S(
        sumout[15]) );
  FADDX1 U8 ( .A(in1[16]), .B(in2[16]), .CI(in3[16]), .CO(cout[16]), .S(
        sumout[16]) );
  FADDX1 U9 ( .A(in1[17]), .B(in2[17]), .CI(in3[17]), .CO(cout[17]), .S(
        sumout[17]) );
  FADDX1 U10 ( .A(in1[18]), .B(in2[18]), .CI(in3[18]), .CO(cout[18]), .S(
        sumout[18]) );
  FADDX1 U11 ( .A(in1[19]), .B(in2[19]), .CI(in3[19]), .CO(cout[19]), .S(
        sumout[19]) );
  FADDX1 U12 ( .A(in1[20]), .B(in2[20]), .CI(in3[20]), .CO(cout[20]), .S(
        sumout[20]) );
  FADDX1 U13 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U14 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U15 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U16 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U17 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U18 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U19 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U20 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U21 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U22 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U23 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U24 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
  FADDX1 U25 ( .A(in1[33]), .B(in2[33]), .CI(in3[33]), .CO(cout[33]), .S(
        sumout[33]) );
  FADDX1 U26 ( .A(in1[34]), .B(in2[34]), .CI(in3[34]), .CO(cout[34]), .S(
        sumout[34]) );
  FADDX1 U27 ( .A(in1[35]), .B(in2[35]), .CI(in3[35]), .CO(cout[35]), .S(
        sumout[35]) );
  FADDX1 U28 ( .A(in1[36]), .B(in2[36]), .CI(in3[36]), .CO(cout[36]), .S(
        sumout[36]) );
  FADDX1 U29 ( .A(in1[37]), .B(in2[37]), .CI(in3[37]), .CO(cout[37]), .S(
        sumout[37]) );
  FADDX1 U30 ( .A(in1[38]), .B(in2[38]), .CI(in3[38]), .CO(cout[38]), .S(
        sumout[38]) );
  FADDX1 U31 ( .A(in1[39]), .B(in2[39]), .CI(in3[39]), .CO(cout[39]), .S(
        sumout[39]) );
  FADDX1 U32 ( .A(in1[40]), .B(in2[40]), .CI(in3[40]), .CO(cout[40]), .S(
        sumout[40]) );
  FADDX1 U33 ( .A(in1[41]), .B(in2[41]), .CI(in3[41]), .CO(cout[41]), .S(
        sumout[41]) );
  FADDX1 U34 ( .A(in1[42]), .B(in2[42]), .CI(in3[42]), .CO(cout[42]), .S(
        sumout[42]) );
  FADDX1 U35 ( .A(in1[43]), .B(in2[43]), .CI(in3[43]), .CO(cout[43]), .S(
        sumout[43]) );
  FADDX1 U36 ( .A(in1[44]), .B(in2[44]), .CI(in3[44]), .CO(cout[44]), .S(
        sumout[44]) );
  FADDX1 U37 ( .A(in1[45]), .B(in2[45]), .CI(in3[45]), .CO(cout[45]), .S(
        sumout[45]) );
  FADDX1 U38 ( .A(in1[46]), .B(in2[46]), .CI(in3[46]), .CO(cout[46]), .S(
        sumout[46]) );
  XOR3X1 U39 ( .IN1(in2[47]), .IN2(in3[47]), .IN3(in1[47]), .Q(sumout[47]) );
  FADDX1 U40 ( .A(in1[7]), .B(in2[7]), .CI(in3[7]), .CO(cout[7]), .S(sumout[7]) );
  FADDX1 U41 ( .A(in1[8]), .B(in2[8]), .CI(in3[8]), .CO(cout[8]), .S(sumout[8]) );
  FADDX1 U42 ( .A(in1[9]), .B(in2[9]), .CI(in3[9]), .CO(cout[9]), .S(sumout[9]) );
endmodule


module csa51squ_51 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14;

  AND2X1 U1 ( .IN1(in2[7]), .IN2(in1[7]), .Q(cout[7]) );
  NOR2X0 U2 ( .IN1(in2[7]), .IN2(in1[7]), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(cout[7]), .QN(sumout[7]) );
  AND2X1 U4 ( .IN1(in2[8]), .IN2(in1[8]), .Q(cout[8]) );
  NOR2X0 U5 ( .IN1(in2[8]), .IN2(in1[8]), .QN(n2) );
  NOR2X0 U6 ( .IN1(n2), .IN2(cout[8]), .QN(sumout[8]) );
  AND2X1 U7 ( .IN1(in2[9]), .IN2(in1[9]), .Q(cout[9]) );
  NOR2X0 U8 ( .IN1(in2[9]), .IN2(in1[9]), .QN(n3) );
  NOR2X0 U9 ( .IN1(n3), .IN2(cout[9]), .QN(sumout[9]) );
  AND2X1 U10 ( .IN1(in2[10]), .IN2(in1[10]), .Q(cout[10]) );
  NOR2X0 U11 ( .IN1(in2[10]), .IN2(in1[10]), .QN(n4) );
  NOR2X0 U12 ( .IN1(n4), .IN2(cout[10]), .QN(sumout[10]) );
  AND2X1 U13 ( .IN1(in2[11]), .IN2(in1[11]), .Q(cout[11]) );
  NOR2X0 U14 ( .IN1(in2[11]), .IN2(in1[11]), .QN(n5) );
  NOR2X0 U15 ( .IN1(n5), .IN2(cout[11]), .QN(sumout[11]) );
  AND2X1 U16 ( .IN1(in2[12]), .IN2(in1[12]), .Q(cout[12]) );
  NOR2X0 U17 ( .IN1(in2[12]), .IN2(in1[12]), .QN(n6) );
  NOR2X0 U18 ( .IN1(n6), .IN2(cout[12]), .QN(sumout[12]) );
  AND2X1 U19 ( .IN1(in3[40]), .IN2(in2[40]), .Q(cout[40]) );
  NOR2X0 U20 ( .IN1(in3[40]), .IN2(in2[40]), .QN(n7) );
  NOR2X0 U21 ( .IN1(n7), .IN2(cout[40]), .QN(sumout[40]) );
  AND2X1 U22 ( .IN1(in3[41]), .IN2(in2[41]), .Q(cout[41]) );
  NOR2X0 U23 ( .IN1(in3[41]), .IN2(in2[41]), .QN(n8) );
  NOR2X0 U24 ( .IN1(n8), .IN2(cout[41]), .QN(sumout[41]) );
  AND2X1 U25 ( .IN1(in3[42]), .IN2(in2[42]), .Q(cout[42]) );
  NOR2X0 U26 ( .IN1(in3[42]), .IN2(in2[42]), .QN(n9) );
  NOR2X0 U27 ( .IN1(n9), .IN2(cout[42]), .QN(sumout[42]) );
  AND2X1 U28 ( .IN1(in3[43]), .IN2(in2[43]), .Q(cout[43]) );
  NOR2X0 U29 ( .IN1(in3[43]), .IN2(in2[43]), .QN(n10) );
  NOR2X0 U30 ( .IN1(n10), .IN2(cout[43]), .QN(sumout[43]) );
  AND2X1 U31 ( .IN1(in3[44]), .IN2(in2[44]), .Q(cout[44]) );
  NOR2X0 U32 ( .IN1(in3[44]), .IN2(in2[44]), .QN(n11) );
  NOR2X0 U33 ( .IN1(n11), .IN2(cout[44]), .QN(sumout[44]) );
  AND2X1 U34 ( .IN1(in3[45]), .IN2(in2[45]), .Q(cout[45]) );
  NOR2X0 U35 ( .IN1(in3[45]), .IN2(in2[45]), .QN(n12) );
  NOR2X0 U36 ( .IN1(n12), .IN2(cout[45]), .QN(sumout[45]) );
  AND2X1 U37 ( .IN1(in3[46]), .IN2(in2[46]), .Q(cout[46]) );
  NOR2X0 U38 ( .IN1(in3[46]), .IN2(in2[46]), .QN(n13) );
  NOR2X0 U39 ( .IN1(n13), .IN2(cout[46]), .QN(sumout[46]) );
  INVX0 U40 ( .INP(in3[47]), .ZN(sumout[47]) );
  AND2X1 U41 ( .IN1(in2[5]), .IN2(in1[5]), .Q(cout[5]) );
  AND2X1 U42 ( .IN1(in2[6]), .IN2(in1[6]), .Q(cout[6]) );
  NOR2X0 U43 ( .IN1(in2[6]), .IN2(in1[6]), .QN(n14) );
  NOR2X0 U44 ( .IN1(n14), .IN2(cout[6]), .QN(sumout[6]) );
  FADDX1 U45 ( .A(in1[13]), .B(in2[13]), .CI(in3[13]), .CO(cout[13]), .S(
        sumout[13]) );
  FADDX1 U46 ( .A(in1[14]), .B(in2[14]), .CI(in3[14]), .CO(cout[14]), .S(
        sumout[14]) );
  FADDX1 U47 ( .A(in1[15]), .B(in2[15]), .CI(in3[15]), .CO(cout[15]), .S(
        sumout[15]) );
  FADDX1 U48 ( .A(in1[16]), .B(in2[16]), .CI(in3[16]), .CO(cout[16]), .S(
        sumout[16]) );
  FADDX1 U49 ( .A(in1[17]), .B(in2[17]), .CI(in3[17]), .CO(cout[17]), .S(
        sumout[17]) );
  FADDX1 U50 ( .A(in1[18]), .B(in2[18]), .CI(in3[18]), .CO(cout[18]), .S(
        sumout[18]) );
  FADDX1 U51 ( .A(in1[19]), .B(in2[19]), .CI(in3[19]), .CO(cout[19]), .S(
        sumout[19]) );
  FADDX1 U52 ( .A(in1[20]), .B(in2[20]), .CI(in3[20]), .CO(cout[20]), .S(
        sumout[20]) );
  FADDX1 U53 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U54 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U55 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U56 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U57 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U58 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U59 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U60 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U61 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U62 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U63 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U64 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
  FADDX1 U65 ( .A(in1[33]), .B(in2[33]), .CI(in3[33]), .CO(cout[33]), .S(
        sumout[33]) );
  FADDX1 U66 ( .A(in1[34]), .B(in2[34]), .CI(in3[34]), .CO(cout[34]), .S(
        sumout[34]) );
  FADDX1 U67 ( .A(in1[35]), .B(in2[35]), .CI(in3[35]), .CO(cout[35]), .S(
        sumout[35]) );
  FADDX1 U68 ( .A(in1[36]), .B(in2[36]), .CI(in3[36]), .CO(cout[36]), .S(
        sumout[36]) );
  FADDX1 U69 ( .A(in1[37]), .B(in2[37]), .CI(in3[37]), .CO(cout[37]), .S(
        sumout[37]) );
  FADDX1 U70 ( .A(in1[38]), .B(in2[38]), .CI(in3[38]), .CO(cout[38]), .S(
        sumout[38]) );
  FADDX1 U71 ( .A(in1[39]), .B(in2[39]), .CI(in3[39]), .CO(cout[39]), .S(
        sumout[39]) );
endmodule


module csa51squ_52 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17;

  NBUFFX2 U1 ( .INP(in1[6]), .Z(sumout[6]) );
  NBUFFX2 U2 ( .INP(in1[7]), .Z(sumout[7]) );
  NBUFFX2 U3 ( .INP(in1[8]), .Z(sumout[8]) );
  NBUFFX2 U4 ( .INP(in1[9]), .Z(sumout[9]) );
  NBUFFX2 U5 ( .INP(in1[10]), .Z(sumout[10]) );
  NBUFFX2 U6 ( .INP(in1[11]), .Z(sumout[11]) );
  AND2X1 U7 ( .IN1(in3[13]), .IN2(in1[13]), .Q(cout[13]) );
  NOR2X0 U8 ( .IN1(in3[13]), .IN2(in1[13]), .QN(n7) );
  NOR2X0 U9 ( .IN1(n7), .IN2(cout[13]), .QN(sumout[13]) );
  AND2X1 U10 ( .IN1(in3[15]), .IN2(in1[15]), .Q(cout[15]) );
  NOR2X0 U11 ( .IN1(in3[15]), .IN2(in1[15]), .QN(n8) );
  NOR2X0 U12 ( .IN1(n8), .IN2(cout[15]), .QN(sumout[15]) );
  AND2X1 U13 ( .IN1(in3[17]), .IN2(in1[17]), .Q(cout[17]) );
  NOR2X0 U14 ( .IN1(in3[17]), .IN2(in1[17]), .QN(n9) );
  NOR2X0 U15 ( .IN1(n9), .IN2(cout[17]), .QN(sumout[17]) );
  AND2X1 U16 ( .IN1(in3[43]), .IN2(in2[43]), .Q(cout[43]) );
  NOR2X0 U17 ( .IN1(in3[43]), .IN2(in2[43]), .QN(n10) );
  NOR2X0 U18 ( .IN1(n10), .IN2(cout[43]), .QN(sumout[43]) );
  AND2X1 U19 ( .IN1(in3[44]), .IN2(in2[44]), .Q(cout[44]) );
  NOR2X0 U20 ( .IN1(in3[44]), .IN2(in2[44]), .QN(n11) );
  NOR2X0 U21 ( .IN1(n11), .IN2(cout[44]), .QN(sumout[44]) );
  AND2X1 U22 ( .IN1(in3[45]), .IN2(in2[45]), .Q(cout[45]) );
  NOR2X0 U23 ( .IN1(in3[45]), .IN2(in2[45]), .QN(n12) );
  NOR2X0 U24 ( .IN1(n12), .IN2(cout[45]), .QN(sumout[45]) );
  AND2X1 U25 ( .IN1(in3[46]), .IN2(in2[46]), .Q(cout[46]) );
  NOR2X0 U26 ( .IN1(in3[46]), .IN2(in2[46]), .QN(n13) );
  NOR2X0 U27 ( .IN1(n13), .IN2(cout[46]), .QN(sumout[46]) );
  XOR2X1 U28 ( .IN1(in3[47]), .IN2(in2[47]), .Q(sumout[47]) );
  AND2X1 U29 ( .IN1(in3[12]), .IN2(in1[12]), .Q(cout[12]) );
  NOR2X0 U30 ( .IN1(in3[12]), .IN2(in1[12]), .QN(n14) );
  NOR2X0 U31 ( .IN1(n14), .IN2(cout[12]), .QN(sumout[12]) );
  AND2X1 U32 ( .IN1(in3[14]), .IN2(in1[14]), .Q(cout[14]) );
  NOR2X0 U33 ( .IN1(in3[14]), .IN2(in1[14]), .QN(n15) );
  NOR2X0 U34 ( .IN1(n15), .IN2(cout[14]), .QN(sumout[14]) );
  AND2X1 U35 ( .IN1(in3[16]), .IN2(in1[16]), .Q(cout[16]) );
  NOR2X0 U36 ( .IN1(in3[16]), .IN2(in1[16]), .QN(n16) );
  NOR2X0 U37 ( .IN1(n16), .IN2(cout[16]), .QN(sumout[16]) );
  AND2X1 U38 ( .IN1(in3[18]), .IN2(in1[18]), .Q(cout[18]) );
  NOR2X0 U39 ( .IN1(in3[18]), .IN2(in1[18]), .QN(n17) );
  NOR2X0 U40 ( .IN1(n17), .IN2(cout[18]), .QN(sumout[18]) );
  FADDX1 U41 ( .A(in1[19]), .B(in2[19]), .CI(in3[19]), .CO(cout[19]), .S(
        sumout[19]) );
  FADDX1 U42 ( .A(in1[20]), .B(in2[20]), .CI(in3[20]), .CO(cout[20]), .S(
        sumout[20]) );
  FADDX1 U43 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U44 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U45 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U46 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U47 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U48 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U49 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U50 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U51 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U52 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U53 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U54 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
  FADDX1 U55 ( .A(in1[33]), .B(in2[33]), .CI(in3[33]), .CO(cout[33]), .S(
        sumout[33]) );
  FADDX1 U56 ( .A(in1[34]), .B(in2[34]), .CI(in3[34]), .CO(cout[34]), .S(
        sumout[34]) );
  FADDX1 U57 ( .A(in1[35]), .B(in2[35]), .CI(in3[35]), .CO(cout[35]), .S(
        sumout[35]) );
  FADDX1 U58 ( .A(in1[36]), .B(in2[36]), .CI(in3[36]), .CO(cout[36]), .S(
        sumout[36]) );
  FADDX1 U59 ( .A(in1[37]), .B(in2[37]), .CI(in3[37]), .CO(cout[37]), .S(
        sumout[37]) );
  FADDX1 U60 ( .A(in1[38]), .B(in2[38]), .CI(in3[38]), .CO(cout[38]), .S(
        sumout[38]) );
  FADDX1 U61 ( .A(in1[39]), .B(in2[39]), .CI(in3[39]), .CO(cout[39]), .S(
        sumout[39]) );
  FADDX1 U62 ( .A(in1[40]), .B(in2[40]), .CI(in3[40]), .CO(cout[40]), .S(
        sumout[40]) );
  FADDX1 U63 ( .A(in1[41]), .B(in2[41]), .CI(in3[41]), .CO(cout[41]), .S(
        sumout[41]) );
  FADDX1 U64 ( .A(in1[42]), .B(in2[42]), .CI(in3[42]), .CO(cout[42]), .S(
        sumout[42]) );
endmodule


module csa51squ_53 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19;

  NBUFFX2 U1 ( .INP(in2[46]), .Z(sumout[46]) );
  NBUFFX2 U2 ( .INP(in2[45]), .Z(sumout[45]) );
  NBUFFX2 U3 ( .INP(in2[44]), .Z(sumout[44]) );
  NBUFFX2 U4 ( .INP(in2[43]), .Z(sumout[43]) );
  NBUFFX2 U5 ( .INP(in2[42]), .Z(sumout[42]) );
  NBUFFX2 U6 ( .INP(in2[41]), .Z(sumout[41]) );
  NBUFFX2 U7 ( .INP(in2[40]), .Z(sumout[40]) );
  NBUFFX2 U8 ( .INP(in2[39]), .Z(sumout[39]) );
  AND2X1 U9 ( .IN1(in2[7]), .IN2(in1[7]), .Q(cout[7]) );
  NOR2X0 U10 ( .IN1(in2[7]), .IN2(in1[7]), .QN(n9) );
  NOR2X0 U11 ( .IN1(n9), .IN2(cout[7]), .QN(sumout[7]) );
  AND2X1 U12 ( .IN1(in2[8]), .IN2(in1[8]), .Q(cout[8]) );
  NOR2X0 U13 ( .IN1(in2[8]), .IN2(in1[8]), .QN(n10) );
  NOR2X0 U14 ( .IN1(n10), .IN2(cout[8]), .QN(sumout[8]) );
  AND2X1 U15 ( .IN1(in2[9]), .IN2(in1[9]), .Q(cout[9]) );
  NOR2X0 U16 ( .IN1(in2[9]), .IN2(in1[9]), .QN(n11) );
  NOR2X0 U17 ( .IN1(n11), .IN2(cout[9]), .QN(sumout[9]) );
  AND2X1 U18 ( .IN1(in3[33]), .IN2(in2[33]), .Q(cout[33]) );
  NOR2X0 U19 ( .IN1(in3[33]), .IN2(in2[33]), .QN(n12) );
  NOR2X0 U20 ( .IN1(n12), .IN2(cout[33]), .QN(sumout[33]) );
  AND2X1 U21 ( .IN1(in3[34]), .IN2(in2[34]), .Q(cout[34]) );
  NOR2X0 U22 ( .IN1(in3[34]), .IN2(in2[34]), .QN(n13) );
  NOR2X0 U23 ( .IN1(n13), .IN2(cout[34]), .QN(sumout[34]) );
  AND2X1 U24 ( .IN1(in3[35]), .IN2(in2[35]), .Q(cout[35]) );
  NOR2X0 U25 ( .IN1(in3[35]), .IN2(in2[35]), .QN(n14) );
  NOR2X0 U26 ( .IN1(n14), .IN2(cout[35]), .QN(sumout[35]) );
  AND2X1 U27 ( .IN1(in3[36]), .IN2(in2[36]), .Q(cout[36]) );
  NOR2X0 U28 ( .IN1(in3[36]), .IN2(in2[36]), .QN(n15) );
  NOR2X0 U29 ( .IN1(n15), .IN2(cout[36]), .QN(sumout[36]) );
  AND2X1 U30 ( .IN1(in3[37]), .IN2(in2[37]), .Q(cout[37]) );
  NOR2X0 U31 ( .IN1(in3[37]), .IN2(in2[37]), .QN(n16) );
  NOR2X0 U32 ( .IN1(n16), .IN2(cout[37]), .QN(sumout[37]) );
  AND2X1 U33 ( .IN1(in3[38]), .IN2(in2[38]), .Q(cout[38]) );
  NOR2X0 U34 ( .IN1(in3[38]), .IN2(in2[38]), .QN(n17) );
  NOR2X0 U35 ( .IN1(n17), .IN2(cout[38]), .QN(sumout[38]) );
  AND2X1 U36 ( .IN1(in2[4]), .IN2(in1[4]), .Q(cout[4]) );
  AND2X1 U37 ( .IN1(in2[5]), .IN2(in1[5]), .Q(cout[5]) );
  NOR2X0 U38 ( .IN1(in2[5]), .IN2(in1[5]), .QN(n18) );
  NOR2X0 U39 ( .IN1(n18), .IN2(cout[5]), .QN(sumout[5]) );
  AND2X1 U40 ( .IN1(in2[6]), .IN2(in1[6]), .Q(cout[6]) );
  NOR2X0 U41 ( .IN1(in2[6]), .IN2(in1[6]), .QN(n19) );
  NOR2X0 U42 ( .IN1(n19), .IN2(cout[6]), .QN(sumout[6]) );
  FADDX1 U43 ( .A(in1[10]), .B(in2[10]), .CI(in3[10]), .CO(cout[10]), .S(
        sumout[10]) );
  FADDX1 U44 ( .A(in1[11]), .B(in2[11]), .CI(in3[11]), .CO(cout[11]), .S(
        sumout[11]) );
  FADDX1 U45 ( .A(in1[12]), .B(in2[12]), .CI(in3[12]), .CO(cout[12]), .S(
        sumout[12]) );
  FADDX1 U46 ( .A(in1[13]), .B(in2[13]), .CI(in3[13]), .CO(cout[13]), .S(
        sumout[13]) );
  FADDX1 U47 ( .A(in1[14]), .B(in2[14]), .CI(in3[14]), .CO(cout[14]), .S(
        sumout[14]) );
  FADDX1 U48 ( .A(in1[15]), .B(in2[15]), .CI(in3[15]), .CO(cout[15]), .S(
        sumout[15]) );
  FADDX1 U49 ( .A(in1[16]), .B(in2[16]), .CI(in3[16]), .CO(cout[16]), .S(
        sumout[16]) );
  FADDX1 U50 ( .A(in1[17]), .B(in2[17]), .CI(in3[17]), .CO(cout[17]), .S(
        sumout[17]) );
  FADDX1 U51 ( .A(in1[18]), .B(in2[18]), .CI(in3[18]), .CO(cout[18]), .S(
        sumout[18]) );
  FADDX1 U52 ( .A(in1[19]), .B(in2[19]), .CI(in3[19]), .CO(cout[19]), .S(
        sumout[19]) );
  FADDX1 U53 ( .A(in1[20]), .B(in2[20]), .CI(in3[20]), .CO(cout[20]), .S(
        sumout[20]) );
  FADDX1 U54 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U55 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U56 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U57 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U58 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U59 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U60 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U61 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U62 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U63 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U64 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U65 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
endmodule


module csa51squ_54 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n7, n8, n9, n10, n11, n12, n13;

  NBUFFX2 U1 ( .INP(in1[12]), .Z(sumout[12]) );
  NBUFFX2 U2 ( .INP(in1[13]), .Z(sumout[13]) );
  NBUFFX2 U3 ( .INP(in1[14]), .Z(sumout[14]) );
  NBUFFX2 U4 ( .INP(in1[15]), .Z(sumout[15]) );
  NBUFFX2 U5 ( .INP(in1[16]), .Z(sumout[16]) );
  NBUFFX2 U6 ( .INP(in1[17]), .Z(sumout[17]) );
  AND2X1 U7 ( .IN1(in3[19]), .IN2(in1[19]), .Q(cout[19]) );
  NOR2X0 U8 ( .IN1(in3[19]), .IN2(in1[19]), .QN(n7) );
  NOR2X0 U9 ( .IN1(n7), .IN2(cout[19]), .QN(sumout[19]) );
  AND2X1 U10 ( .IN1(in3[44]), .IN2(in2[44]), .Q(cout[44]) );
  NOR2X0 U11 ( .IN1(in3[44]), .IN2(in2[44]), .QN(n8) );
  NOR2X0 U12 ( .IN1(n8), .IN2(cout[44]), .QN(sumout[44]) );
  AND2X1 U13 ( .IN1(in3[45]), .IN2(in2[45]), .Q(cout[45]) );
  NOR2X0 U14 ( .IN1(in3[45]), .IN2(in2[45]), .QN(n9) );
  NOR2X0 U15 ( .IN1(n9), .IN2(cout[45]), .QN(sumout[45]) );
  AND2X1 U16 ( .IN1(in3[46]), .IN2(in2[46]), .Q(cout[46]) );
  NOR2X0 U17 ( .IN1(in3[46]), .IN2(in2[46]), .QN(n10) );
  NOR2X0 U18 ( .IN1(n10), .IN2(cout[46]), .QN(sumout[46]) );
  XOR2X1 U19 ( .IN1(in3[47]), .IN2(in2[47]), .Q(sumout[47]) );
  AND2X1 U20 ( .IN1(in3[18]), .IN2(in1[18]), .Q(cout[18]) );
  NOR2X0 U21 ( .IN1(in3[18]), .IN2(in1[18]), .QN(n11) );
  NOR2X0 U22 ( .IN1(n11), .IN2(cout[18]), .QN(sumout[18]) );
  AND2X1 U23 ( .IN1(in3[20]), .IN2(in1[20]), .Q(cout[20]) );
  NOR2X0 U24 ( .IN1(in3[20]), .IN2(in1[20]), .QN(n12) );
  NOR2X0 U25 ( .IN1(n12), .IN2(cout[20]), .QN(sumout[20]) );
  INVX0 U26 ( .INP(in1[42]), .ZN(n13) );
  FADDX1 U27 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U28 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U29 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U30 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U31 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U32 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U33 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U34 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U35 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U36 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U37 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U38 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
  FADDX1 U39 ( .A(in1[33]), .B(in2[33]), .CI(in3[33]), .CO(cout[33]), .S(
        sumout[33]) );
  FADDX1 U40 ( .A(in1[34]), .B(in2[34]), .CI(in3[34]), .CO(cout[34]), .S(
        sumout[34]) );
  FADDX1 U41 ( .A(in1[35]), .B(in2[35]), .CI(in3[35]), .CO(cout[35]), .S(
        sumout[35]) );
  FADDX1 U42 ( .A(in1[36]), .B(in2[36]), .CI(in3[36]), .CO(cout[36]), .S(
        sumout[36]) );
  FADDX1 U43 ( .A(in1[37]), .B(in2[37]), .CI(in3[37]), .CO(cout[37]), .S(
        sumout[37]) );
  FADDX1 U44 ( .A(in1[38]), .B(in2[38]), .CI(in3[38]), .CO(cout[38]), .S(
        sumout[38]) );
  FADDX1 U45 ( .A(in1[39]), .B(in2[39]), .CI(in3[39]), .CO(cout[39]), .S(
        sumout[39]) );
  FADDX1 U46 ( .A(in1[40]), .B(in2[40]), .CI(in3[40]), .CO(cout[40]), .S(
        sumout[40]) );
  FADDX1 U47 ( .A(in1[41]), .B(in2[41]), .CI(in3[41]), .CO(cout[41]), .S(
        sumout[41]) );
  FADDX1 U48 ( .A(in1[42]), .B(in2[42]), .CI(in3[42]), .CO(cout[42]), .S(
        sumout[42]) );
  FADDX1 U49 ( .A(in2[43]), .B(in3[43]), .CI(n13), .CO(cout[43]), .S(
        sumout[43]) );
endmodule


module csa51squ_55 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n9, n10, n11, n12, n13, n14, n15;

  NBUFFX2 U1 ( .INP(in2[6]), .Z(sumout[6]) );
  NBUFFX2 U2 ( .INP(in2[7]), .Z(sumout[7]) );
  NBUFFX2 U3 ( .INP(in2[8]), .Z(sumout[8]) );
  NBUFFX2 U4 ( .INP(in3[42]), .Z(sumout[42]) );
  NBUFFX2 U5 ( .INP(in3[41]), .Z(sumout[41]) );
  NBUFFX2 U6 ( .INP(in3[39]), .Z(sumout[39]) );
  NBUFFX2 U7 ( .INP(in3[38]), .Z(sumout[38]) );
  NBUFFX2 U8 ( .INP(in3[40]), .Z(sumout[40]) );
  AND2X1 U9 ( .IN1(in2[13]), .IN2(in1[13]), .Q(cout[13]) );
  NOR2X0 U10 ( .IN1(in2[13]), .IN2(in1[13]), .QN(n9) );
  NOR2X0 U11 ( .IN1(n9), .IN2(cout[13]), .QN(sumout[13]) );
  AND2X1 U12 ( .IN1(in2[37]), .IN2(in3[37]), .Q(cout[37]) );
  INVX0 U13 ( .INP(in2[37]), .ZN(n15) );
  MUX21X1 U14 ( .IN1(in2[37]), .IN2(n15), .S(in3[37]), .Q(sumout[37]) );
  AND2X1 U15 ( .IN1(in2[9]), .IN2(in1[9]), .Q(cout[9]) );
  NOR2X0 U16 ( .IN1(in2[9]), .IN2(in1[9]), .QN(n10) );
  NOR2X0 U17 ( .IN1(n10), .IN2(cout[9]), .QN(sumout[9]) );
  AND2X1 U18 ( .IN1(in2[10]), .IN2(in1[10]), .Q(cout[10]) );
  NOR2X0 U19 ( .IN1(in2[10]), .IN2(in1[10]), .QN(n11) );
  NOR2X0 U20 ( .IN1(n11), .IN2(cout[10]), .QN(sumout[10]) );
  AND2X1 U21 ( .IN1(in2[11]), .IN2(in1[11]), .Q(cout[11]) );
  NOR2X0 U22 ( .IN1(in2[11]), .IN2(in1[11]), .QN(n12) );
  NOR2X0 U23 ( .IN1(n12), .IN2(cout[11]), .QN(sumout[11]) );
  AND2X1 U24 ( .IN1(in2[12]), .IN2(in1[12]), .Q(cout[12]) );
  NOR2X0 U25 ( .IN1(in2[12]), .IN2(in1[12]), .QN(n13) );
  NOR2X0 U26 ( .IN1(n13), .IN2(cout[12]), .QN(sumout[12]) );
  AND2X1 U27 ( .IN1(in2[14]), .IN2(in1[14]), .Q(cout[14]) );
  NOR2X0 U28 ( .IN1(in2[14]), .IN2(in1[14]), .QN(n14) );
  NOR2X0 U29 ( .IN1(n14), .IN2(cout[14]), .QN(sumout[14]) );
  FADDX1 U30 ( .A(in1[15]), .B(in2[15]), .CI(in3[15]), .CO(cout[15]), .S(
        sumout[15]) );
  FADDX1 U31 ( .A(in1[16]), .B(in2[16]), .CI(in3[16]), .CO(cout[16]), .S(
        sumout[16]) );
  FADDX1 U32 ( .A(in1[17]), .B(in2[17]), .CI(in3[17]), .CO(cout[17]), .S(
        sumout[17]) );
  FADDX1 U33 ( .A(in1[18]), .B(in2[18]), .CI(in3[18]), .CO(cout[18]), .S(
        sumout[18]) );
  FADDX1 U34 ( .A(in1[19]), .B(in2[19]), .CI(in3[19]), .CO(cout[19]), .S(
        sumout[19]) );
  FADDX1 U35 ( .A(in1[20]), .B(in2[20]), .CI(in3[20]), .CO(cout[20]), .S(
        sumout[20]) );
  FADDX1 U36 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U37 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U38 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U39 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U40 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U41 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U42 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U43 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U44 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U45 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U46 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U47 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
  FADDX1 U48 ( .A(in1[33]), .B(in2[33]), .CI(in3[33]), .CO(cout[33]), .S(
        sumout[33]) );
  FADDX1 U49 ( .A(in1[34]), .B(in2[34]), .CI(in3[34]), .CO(cout[34]), .S(
        sumout[34]) );
  FADDX1 U50 ( .A(in1[35]), .B(in2[35]), .CI(in3[35]), .CO(cout[35]), .S(
        sumout[35]) );
  FADDX1 U51 ( .A(in1[36]), .B(in3[36]), .CI(n15), .CO(cout[36]), .S(
        sumout[36]) );
endmodule


module csa51squ_56 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36;

  NBUFFX2 U1 ( .INP(in3[46]), .Z(sumout[46]) );
  NBUFFX2 U2 ( .INP(in3[45]), .Z(sumout[45]) );
  NBUFFX2 U3 ( .INP(in3[44]), .Z(sumout[44]) );
  NBUFFX2 U4 ( .INP(in3[43]), .Z(sumout[43]) );
  NBUFFX2 U5 ( .INP(in3[42]), .Z(sumout[42]) );
  NBUFFX2 U6 ( .INP(in3[37]), .Z(sumout[37]) );
  NBUFFX2 U7 ( .INP(in3[36]), .Z(sumout[36]) );
  NBUFFX2 U8 ( .INP(in3[35]), .Z(sumout[35]) );
  NBUFFX2 U9 ( .INP(in3[34]), .Z(sumout[34]) );
  NBUFFX2 U10 ( .INP(in3[33]), .Z(sumout[33]) );
  NBUFFX2 U11 ( .INP(in3[32]), .Z(sumout[32]) );
  NBUFFX2 U12 ( .INP(in3[41]), .Z(sumout[41]) );
  NBUFFX2 U13 ( .INP(in3[40]), .Z(sumout[40]) );
  NBUFFX2 U14 ( .INP(in3[39]), .Z(sumout[39]) );
  NBUFFX2 U15 ( .INP(in3[38]), .Z(sumout[38]) );
  AND2X1 U16 ( .IN1(in2[31]), .IN2(in3[31]), .Q(cout[31]) );
  INVX0 U17 ( .INP(in2[31]), .ZN(n36) );
  MUX21X1 U18 ( .IN1(in2[31]), .IN2(n36), .S(in3[31]), .Q(sumout[31]) );
  AND2X1 U19 ( .IN1(in2[3]), .IN2(in1[3]), .Q(cout[3]) );
  AND2X1 U20 ( .IN1(in2[4]), .IN2(in1[4]), .Q(cout[4]) );
  NOR2X0 U21 ( .IN1(in2[4]), .IN2(in1[4]), .QN(n16) );
  NOR2X0 U22 ( .IN1(n16), .IN2(cout[4]), .QN(sumout[4]) );
  AND2X1 U23 ( .IN1(in2[5]), .IN2(in1[5]), .Q(cout[5]) );
  NOR2X0 U24 ( .IN1(in2[5]), .IN2(in1[5]), .QN(n17) );
  NOR2X0 U25 ( .IN1(n17), .IN2(cout[5]), .QN(sumout[5]) );
  AND2X1 U26 ( .IN1(in2[6]), .IN2(in1[6]), .Q(cout[6]) );
  NOR2X0 U27 ( .IN1(in2[6]), .IN2(in1[6]), .QN(n18) );
  NOR2X0 U28 ( .IN1(n18), .IN2(cout[6]), .QN(sumout[6]) );
  AND2X1 U29 ( .IN1(in2[7]), .IN2(in1[7]), .Q(cout[7]) );
  NOR2X0 U30 ( .IN1(in2[7]), .IN2(in1[7]), .QN(n19) );
  NOR2X0 U31 ( .IN1(n19), .IN2(cout[7]), .QN(sumout[7]) );
  AND2X1 U32 ( .IN1(in2[8]), .IN2(in1[8]), .Q(cout[8]) );
  NOR2X0 U33 ( .IN1(in2[8]), .IN2(in1[8]), .QN(n20) );
  NOR2X0 U34 ( .IN1(n20), .IN2(cout[8]), .QN(sumout[8]) );
  AND2X1 U35 ( .IN1(in2[9]), .IN2(in1[9]), .Q(cout[9]) );
  NOR2X0 U36 ( .IN1(in2[9]), .IN2(in1[9]), .QN(n21) );
  NOR2X0 U37 ( .IN1(n21), .IN2(cout[9]), .QN(sumout[9]) );
  AND2X1 U38 ( .IN1(in2[10]), .IN2(in1[10]), .Q(cout[10]) );
  NOR2X0 U39 ( .IN1(in2[10]), .IN2(in1[10]), .QN(n22) );
  NOR2X0 U40 ( .IN1(n22), .IN2(cout[10]), .QN(sumout[10]) );
  AND2X1 U41 ( .IN1(in2[11]), .IN2(in1[11]), .Q(cout[11]) );
  NOR2X0 U42 ( .IN1(in2[11]), .IN2(in1[11]), .QN(n23) );
  NOR2X0 U43 ( .IN1(n23), .IN2(cout[11]), .QN(sumout[11]) );
  AND2X1 U44 ( .IN1(in2[12]), .IN2(in1[12]), .Q(cout[12]) );
  NOR2X0 U45 ( .IN1(in2[12]), .IN2(in1[12]), .QN(n24) );
  NOR2X0 U46 ( .IN1(n24), .IN2(cout[12]), .QN(sumout[12]) );
  AND2X1 U47 ( .IN1(in2[13]), .IN2(in1[13]), .Q(cout[13]) );
  NOR2X0 U48 ( .IN1(in2[13]), .IN2(in1[13]), .QN(n25) );
  NOR2X0 U49 ( .IN1(n25), .IN2(cout[13]), .QN(sumout[13]) );
  AND2X1 U50 ( .IN1(in2[14]), .IN2(in1[14]), .Q(cout[14]) );
  NOR2X0 U51 ( .IN1(in2[14]), .IN2(in1[14]), .QN(n26) );
  NOR2X0 U52 ( .IN1(n26), .IN2(cout[14]), .QN(sumout[14]) );
  AND2X1 U53 ( .IN1(in2[15]), .IN2(in1[15]), .Q(cout[15]) );
  NOR2X0 U54 ( .IN1(in2[15]), .IN2(in1[15]), .QN(n27) );
  NOR2X0 U55 ( .IN1(n27), .IN2(cout[15]), .QN(sumout[15]) );
  AND2X1 U56 ( .IN1(in2[16]), .IN2(in1[16]), .Q(cout[16]) );
  NOR2X0 U57 ( .IN1(in2[16]), .IN2(in1[16]), .QN(n28) );
  NOR2X0 U58 ( .IN1(n28), .IN2(cout[16]), .QN(sumout[16]) );
  AND2X1 U59 ( .IN1(in2[17]), .IN2(in1[17]), .Q(cout[17]) );
  NOR2X0 U60 ( .IN1(in2[17]), .IN2(in1[17]), .QN(n29) );
  NOR2X0 U61 ( .IN1(n29), .IN2(cout[17]), .QN(sumout[17]) );
  AND2X1 U62 ( .IN1(in2[18]), .IN2(in1[18]), .Q(cout[18]) );
  NOR2X0 U63 ( .IN1(in2[18]), .IN2(in1[18]), .QN(n30) );
  NOR2X0 U64 ( .IN1(n30), .IN2(cout[18]), .QN(sumout[18]) );
  AND2X1 U65 ( .IN1(in2[19]), .IN2(in1[19]), .Q(cout[19]) );
  NOR2X0 U66 ( .IN1(in2[19]), .IN2(in1[19]), .QN(n31) );
  NOR2X0 U67 ( .IN1(n31), .IN2(cout[19]), .QN(sumout[19]) );
  AND2X1 U68 ( .IN1(in2[20]), .IN2(in1[20]), .Q(cout[20]) );
  NOR2X0 U69 ( .IN1(in2[20]), .IN2(in1[20]), .QN(n32) );
  NOR2X0 U70 ( .IN1(n32), .IN2(cout[20]), .QN(sumout[20]) );
  AND2X1 U71 ( .IN1(in2[21]), .IN2(in1[21]), .Q(cout[21]) );
  NOR2X0 U72 ( .IN1(in2[21]), .IN2(in1[21]), .QN(n33) );
  NOR2X0 U73 ( .IN1(n33), .IN2(cout[21]), .QN(sumout[21]) );
  AND2X1 U74 ( .IN1(in2[22]), .IN2(in1[22]), .Q(cout[22]) );
  NOR2X0 U75 ( .IN1(in2[22]), .IN2(in1[22]), .QN(n34) );
  NOR2X0 U76 ( .IN1(n34), .IN2(cout[22]), .QN(sumout[22]) );
  AND2X1 U77 ( .IN1(in2[23]), .IN2(in1[23]), .Q(cout[23]) );
  NOR2X0 U78 ( .IN1(in2[23]), .IN2(in1[23]), .QN(n35) );
  NOR2X0 U79 ( .IN1(n35), .IN2(cout[23]), .QN(sumout[23]) );
  FADDX1 U80 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U81 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U82 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U83 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U84 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U85 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U86 ( .A(in1[30]), .B(in3[30]), .CI(n36), .CO(cout[30]), .S(
        sumout[30]) );
endmodule


module csa51squ_57 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n3, n4, n5, n6, n7;

  NBUFFX2 U1 ( .INP(in1[18]), .Z(sumout[18]) );
  NBUFFX2 U2 ( .INP(in1[19]), .Z(sumout[19]) );
  AND2X1 U3 ( .IN1(in2[20]), .IN2(in1[20]), .Q(cout[20]) );
  NOR2X0 U4 ( .IN1(in2[20]), .IN2(in1[20]), .QN(n3) );
  NOR2X0 U5 ( .IN1(n3), .IN2(cout[20]), .QN(sumout[20]) );
  AND2X1 U6 ( .IN1(in2[21]), .IN2(in1[21]), .Q(cout[21]) );
  NOR2X0 U7 ( .IN1(in2[21]), .IN2(in1[21]), .QN(n4) );
  NOR2X0 U8 ( .IN1(n4), .IN2(cout[21]), .QN(sumout[21]) );
  AND2X1 U9 ( .IN1(in2[46]), .IN2(in3[46]), .Q(cout[46]) );
  NOR2X0 U10 ( .IN1(in2[46]), .IN2(in3[46]), .QN(n5) );
  NOR2X0 U11 ( .IN1(n5), .IN2(cout[46]), .QN(sumout[46]) );
  INVX0 U12 ( .INP(in2[46]), .ZN(n6) );
  MUX21X1 U13 ( .IN1(n6), .IN2(in2[46]), .S(in3[47]), .Q(sumout[47]) );
  INVX0 U14 ( .INP(in1[44]), .ZN(n7) );
  FADDX1 U15 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U16 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U17 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U18 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U19 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U20 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U21 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U22 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U23 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U24 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U25 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
  FADDX1 U26 ( .A(in1[33]), .B(in2[33]), .CI(in3[33]), .CO(cout[33]), .S(
        sumout[33]) );
  FADDX1 U27 ( .A(in1[34]), .B(in2[34]), .CI(in3[34]), .CO(cout[34]), .S(
        sumout[34]) );
  FADDX1 U28 ( .A(in1[35]), .B(in2[35]), .CI(in3[35]), .CO(cout[35]), .S(
        sumout[35]) );
  FADDX1 U29 ( .A(in1[36]), .B(in2[36]), .CI(in3[36]), .CO(cout[36]), .S(
        sumout[36]) );
  FADDX1 U30 ( .A(in1[37]), .B(in2[37]), .CI(in3[37]), .CO(cout[37]), .S(
        sumout[37]) );
  FADDX1 U31 ( .A(in1[38]), .B(in2[38]), .CI(in3[38]), .CO(cout[38]), .S(
        sumout[38]) );
  FADDX1 U32 ( .A(in1[39]), .B(in2[39]), .CI(in3[39]), .CO(cout[39]), .S(
        sumout[39]) );
  FADDX1 U33 ( .A(in1[40]), .B(in2[40]), .CI(in3[40]), .CO(cout[40]), .S(
        sumout[40]) );
  FADDX1 U34 ( .A(in1[41]), .B(in2[41]), .CI(in3[41]), .CO(cout[41]), .S(
        sumout[41]) );
  FADDX1 U35 ( .A(in1[42]), .B(in2[42]), .CI(in3[42]), .CO(cout[42]), .S(
        sumout[42]) );
  FADDX1 U36 ( .A(in1[43]), .B(in2[43]), .CI(in3[43]), .CO(cout[43]), .S(
        sumout[43]) );
  FADDX1 U37 ( .A(in1[44]), .B(in2[44]), .CI(in3[44]), .CO(cout[44]), .S(
        sumout[44]) );
  FADDX1 U38 ( .A(in2[45]), .B(in3[45]), .CI(n7), .CO(cout[45]), .S(sumout[45]) );
endmodule


module csa51squ_58 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n4, n5, n6, n7, n8;

  NBUFFX2 U1 ( .INP(in1[12]), .Z(sumout[12]) );
  NBUFFX2 U2 ( .INP(in1[13]), .Z(sumout[13]) );
  NBUFFX2 U3 ( .INP(in3[42]), .Z(sumout[42]) );
  AND2X1 U4 ( .IN1(in2[14]), .IN2(in1[14]), .Q(cout[14]) );
  NOR2X0 U5 ( .IN1(in2[14]), .IN2(in1[14]), .QN(n4) );
  NOR2X0 U6 ( .IN1(n4), .IN2(cout[14]), .QN(sumout[14]) );
  AND2X1 U7 ( .IN1(in2[15]), .IN2(in1[15]), .Q(cout[15]) );
  NOR2X0 U8 ( .IN1(in2[15]), .IN2(in1[15]), .QN(n5) );
  NOR2X0 U9 ( .IN1(n5), .IN2(cout[15]), .QN(sumout[15]) );
  AND2X1 U10 ( .IN1(in2[40]), .IN2(in3[40]), .Q(cout[40]) );
  NOR2X0 U11 ( .IN1(in2[40]), .IN2(in3[40]), .QN(n6) );
  NOR2X0 U12 ( .IN1(n6), .IN2(cout[40]), .QN(sumout[40]) );
  INVX0 U13 ( .INP(in3[41]), .ZN(n7) );
  NOR2X0 U14 ( .IN1(in2[40]), .IN2(n7), .QN(cout[41]) );
  MUX21X1 U15 ( .IN1(n7), .IN2(in3[41]), .S(in2[40]), .Q(sumout[41]) );
  INVX0 U16 ( .INP(in1[38]), .ZN(n8) );
  FADDX1 U17 ( .A(in1[16]), .B(in2[16]), .CI(in3[16]), .CO(cout[16]), .S(
        sumout[16]) );
  FADDX1 U18 ( .A(in1[17]), .B(in2[17]), .CI(in3[17]), .CO(cout[17]), .S(
        sumout[17]) );
  FADDX1 U19 ( .A(in1[18]), .B(in2[18]), .CI(in3[18]), .CO(cout[18]), .S(
        sumout[18]) );
  FADDX1 U20 ( .A(in1[19]), .B(in2[19]), .CI(in3[19]), .CO(cout[19]), .S(
        sumout[19]) );
  FADDX1 U21 ( .A(in1[20]), .B(in2[20]), .CI(in3[20]), .CO(cout[20]), .S(
        sumout[20]) );
  FADDX1 U22 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U23 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U24 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U25 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U26 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U27 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U28 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U29 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U30 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U31 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U32 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U33 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
  FADDX1 U34 ( .A(in1[33]), .B(in2[33]), .CI(in3[33]), .CO(cout[33]), .S(
        sumout[33]) );
  FADDX1 U35 ( .A(in1[34]), .B(in2[34]), .CI(in3[34]), .CO(cout[34]), .S(
        sumout[34]) );
  FADDX1 U36 ( .A(in1[35]), .B(in2[35]), .CI(in3[35]), .CO(cout[35]), .S(
        sumout[35]) );
  FADDX1 U37 ( .A(in1[36]), .B(in2[36]), .CI(in3[36]), .CO(cout[36]), .S(
        sumout[36]) );
  FADDX1 U38 ( .A(in1[37]), .B(in2[37]), .CI(in3[37]), .CO(cout[37]), .S(
        sumout[37]) );
  FADDX1 U39 ( .A(in1[38]), .B(in2[38]), .CI(in3[38]), .CO(cout[38]), .S(
        sumout[38]) );
  FADDX1 U40 ( .A(in2[39]), .B(in3[39]), .CI(n8), .CO(cout[39]), .S(sumout[39]) );
endmodule


module csa51squ_59 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n4, n5, n6, n7, n8;

  NBUFFX2 U1 ( .INP(in1[6]), .Z(sumout[6]) );
  NBUFFX2 U2 ( .INP(in1[7]), .Z(sumout[7]) );
  NBUFFX2 U3 ( .INP(in3[37]), .Z(sumout[37]) );
  AND2X1 U4 ( .IN1(in2[8]), .IN2(in1[8]), .Q(cout[8]) );
  NOR2X0 U5 ( .IN1(in2[8]), .IN2(in1[8]), .QN(n4) );
  NOR2X0 U6 ( .IN1(n4), .IN2(cout[8]), .QN(sumout[8]) );
  AND2X1 U7 ( .IN1(in2[9]), .IN2(in1[9]), .Q(cout[9]) );
  NOR2X0 U8 ( .IN1(in2[9]), .IN2(in1[9]), .QN(n5) );
  NOR2X0 U9 ( .IN1(n5), .IN2(cout[9]), .QN(sumout[9]) );
  AND2X1 U10 ( .IN1(in2[34]), .IN2(in3[34]), .Q(cout[34]) );
  NOR2X0 U11 ( .IN1(in2[34]), .IN2(in3[34]), .QN(n6) );
  NOR2X0 U12 ( .IN1(n6), .IN2(cout[34]), .QN(sumout[34]) );
  INVX0 U13 ( .INP(in3[35]), .ZN(n7) );
  NOR2X0 U14 ( .IN1(in2[34]), .IN2(n7), .QN(cout[35]) );
  MUX21X1 U15 ( .IN1(n7), .IN2(in3[35]), .S(in2[34]), .Q(sumout[35]) );
  INVX0 U16 ( .INP(in1[32]), .ZN(n8) );
  FADDX1 U17 ( .A(in1[10]), .B(in2[10]), .CI(in3[10]), .CO(cout[10]), .S(
        sumout[10]) );
  FADDX1 U18 ( .A(in1[11]), .B(in2[11]), .CI(in3[11]), .CO(cout[11]), .S(
        sumout[11]) );
  FADDX1 U19 ( .A(in1[12]), .B(in2[12]), .CI(in3[12]), .CO(cout[12]), .S(
        sumout[12]) );
  FADDX1 U20 ( .A(in1[13]), .B(in2[13]), .CI(in3[13]), .CO(cout[13]), .S(
        sumout[13]) );
  FADDX1 U21 ( .A(in1[14]), .B(in2[14]), .CI(in3[14]), .CO(cout[14]), .S(
        sumout[14]) );
  FADDX1 U22 ( .A(in1[15]), .B(in2[15]), .CI(in3[15]), .CO(cout[15]), .S(
        sumout[15]) );
  FADDX1 U23 ( .A(in1[16]), .B(in2[16]), .CI(in3[16]), .CO(cout[16]), .S(
        sumout[16]) );
  FADDX1 U24 ( .A(in1[17]), .B(in2[17]), .CI(in3[17]), .CO(cout[17]), .S(
        sumout[17]) );
  FADDX1 U25 ( .A(in1[18]), .B(in2[18]), .CI(in3[18]), .CO(cout[18]), .S(
        sumout[18]) );
  FADDX1 U26 ( .A(in1[19]), .B(in2[19]), .CI(in3[19]), .CO(cout[19]), .S(
        sumout[19]) );
  FADDX1 U27 ( .A(in1[20]), .B(in2[20]), .CI(in3[20]), .CO(cout[20]), .S(
        sumout[20]) );
  FADDX1 U28 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U29 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U30 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U31 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U32 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U33 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U34 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U35 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U36 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U37 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U38 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U39 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
  FADDX1 U40 ( .A(in2[33]), .B(in3[33]), .CI(n8), .CO(cout[33]), .S(sumout[33]) );
endmodule


module csa51squ_60 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n2, n3, n4, n5;

  NBUFFX2 U1 ( .INP(in3[31]), .Z(sumout[31]) );
  AND2X1 U2 ( .IN1(in2[2]), .IN2(in1[2]), .Q(cout[2]) );
  AND2X1 U3 ( .IN1(in2[3]), .IN2(in1[3]), .Q(cout[3]) );
  NOR2X0 U4 ( .IN1(in2[3]), .IN2(in1[3]), .QN(n2) );
  NOR2X0 U5 ( .IN1(n2), .IN2(cout[3]), .QN(sumout[3]) );
  AND2X1 U6 ( .IN1(in2[28]), .IN2(in3[28]), .Q(cout[28]) );
  NOR2X0 U7 ( .IN1(in2[28]), .IN2(in3[28]), .QN(n3) );
  NOR2X0 U8 ( .IN1(n3), .IN2(cout[28]), .QN(sumout[28]) );
  INVX0 U9 ( .INP(in3[29]), .ZN(n4) );
  NOR2X0 U10 ( .IN1(in2[28]), .IN2(n4), .QN(cout[29]) );
  MUX21X1 U11 ( .IN1(n4), .IN2(in3[29]), .S(in2[28]), .Q(sumout[29]) );
  INVX0 U12 ( .INP(in1[26]), .ZN(n5) );
  FADDX1 U13 ( .A(in1[10]), .B(in2[10]), .CI(in3[10]), .CO(cout[10]), .S(
        sumout[10]) );
  FADDX1 U14 ( .A(in1[11]), .B(in2[11]), .CI(in3[11]), .CO(cout[11]), .S(
        sumout[11]) );
  FADDX1 U15 ( .A(in1[12]), .B(in2[12]), .CI(in3[12]), .CO(cout[12]), .S(
        sumout[12]) );
  FADDX1 U16 ( .A(in1[13]), .B(in2[13]), .CI(in3[13]), .CO(cout[13]), .S(
        sumout[13]) );
  FADDX1 U17 ( .A(in1[14]), .B(in2[14]), .CI(in3[14]), .CO(cout[14]), .S(
        sumout[14]) );
  FADDX1 U18 ( .A(in1[15]), .B(in2[15]), .CI(in3[15]), .CO(cout[15]), .S(
        sumout[15]) );
  FADDX1 U19 ( .A(in1[16]), .B(in2[16]), .CI(in3[16]), .CO(cout[16]), .S(
        sumout[16]) );
  FADDX1 U20 ( .A(in1[17]), .B(in2[17]), .CI(in3[17]), .CO(cout[17]), .S(
        sumout[17]) );
  FADDX1 U21 ( .A(in1[18]), .B(in2[18]), .CI(in3[18]), .CO(cout[18]), .S(
        sumout[18]) );
  FADDX1 U22 ( .A(in1[19]), .B(in2[19]), .CI(in3[19]), .CO(cout[19]), .S(
        sumout[19]) );
  FADDX1 U23 ( .A(in1[20]), .B(in2[20]), .CI(in3[20]), .CO(cout[20]), .S(
        sumout[20]) );
  FADDX1 U24 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U25 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U26 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U27 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U28 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U29 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U30 ( .A(in2[27]), .B(in3[27]), .CI(n5), .CO(cout[27]), .S(sumout[27]) );
  FADDX1 U31 ( .A(in1[4]), .B(in2[4]), .CI(in3[4]), .CO(cout[4]), .S(sumout[4]) );
  FADDX1 U32 ( .A(in1[5]), .B(in2[5]), .CI(in3[5]), .CO(cout[5]), .S(sumout[5]) );
  FADDX1 U33 ( .A(in1[6]), .B(in2[6]), .CI(in3[6]), .CO(cout[6]), .S(sumout[6]) );
  FADDX1 U34 ( .A(in1[7]), .B(in2[7]), .CI(in3[7]), .CO(cout[7]), .S(sumout[7]) );
  FADDX1 U35 ( .A(in1[8]), .B(in2[8]), .CI(in3[8]), .CO(cout[8]), .S(sumout[8]) );
  FADDX1 U36 ( .A(in1[9]), .B(in2[9]), .CI(in3[9]), .CO(cout[9]), .S(sumout[9]) );
endmodule


module booth27_53 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;


  NBUFFX2 U3 ( .INP(in2[22]), .Z(out1[22]) );
  NBUFFX2 U4 ( .INP(in2[21]), .Z(out1[21]) );
  NBUFFX2 U5 ( .INP(in2[20]), .Z(out1[20]) );
  NBUFFX2 U6 ( .INP(in2[0]), .Z(out1[0]) );
  NBUFFX2 U7 ( .INP(in2[19]), .Z(out1[19]) );
  NBUFFX2 U8 ( .INP(in2[18]), .Z(out1[18]) );
  NBUFFX2 U9 ( .INP(in2[2]), .Z(out1[2]) );
  NBUFFX2 U10 ( .INP(in2[1]), .Z(out1[1]) );
  NBUFFX2 U11 ( .INP(in2[4]), .Z(out1[4]) );
  NBUFFX2 U12 ( .INP(in2[3]), .Z(out1[3]) );
  NBUFFX2 U13 ( .INP(in2[13]), .Z(out1[13]) );
  NBUFFX2 U14 ( .INP(in2[12]), .Z(out1[12]) );
  NBUFFX2 U15 ( .INP(in2[11]), .Z(out1[11]) );
  NBUFFX2 U16 ( .INP(in2[10]), .Z(out1[10]) );
  NBUFFX2 U17 ( .INP(in2[9]), .Z(out1[9]) );
  NBUFFX2 U18 ( .INP(in2[8]), .Z(out1[8]) );
  NBUFFX2 U19 ( .INP(in2[7]), .Z(out1[7]) );
  NBUFFX2 U20 ( .INP(in2[6]), .Z(out1[6]) );
  NBUFFX2 U21 ( .INP(in2[5]), .Z(out1[5]) );
  NBUFFX2 U22 ( .INP(in2[17]), .Z(out1[17]) );
  NBUFFX2 U23 ( .INP(in2[16]), .Z(out1[16]) );
  NBUFFX2 U24 ( .INP(in2[15]), .Z(out1[15]) );
  NBUFFX2 U25 ( .INP(in2[14]), .Z(out1[14]) );
endmodule


module booth27_54 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76;

  NAND2X0 U3 ( .IN1(n1), .IN2(n2), .QN(n8) );
  NAND2X0 U4 ( .IN1(n71), .IN2(in2[0]), .QN(n15) );
  NAND2X0 U5 ( .IN1(n19), .IN2(in2[5]), .QN(n20) );
  NAND2X0 U6 ( .IN1(n25), .IN2(in2[7]), .QN(n26) );
  NAND2X0 U7 ( .IN1(n31), .IN2(in2[9]), .QN(n32) );
  NAND2X0 U8 ( .IN1(n37), .IN2(in2[11]), .QN(n38) );
  NAND2X0 U9 ( .IN1(n43), .IN2(in2[13]), .QN(n44) );
  NAND2X0 U10 ( .IN1(n46), .IN2(in2[14]), .QN(n47) );
  NAND2X0 U11 ( .IN1(n49), .IN2(in2[15]), .QN(n50) );
  NAND2X0 U12 ( .IN1(n52), .IN2(in2[16]), .QN(n53) );
  NAND2X0 U13 ( .IN1(n55), .IN2(in2[17]), .QN(n56) );
  NAND2X0 U14 ( .IN1(n7), .IN2(n15), .QN(out1[1]) );
  NAND2X0 U15 ( .IN1(n10), .IN2(n9), .QN(out1[2]) );
  NAND2X0 U16 ( .IN1(n58), .IN2(in2[18]), .QN(n59) );
  NAND2X0 U17 ( .IN1(n61), .IN2(in2[19]), .QN(n62) );
  NAND2X0 U18 ( .IN1(in1[1]), .IN2(in1[0]), .QN(out1[25]) );
  NOR2X0 U19 ( .IN1(in1[1]), .IN2(in1[0]), .QN(n71) );
  INVX0 U20 ( .INP(in2[0]), .ZN(n1) );
  INVX0 U21 ( .INP(in2[1]), .ZN(n2) );
  INVX0 U22 ( .INP(in2[3]), .ZN(n3) );
  INVX0 U23 ( .INP(in2[21]), .ZN(n4) );
  INVX0 U24 ( .INP(in2[22]), .ZN(n5) );
  INVX0 U25 ( .INP(in1[1]), .ZN(n6) );
  MUX21X1 U26 ( .IN1(in1[1]), .IN2(n6), .S(in1[0]), .Q(n74) );
  INVX0 U27 ( .INP(n74), .ZN(n76) );
  AO221X1 U28 ( .IN1(in2[0]), .IN2(in2[1]), .IN3(n1), .IN4(n2), .IN5(n76), .Q(
        n7) );
  MUX21X1 U29 ( .IN1(n2), .IN2(n8), .S(in2[2]), .Q(n12) );
  AO221X1 U30 ( .IN1(n12), .IN2(in2[2]), .IN3(n12), .IN4(n1), .IN5(n76), .Q(
        n10) );
  INVX0 U31 ( .INP(n71), .ZN(n13) );
  AO221X1 U32 ( .IN1(in2[0]), .IN2(in2[1]), .IN3(n1), .IN4(n2), .IN5(n13), .Q(
        n9) );
  NOR3X0 U33 ( .IN1(in2[0]), .IN2(in2[2]), .IN3(in2[1]), .QN(n11) );
  OR4X1 U34 ( .IN1(in2[3]), .IN2(in2[0]), .IN3(in2[2]), .IN4(in2[1]), .Q(n16)
         );
  OA21X1 U35 ( .IN1(n11), .IN2(n3), .IN3(n16), .Q(n18) );
  INVX0 U36 ( .INP(n18), .ZN(n14) );
  OAI222X1 U37 ( .IN1(n15), .IN2(in2[2]), .IN3(n14), .IN4(n76), .IN5(n13), 
        .IN6(n12), .QN(out1[3]) );
  OR2X1 U38 ( .IN1(in2[4]), .IN2(n16), .Q(n19) );
  NAND2X0 U39 ( .IN1(n16), .IN2(in2[4]), .QN(n17) );
  AND2X1 U40 ( .IN1(n19), .IN2(n17), .Q(n21) );
  AO22X1 U41 ( .IN1(n71), .IN2(n18), .IN3(n21), .IN4(n74), .Q(out1[4]) );
  OR2X1 U42 ( .IN1(in2[5]), .IN2(n19), .Q(n22) );
  AND2X1 U43 ( .IN1(n22), .IN2(n20), .Q(n24) );
  AO22X1 U44 ( .IN1(n71), .IN2(n21), .IN3(n24), .IN4(n74), .Q(out1[5]) );
  OR2X1 U45 ( .IN1(in2[6]), .IN2(n22), .Q(n25) );
  NAND2X0 U46 ( .IN1(n22), .IN2(in2[6]), .QN(n23) );
  AND2X1 U47 ( .IN1(n25), .IN2(n23), .Q(n27) );
  AO22X1 U48 ( .IN1(n71), .IN2(n24), .IN3(n27), .IN4(n74), .Q(out1[6]) );
  OR2X1 U49 ( .IN1(in2[7]), .IN2(n25), .Q(n28) );
  AND2X1 U50 ( .IN1(n28), .IN2(n26), .Q(n30) );
  AO22X1 U51 ( .IN1(n71), .IN2(n27), .IN3(n30), .IN4(n74), .Q(out1[7]) );
  OR2X1 U52 ( .IN1(in2[8]), .IN2(n28), .Q(n31) );
  NAND2X0 U53 ( .IN1(n28), .IN2(in2[8]), .QN(n29) );
  AND2X1 U54 ( .IN1(n31), .IN2(n29), .Q(n33) );
  AO22X1 U55 ( .IN1(n71), .IN2(n30), .IN3(n33), .IN4(n74), .Q(out1[8]) );
  OR2X1 U56 ( .IN1(in2[9]), .IN2(n31), .Q(n34) );
  AND2X1 U57 ( .IN1(n34), .IN2(n32), .Q(n36) );
  AO22X1 U58 ( .IN1(n71), .IN2(n33), .IN3(n36), .IN4(n74), .Q(out1[9]) );
  OR2X1 U59 ( .IN1(in2[10]), .IN2(n34), .Q(n37) );
  NAND2X0 U60 ( .IN1(n34), .IN2(in2[10]), .QN(n35) );
  AND2X1 U61 ( .IN1(n37), .IN2(n35), .Q(n39) );
  AO22X1 U62 ( .IN1(n71), .IN2(n36), .IN3(n39), .IN4(n74), .Q(out1[10]) );
  OR2X1 U63 ( .IN1(in2[11]), .IN2(n37), .Q(n40) );
  AND2X1 U64 ( .IN1(n40), .IN2(n38), .Q(n42) );
  AO22X1 U65 ( .IN1(n71), .IN2(n39), .IN3(n42), .IN4(n74), .Q(out1[11]) );
  OR2X1 U66 ( .IN1(in2[12]), .IN2(n40), .Q(n43) );
  NAND2X0 U67 ( .IN1(n40), .IN2(in2[12]), .QN(n41) );
  AND2X1 U68 ( .IN1(n43), .IN2(n41), .Q(n45) );
  AO22X1 U69 ( .IN1(n71), .IN2(n42), .IN3(n45), .IN4(n74), .Q(out1[12]) );
  OR2X1 U70 ( .IN1(in2[13]), .IN2(n43), .Q(n46) );
  AND2X1 U71 ( .IN1(n46), .IN2(n44), .Q(n48) );
  AO22X1 U72 ( .IN1(n71), .IN2(n45), .IN3(n48), .IN4(n74), .Q(out1[13]) );
  OR2X1 U73 ( .IN1(in2[14]), .IN2(n46), .Q(n49) );
  AND2X1 U74 ( .IN1(n49), .IN2(n47), .Q(n51) );
  AO22X1 U75 ( .IN1(n71), .IN2(n48), .IN3(n51), .IN4(n74), .Q(out1[14]) );
  OR2X1 U76 ( .IN1(in2[15]), .IN2(n49), .Q(n52) );
  AND2X1 U77 ( .IN1(n52), .IN2(n50), .Q(n54) );
  AO22X1 U78 ( .IN1(n71), .IN2(n51), .IN3(n54), .IN4(n74), .Q(out1[15]) );
  OR2X1 U79 ( .IN1(in2[16]), .IN2(n52), .Q(n55) );
  AND2X1 U80 ( .IN1(n55), .IN2(n53), .Q(n57) );
  AO22X1 U81 ( .IN1(n71), .IN2(n54), .IN3(n57), .IN4(n74), .Q(out1[16]) );
  OR2X1 U82 ( .IN1(in2[17]), .IN2(n55), .Q(n58) );
  AND2X1 U83 ( .IN1(n58), .IN2(n56), .Q(n60) );
  AO22X1 U84 ( .IN1(n71), .IN2(n57), .IN3(n60), .IN4(n74), .Q(out1[17]) );
  OR2X1 U85 ( .IN1(in2[18]), .IN2(n58), .Q(n61) );
  AND2X1 U86 ( .IN1(n61), .IN2(n59), .Q(n63) );
  AO22X1 U87 ( .IN1(n71), .IN2(n60), .IN3(n63), .IN4(n74), .Q(out1[18]) );
  OR2X1 U88 ( .IN1(in2[19]), .IN2(n61), .Q(n64) );
  AND2X1 U89 ( .IN1(n64), .IN2(n62), .Q(n65) );
  AO22X1 U90 ( .IN1(n71), .IN2(n63), .IN3(n65), .IN4(n74), .Q(out1[19]) );
  NOR2X0 U91 ( .IN1(in2[20]), .IN2(n64), .QN(n72) );
  AOI21X1 U92 ( .IN1(in2[20]), .IN2(n64), .IN3(n72), .QN(n66) );
  AO22X1 U93 ( .IN1(n71), .IN2(n65), .IN3(n66), .IN4(n74), .Q(out1[20]) );
  MUX21X1 U94 ( .IN1(n4), .IN2(in2[21]), .S(n72), .Q(n69) );
  AO22X1 U95 ( .IN1(n71), .IN2(n66), .IN3(n69), .IN4(n74), .Q(out1[21]) );
  INVX0 U96 ( .INP(n72), .ZN(n67) );
  NOR2X0 U97 ( .IN1(in2[21]), .IN2(n67), .QN(n70) );
  MUX21X1 U98 ( .IN1(n5), .IN2(in2[22]), .S(n70), .Q(n68) );
  AO22X1 U99 ( .IN1(n71), .IN2(n69), .IN3(n68), .IN4(n74), .Q(out1[22]) );
  MUX21X1 U100 ( .IN1(n71), .IN2(n74), .S(n70), .Q(n73) );
  AND3X1 U101 ( .IN1(n72), .IN2(n71), .IN3(n4), .Q(n75) );
  MUX21X1 U102 ( .IN1(n73), .IN2(n75), .S(in2[22]), .Q(out1[23]) );
  AO21X1 U103 ( .IN1(n75), .IN2(n5), .IN3(n74), .Q(out1[24]) );
  NOR2X0 U104 ( .IN1(n76), .IN2(n1), .QN(out1[0]) );
endmodule


module booth27_55 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n25), .IN2(n6), .QN(n30) );
  NAND2X0 U4 ( .IN1(n33), .IN2(n7), .QN(n37) );
  NAND2X0 U5 ( .IN1(n41), .IN2(n8), .QN(n45) );
  NAND2X0 U6 ( .IN1(n49), .IN2(n9), .QN(n53) );
  NAND2X0 U7 ( .IN1(n57), .IN2(n10), .QN(n61) );
  NAND2X0 U8 ( .IN1(n65), .IN2(n11), .QN(n77) );
  NAND2X0 U9 ( .IN1(n81), .IN2(n13), .QN(n89) );
  NAND2X0 U10 ( .IN1(n93), .IN2(n15), .QN(n101) );
  NAND2X0 U11 ( .IN1(n105), .IN2(n17), .QN(n114) );
  NAND2X0 U12 ( .IN1(n27), .IN2(n132), .QN(n4) );
  NAND2X0 U13 ( .IN1(in1[2]), .IN2(n77), .QN(n71) );
  NAND2X0 U14 ( .IN1(n70), .IN2(n132), .QN(n74) );
  NAND2X0 U15 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U16 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U17 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U18 ( .IN1(n118), .IN2(n19), .QN(n125) );
  NAND2X0 U19 ( .IN1(n141), .IN2(n130), .QN(n24) );
  NAND2X0 U20 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NAND2X0 U21 ( .IN1(n32), .IN2(n31), .QN(out1[3]) );
  NAND2X0 U22 ( .IN1(n36), .IN2(n35), .QN(out1[4]) );
  NAND2X0 U23 ( .IN1(n40), .IN2(n39), .QN(out1[5]) );
  NAND2X0 U24 ( .IN1(n44), .IN2(n43), .QN(out1[6]) );
  NAND2X0 U25 ( .IN1(n48), .IN2(n47), .QN(out1[7]) );
  NAND2X0 U26 ( .IN1(n52), .IN2(n51), .QN(out1[8]) );
  NAND2X0 U27 ( .IN1(n56), .IN2(n55), .QN(out1[9]) );
  NAND2X0 U28 ( .IN1(n60), .IN2(n59), .QN(out1[10]) );
  NAND2X0 U29 ( .IN1(n64), .IN2(n63), .QN(out1[11]) );
  NAND2X0 U30 ( .IN1(n69), .IN2(n68), .QN(out1[12]) );
  NAND2X0 U31 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U32 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U33 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U34 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U35 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U36 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U37 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U38 ( .IN1(n23), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U39 ( .IN1(in1[2]), .IN2(n22), .QN(n23) );
  NOR2X0 U40 ( .IN1(n28), .IN2(n26), .QN(n3) );
  NOR2X0 U41 ( .IN1(n142), .IN2(n21), .QN(n1) );
  NOR2X0 U42 ( .IN1(n142), .IN2(n111), .QN(n138) );
  INVX0 U43 ( .INP(n130), .ZN(n137) );
  INVX0 U44 ( .INP(n132), .ZN(n141) );
  NOR3X0 U45 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  NAND3X0 U46 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  MUX21X1 U47 ( .IN1(n22), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  INVX0 U48 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U49 ( .INP(in2[2]), .ZN(n6) );
  INVX0 U50 ( .INP(in2[4]), .ZN(n7) );
  INVX0 U51 ( .INP(in2[6]), .ZN(n8) );
  INVX0 U52 ( .INP(in2[8]), .ZN(n9) );
  INVX0 U53 ( .INP(in2[10]), .ZN(n10) );
  INVX0 U54 ( .INP(in2[12]), .ZN(n11) );
  INVX0 U55 ( .INP(in2[13]), .ZN(n12) );
  INVX0 U56 ( .INP(in2[14]), .ZN(n13) );
  INVX0 U57 ( .INP(in2[15]), .ZN(n14) );
  INVX0 U58 ( .INP(in2[16]), .ZN(n15) );
  INVX0 U59 ( .INP(in2[17]), .ZN(n16) );
  INVX0 U60 ( .INP(in2[18]), .ZN(n17) );
  INVX0 U61 ( .INP(in2[19]), .ZN(n18) );
  INVX0 U62 ( .INP(in2[20]), .ZN(n19) );
  INVX0 U63 ( .INP(in2[21]), .ZN(n20) );
  INVX0 U64 ( .INP(in2[22]), .ZN(n21) );
  INVX0 U65 ( .INP(in1[1]), .ZN(n22) );
  INVX0 U66 ( .INP(in1[2]), .ZN(n111) );
  INVX0 U67 ( .INP(n138), .ZN(n140) );
  NOR2X0 U68 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n25) );
  AOI21X1 U69 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n25), .QN(n27) );
  NOR2X0 U70 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U71 ( .IN1(n24), .IN2(in2[0]), .IN3(n138), .IN4(n27), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U72 ( .INP(n133), .ZN(n67) );
  NOR2X0 U73 ( .IN1(n67), .IN2(n6), .QN(n28) );
  OA21X1 U74 ( .IN1(n25), .IN2(n6), .IN3(n30), .Q(n29) );
  AO22X1 U75 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n29), .Q(n26) );
  AOI22X1 U76 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n29), .QN(n32) );
  NOR2X0 U77 ( .IN1(in2[3]), .IN2(n30), .QN(n33) );
  AO21X1 U78 ( .IN1(in2[3]), .IN2(n30), .IN3(n33), .Q(n34) );
  OA22X1 U79 ( .IN1(n6), .IN2(n130), .IN3(n140), .IN4(n34), .Q(n31) );
  OA21X1 U80 ( .IN1(n33), .IN2(n7), .IN3(n37), .Q(n38) );
  AOI22X1 U81 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n38), .QN(n36) );
  OA22X1 U82 ( .IN1(n67), .IN2(n7), .IN3(n141), .IN4(n34), .Q(n35) );
  NOR2X0 U83 ( .IN1(in2[5]), .IN2(n37), .QN(n41) );
  AO21X1 U84 ( .IN1(in2[5]), .IN2(n37), .IN3(n41), .Q(n42) );
  OA22X1 U85 ( .IN1(n7), .IN2(n130), .IN3(n140), .IN4(n42), .Q(n40) );
  AOI22X1 U86 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n38), .QN(n39) );
  OA21X1 U87 ( .IN1(n41), .IN2(n8), .IN3(n45), .Q(n46) );
  AOI22X1 U88 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n46), .QN(n44) );
  OA22X1 U89 ( .IN1(n67), .IN2(n8), .IN3(n141), .IN4(n42), .Q(n43) );
  NOR2X0 U90 ( .IN1(in2[7]), .IN2(n45), .QN(n49) );
  AO21X1 U91 ( .IN1(in2[7]), .IN2(n45), .IN3(n49), .Q(n50) );
  OA22X1 U92 ( .IN1(n8), .IN2(n130), .IN3(n140), .IN4(n50), .Q(n48) );
  AOI22X1 U93 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n46), .QN(n47) );
  OA21X1 U94 ( .IN1(n49), .IN2(n9), .IN3(n53), .Q(n54) );
  AOI22X1 U95 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n54), .QN(n52) );
  OA22X1 U96 ( .IN1(n67), .IN2(n9), .IN3(n141), .IN4(n50), .Q(n51) );
  NOR2X0 U97 ( .IN1(in2[9]), .IN2(n53), .QN(n57) );
  AO21X1 U98 ( .IN1(in2[9]), .IN2(n53), .IN3(n57), .Q(n58) );
  OA22X1 U99 ( .IN1(n9), .IN2(n130), .IN3(n140), .IN4(n58), .Q(n56) );
  AOI22X1 U100 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n54), .QN(n55) );
  OA21X1 U101 ( .IN1(n57), .IN2(n10), .IN3(n61), .Q(n62) );
  AOI22X1 U102 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n62), .QN(n60) );
  OA22X1 U103 ( .IN1(n67), .IN2(n10), .IN3(n141), .IN4(n58), .Q(n59) );
  NOR2X0 U104 ( .IN1(in2[11]), .IN2(n61), .QN(n65) );
  AO21X1 U105 ( .IN1(in2[11]), .IN2(n61), .IN3(n65), .Q(n66) );
  OA22X1 U106 ( .IN1(n10), .IN2(n130), .IN3(n140), .IN4(n66), .Q(n64) );
  AOI22X1 U107 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n62), .QN(n63) );
  OA21X1 U108 ( .IN1(n65), .IN2(n11), .IN3(n77), .Q(n70) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n70), .QN(n69) );
  OA22X1 U110 ( .IN1(n67), .IN2(n11), .IN3(n141), .IN4(n66), .Q(n68) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n12), .S(n71), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n11), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n13), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n12), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n12), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n14), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n13), .IN4(n85), .IN5(n84), 
        .Q(out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n15), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n14), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n14), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n16), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n15), .IN4(n97), .IN5(n96), 
        .Q(out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n17), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n16), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n16), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n18), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n17), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n19), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n18), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n18), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n20), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n19), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n21), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n20), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n20), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n21), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_56 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n33), .IN2(n7), .QN(n37) );
  NAND2X0 U4 ( .IN1(n41), .IN2(n8), .QN(n45) );
  NAND2X0 U5 ( .IN1(n49), .IN2(n9), .QN(n53) );
  NAND2X0 U6 ( .IN1(n57), .IN2(n10), .QN(n61) );
  NAND2X0 U7 ( .IN1(n25), .IN2(n6), .QN(n30) );
  NAND2X0 U8 ( .IN1(n65), .IN2(n11), .QN(n77) );
  NAND2X0 U9 ( .IN1(n81), .IN2(n13), .QN(n89) );
  NAND2X0 U10 ( .IN1(n93), .IN2(n15), .QN(n101) );
  NAND2X0 U11 ( .IN1(n105), .IN2(n17), .QN(n114) );
  NAND2X0 U12 ( .IN1(n118), .IN2(n19), .QN(n125) );
  NAND2X0 U13 ( .IN1(in1[2]), .IN2(n77), .QN(n71) );
  NAND2X0 U14 ( .IN1(n70), .IN2(n132), .QN(n74) );
  NAND2X0 U15 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U16 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U17 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U18 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U19 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U20 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U21 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U22 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NAND2X0 U23 ( .IN1(n27), .IN2(n132), .QN(n4) );
  NAND2X0 U24 ( .IN1(n32), .IN2(n31), .QN(out1[3]) );
  NAND2X0 U25 ( .IN1(n36), .IN2(n35), .QN(out1[4]) );
  NAND2X0 U26 ( .IN1(n40), .IN2(n39), .QN(out1[5]) );
  NAND2X0 U27 ( .IN1(n44), .IN2(n43), .QN(out1[6]) );
  NAND2X0 U28 ( .IN1(n48), .IN2(n47), .QN(out1[7]) );
  NAND2X0 U29 ( .IN1(n52), .IN2(n51), .QN(out1[8]) );
  NAND2X0 U30 ( .IN1(n56), .IN2(n55), .QN(out1[9]) );
  NAND2X0 U31 ( .IN1(n60), .IN2(n59), .QN(out1[10]) );
  NAND2X0 U32 ( .IN1(n64), .IN2(n63), .QN(out1[11]) );
  NAND2X0 U33 ( .IN1(n69), .IN2(n68), .QN(out1[12]) );
  NAND2X0 U34 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U35 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U36 ( .IN1(n141), .IN2(n130), .QN(n24) );
  NAND2X0 U37 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U38 ( .IN1(n23), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U39 ( .IN1(in1[2]), .IN2(n22), .QN(n23) );
  NOR2X0 U40 ( .IN1(n28), .IN2(n26), .QN(n3) );
  NOR2X0 U41 ( .IN1(n142), .IN2(n111), .QN(n138) );
  NOR2X0 U42 ( .IN1(n142), .IN2(n21), .QN(n1) );
  INVX0 U43 ( .INP(n130), .ZN(n137) );
  INVX0 U44 ( .INP(n132), .ZN(n141) );
  NOR3X0 U45 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  NAND3X0 U46 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  MUX21X1 U47 ( .IN1(n22), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  INVX0 U48 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U49 ( .INP(in2[2]), .ZN(n6) );
  INVX0 U50 ( .INP(in2[4]), .ZN(n7) );
  INVX0 U51 ( .INP(in2[6]), .ZN(n8) );
  INVX0 U52 ( .INP(in2[8]), .ZN(n9) );
  INVX0 U53 ( .INP(in2[10]), .ZN(n10) );
  INVX0 U54 ( .INP(in2[12]), .ZN(n11) );
  INVX0 U55 ( .INP(in2[13]), .ZN(n12) );
  INVX0 U56 ( .INP(in2[14]), .ZN(n13) );
  INVX0 U57 ( .INP(in2[15]), .ZN(n14) );
  INVX0 U58 ( .INP(in2[16]), .ZN(n15) );
  INVX0 U59 ( .INP(in2[17]), .ZN(n16) );
  INVX0 U60 ( .INP(in2[18]), .ZN(n17) );
  INVX0 U61 ( .INP(in2[19]), .ZN(n18) );
  INVX0 U62 ( .INP(in2[20]), .ZN(n19) );
  INVX0 U63 ( .INP(in2[21]), .ZN(n20) );
  INVX0 U64 ( .INP(in2[22]), .ZN(n21) );
  INVX0 U65 ( .INP(in1[1]), .ZN(n22) );
  INVX0 U66 ( .INP(in1[2]), .ZN(n111) );
  INVX0 U67 ( .INP(n138), .ZN(n140) );
  NOR2X0 U68 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n25) );
  AOI21X1 U69 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n25), .QN(n27) );
  NOR2X0 U70 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U71 ( .IN1(n24), .IN2(in2[0]), .IN3(n138), .IN4(n27), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U72 ( .INP(n133), .ZN(n67) );
  NOR2X0 U73 ( .IN1(n67), .IN2(n6), .QN(n28) );
  OA21X1 U74 ( .IN1(n25), .IN2(n6), .IN3(n30), .Q(n29) );
  AO22X1 U75 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n29), .Q(n26) );
  AOI22X1 U76 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n29), .QN(n32) );
  NOR2X0 U77 ( .IN1(in2[3]), .IN2(n30), .QN(n33) );
  AO21X1 U78 ( .IN1(in2[3]), .IN2(n30), .IN3(n33), .Q(n34) );
  OA22X1 U79 ( .IN1(n6), .IN2(n130), .IN3(n140), .IN4(n34), .Q(n31) );
  OA21X1 U80 ( .IN1(n33), .IN2(n7), .IN3(n37), .Q(n38) );
  AOI22X1 U81 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n38), .QN(n36) );
  OA22X1 U82 ( .IN1(n67), .IN2(n7), .IN3(n141), .IN4(n34), .Q(n35) );
  NOR2X0 U83 ( .IN1(in2[5]), .IN2(n37), .QN(n41) );
  AO21X1 U84 ( .IN1(in2[5]), .IN2(n37), .IN3(n41), .Q(n42) );
  OA22X1 U85 ( .IN1(n7), .IN2(n130), .IN3(n140), .IN4(n42), .Q(n40) );
  AOI22X1 U86 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n38), .QN(n39) );
  OA21X1 U87 ( .IN1(n41), .IN2(n8), .IN3(n45), .Q(n46) );
  AOI22X1 U88 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n46), .QN(n44) );
  OA22X1 U89 ( .IN1(n67), .IN2(n8), .IN3(n141), .IN4(n42), .Q(n43) );
  NOR2X0 U90 ( .IN1(in2[7]), .IN2(n45), .QN(n49) );
  AO21X1 U91 ( .IN1(in2[7]), .IN2(n45), .IN3(n49), .Q(n50) );
  OA22X1 U92 ( .IN1(n8), .IN2(n130), .IN3(n140), .IN4(n50), .Q(n48) );
  AOI22X1 U93 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n46), .QN(n47) );
  OA21X1 U94 ( .IN1(n49), .IN2(n9), .IN3(n53), .Q(n54) );
  AOI22X1 U95 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n54), .QN(n52) );
  OA22X1 U96 ( .IN1(n67), .IN2(n9), .IN3(n141), .IN4(n50), .Q(n51) );
  NOR2X0 U97 ( .IN1(in2[9]), .IN2(n53), .QN(n57) );
  AO21X1 U98 ( .IN1(in2[9]), .IN2(n53), .IN3(n57), .Q(n58) );
  OA22X1 U99 ( .IN1(n9), .IN2(n130), .IN3(n140), .IN4(n58), .Q(n56) );
  AOI22X1 U100 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n54), .QN(n55) );
  OA21X1 U101 ( .IN1(n57), .IN2(n10), .IN3(n61), .Q(n62) );
  AOI22X1 U102 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n62), .QN(n60) );
  OA22X1 U103 ( .IN1(n67), .IN2(n10), .IN3(n141), .IN4(n58), .Q(n59) );
  NOR2X0 U104 ( .IN1(in2[11]), .IN2(n61), .QN(n65) );
  AO21X1 U105 ( .IN1(in2[11]), .IN2(n61), .IN3(n65), .Q(n66) );
  OA22X1 U106 ( .IN1(n10), .IN2(n130), .IN3(n140), .IN4(n66), .Q(n64) );
  AOI22X1 U107 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n62), .QN(n63) );
  OA21X1 U108 ( .IN1(n65), .IN2(n11), .IN3(n77), .Q(n70) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n70), .QN(n69) );
  OA22X1 U110 ( .IN1(n67), .IN2(n11), .IN3(n141), .IN4(n66), .Q(n68) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n12), .S(n71), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n11), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n13), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n12), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n12), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n14), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n13), .IN4(n85), .IN5(n84), 
        .Q(out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n15), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n14), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n14), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n16), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n15), .IN4(n97), .IN5(n96), 
        .Q(out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n17), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n16), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n16), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n18), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n17), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n19), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n18), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n18), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n20), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n19), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n21), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n20), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n20), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n21), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_57 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n41), .IN2(n8), .QN(n45) );
  NAND2X0 U4 ( .IN1(n49), .IN2(n9), .QN(n53) );
  NAND2X0 U5 ( .IN1(n57), .IN2(n10), .QN(n61) );
  NAND2X0 U6 ( .IN1(n33), .IN2(n7), .QN(n37) );
  NAND2X0 U7 ( .IN1(n25), .IN2(n6), .QN(n30) );
  NAND2X0 U8 ( .IN1(n65), .IN2(n11), .QN(n77) );
  NAND2X0 U9 ( .IN1(n81), .IN2(n13), .QN(n89) );
  NAND2X0 U10 ( .IN1(n93), .IN2(n15), .QN(n101) );
  NAND2X0 U11 ( .IN1(in1[2]), .IN2(n77), .QN(n71) );
  NAND2X0 U12 ( .IN1(n70), .IN2(n132), .QN(n74) );
  NAND2X0 U13 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U14 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U15 ( .IN1(n105), .IN2(n17), .QN(n114) );
  NAND2X0 U16 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U17 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U18 ( .IN1(n27), .IN2(n132), .QN(n4) );
  NAND2X0 U19 ( .IN1(n141), .IN2(n130), .QN(n24) );
  NAND2X0 U20 ( .IN1(n40), .IN2(n39), .QN(out1[5]) );
  NAND2X0 U21 ( .IN1(n44), .IN2(n43), .QN(out1[6]) );
  NAND2X0 U22 ( .IN1(n48), .IN2(n47), .QN(out1[7]) );
  NAND2X0 U23 ( .IN1(n52), .IN2(n51), .QN(out1[8]) );
  NAND2X0 U24 ( .IN1(n56), .IN2(n55), .QN(out1[9]) );
  NAND2X0 U25 ( .IN1(n60), .IN2(n59), .QN(out1[10]) );
  NAND2X0 U26 ( .IN1(n64), .IN2(n63), .QN(out1[11]) );
  NAND2X0 U27 ( .IN1(n69), .IN2(n68), .QN(out1[12]) );
  NAND2X0 U28 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U29 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U30 ( .IN1(n118), .IN2(n19), .QN(n125) );
  NAND2X0 U31 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U32 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U33 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U34 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U35 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NAND2X0 U36 ( .IN1(n32), .IN2(n31), .QN(out1[3]) );
  NAND2X0 U37 ( .IN1(n36), .IN2(n35), .QN(out1[4]) );
  NAND2X0 U38 ( .IN1(n23), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U39 ( .IN1(in1[2]), .IN2(n22), .QN(n23) );
  INVX0 U40 ( .INP(in1[2]), .ZN(n111) );
  NOR2X0 U41 ( .IN1(n28), .IN2(n26), .QN(n3) );
  NOR2X0 U42 ( .IN1(n142), .IN2(n21), .QN(n1) );
  INVX0 U43 ( .INP(n132), .ZN(n141) );
  INVX0 U44 ( .INP(n130), .ZN(n137) );
  NOR2X0 U45 ( .IN1(n142), .IN2(n111), .QN(n138) );
  MUX21X1 U46 ( .IN1(n22), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  NAND3X0 U47 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  NOR3X0 U48 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  INVX0 U49 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U50 ( .INP(in2[2]), .ZN(n6) );
  INVX0 U51 ( .INP(in2[4]), .ZN(n7) );
  INVX0 U52 ( .INP(in2[6]), .ZN(n8) );
  INVX0 U53 ( .INP(in2[8]), .ZN(n9) );
  INVX0 U54 ( .INP(in2[10]), .ZN(n10) );
  INVX0 U55 ( .INP(in2[12]), .ZN(n11) );
  INVX0 U56 ( .INP(in2[13]), .ZN(n12) );
  INVX0 U57 ( .INP(in2[14]), .ZN(n13) );
  INVX0 U58 ( .INP(in2[15]), .ZN(n14) );
  INVX0 U59 ( .INP(in2[16]), .ZN(n15) );
  INVX0 U60 ( .INP(in2[17]), .ZN(n16) );
  INVX0 U61 ( .INP(in2[18]), .ZN(n17) );
  INVX0 U62 ( .INP(in2[19]), .ZN(n18) );
  INVX0 U63 ( .INP(in2[20]), .ZN(n19) );
  INVX0 U64 ( .INP(in2[21]), .ZN(n20) );
  INVX0 U65 ( .INP(in2[22]), .ZN(n21) );
  INVX0 U66 ( .INP(in1[1]), .ZN(n22) );
  INVX0 U67 ( .INP(n138), .ZN(n140) );
  NOR2X0 U68 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n25) );
  AOI21X1 U69 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n25), .QN(n27) );
  NOR2X0 U70 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U71 ( .IN1(n24), .IN2(in2[0]), .IN3(n138), .IN4(n27), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U72 ( .INP(n133), .ZN(n67) );
  NOR2X0 U73 ( .IN1(n67), .IN2(n6), .QN(n28) );
  OA21X1 U74 ( .IN1(n25), .IN2(n6), .IN3(n30), .Q(n29) );
  AO22X1 U75 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n29), .Q(n26) );
  AOI22X1 U76 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n29), .QN(n32) );
  NOR2X0 U77 ( .IN1(in2[3]), .IN2(n30), .QN(n33) );
  AO21X1 U78 ( .IN1(in2[3]), .IN2(n30), .IN3(n33), .Q(n34) );
  OA22X1 U79 ( .IN1(n6), .IN2(n130), .IN3(n140), .IN4(n34), .Q(n31) );
  OA21X1 U80 ( .IN1(n33), .IN2(n7), .IN3(n37), .Q(n38) );
  AOI22X1 U81 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n38), .QN(n36) );
  OA22X1 U82 ( .IN1(n67), .IN2(n7), .IN3(n141), .IN4(n34), .Q(n35) );
  NOR2X0 U83 ( .IN1(in2[5]), .IN2(n37), .QN(n41) );
  AO21X1 U84 ( .IN1(in2[5]), .IN2(n37), .IN3(n41), .Q(n42) );
  OA22X1 U85 ( .IN1(n7), .IN2(n130), .IN3(n140), .IN4(n42), .Q(n40) );
  AOI22X1 U86 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n38), .QN(n39) );
  OA21X1 U87 ( .IN1(n41), .IN2(n8), .IN3(n45), .Q(n46) );
  AOI22X1 U88 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n46), .QN(n44) );
  OA22X1 U89 ( .IN1(n67), .IN2(n8), .IN3(n141), .IN4(n42), .Q(n43) );
  NOR2X0 U90 ( .IN1(in2[7]), .IN2(n45), .QN(n49) );
  AO21X1 U91 ( .IN1(in2[7]), .IN2(n45), .IN3(n49), .Q(n50) );
  OA22X1 U92 ( .IN1(n8), .IN2(n130), .IN3(n140), .IN4(n50), .Q(n48) );
  AOI22X1 U93 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n46), .QN(n47) );
  OA21X1 U94 ( .IN1(n49), .IN2(n9), .IN3(n53), .Q(n54) );
  AOI22X1 U95 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n54), .QN(n52) );
  OA22X1 U96 ( .IN1(n67), .IN2(n9), .IN3(n141), .IN4(n50), .Q(n51) );
  NOR2X0 U97 ( .IN1(in2[9]), .IN2(n53), .QN(n57) );
  AO21X1 U98 ( .IN1(in2[9]), .IN2(n53), .IN3(n57), .Q(n58) );
  OA22X1 U99 ( .IN1(n9), .IN2(n130), .IN3(n140), .IN4(n58), .Q(n56) );
  AOI22X1 U100 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n54), .QN(n55) );
  OA21X1 U101 ( .IN1(n57), .IN2(n10), .IN3(n61), .Q(n62) );
  AOI22X1 U102 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n62), .QN(n60) );
  OA22X1 U103 ( .IN1(n67), .IN2(n10), .IN3(n141), .IN4(n58), .Q(n59) );
  NOR2X0 U104 ( .IN1(in2[11]), .IN2(n61), .QN(n65) );
  AO21X1 U105 ( .IN1(in2[11]), .IN2(n61), .IN3(n65), .Q(n66) );
  OA22X1 U106 ( .IN1(n10), .IN2(n130), .IN3(n140), .IN4(n66), .Q(n64) );
  AOI22X1 U107 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n62), .QN(n63) );
  OA21X1 U108 ( .IN1(n65), .IN2(n11), .IN3(n77), .Q(n70) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n70), .QN(n69) );
  OA22X1 U110 ( .IN1(n67), .IN2(n11), .IN3(n141), .IN4(n66), .Q(n68) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n12), .S(n71), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n11), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n13), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n12), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n12), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n14), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n13), .IN4(n85), .IN5(n84), 
        .Q(out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n15), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n14), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n14), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n16), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n15), .IN4(n97), .IN5(n96), 
        .Q(out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n17), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n16), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n16), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n18), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n17), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n19), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n18), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n18), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n20), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n19), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n21), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n20), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n20), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n21), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_58 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n49), .IN2(n9), .QN(n53) );
  NAND2X0 U4 ( .IN1(n57), .IN2(n10), .QN(n61) );
  NAND2X0 U5 ( .IN1(n25), .IN2(n6), .QN(n30) );
  NAND2X0 U6 ( .IN1(n41), .IN2(n8), .QN(n45) );
  NAND2X0 U7 ( .IN1(n33), .IN2(n7), .QN(n37) );
  NAND2X0 U8 ( .IN1(n65), .IN2(n11), .QN(n77) );
  NAND2X0 U9 ( .IN1(n81), .IN2(n13), .QN(n89) );
  NAND2X0 U10 ( .IN1(n93), .IN2(n15), .QN(n101) );
  NAND2X0 U11 ( .IN1(n105), .IN2(n17), .QN(n114) );
  NAND2X0 U12 ( .IN1(in1[2]), .IN2(n77), .QN(n71) );
  NAND2X0 U13 ( .IN1(n70), .IN2(n132), .QN(n74) );
  NAND2X0 U14 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U15 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U16 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U17 ( .IN1(n118), .IN2(n19), .QN(n125) );
  NAND2X0 U18 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U19 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U20 ( .IN1(n27), .IN2(n132), .QN(n4) );
  NAND2X0 U21 ( .IN1(n48), .IN2(n47), .QN(out1[7]) );
  NAND2X0 U22 ( .IN1(n52), .IN2(n51), .QN(out1[8]) );
  NAND2X0 U23 ( .IN1(n56), .IN2(n55), .QN(out1[9]) );
  NAND2X0 U24 ( .IN1(n60), .IN2(n59), .QN(out1[10]) );
  NAND2X0 U25 ( .IN1(n64), .IN2(n63), .QN(out1[11]) );
  NAND2X0 U26 ( .IN1(n69), .IN2(n68), .QN(out1[12]) );
  NAND2X0 U27 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U28 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U29 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U30 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U31 ( .IN1(n141), .IN2(n130), .QN(n24) );
  NAND2X0 U32 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NAND2X0 U33 ( .IN1(n36), .IN2(n35), .QN(out1[4]) );
  NAND2X0 U34 ( .IN1(n32), .IN2(n31), .QN(out1[3]) );
  NAND2X0 U35 ( .IN1(n40), .IN2(n39), .QN(out1[5]) );
  NAND2X0 U36 ( .IN1(n44), .IN2(n43), .QN(out1[6]) );
  NAND2X0 U37 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U38 ( .IN1(n23), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U39 ( .IN1(in1[2]), .IN2(n22), .QN(n23) );
  NOR2X0 U40 ( .IN1(n28), .IN2(n26), .QN(n3) );
  INVX0 U41 ( .INP(n130), .ZN(n137) );
  NAND3X0 U42 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  NOR2X0 U43 ( .IN1(n142), .IN2(n21), .QN(n1) );
  NOR2X0 U44 ( .IN1(n142), .IN2(n111), .QN(n138) );
  MUX21X1 U45 ( .IN1(n22), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  INVX0 U46 ( .INP(n132), .ZN(n141) );
  NOR3X0 U47 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  INVX0 U48 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U49 ( .INP(in2[2]), .ZN(n6) );
  INVX0 U50 ( .INP(in2[4]), .ZN(n7) );
  INVX0 U51 ( .INP(in2[6]), .ZN(n8) );
  INVX0 U52 ( .INP(in2[8]), .ZN(n9) );
  INVX0 U53 ( .INP(in2[10]), .ZN(n10) );
  INVX0 U54 ( .INP(in2[12]), .ZN(n11) );
  INVX0 U55 ( .INP(in2[13]), .ZN(n12) );
  INVX0 U56 ( .INP(in2[14]), .ZN(n13) );
  INVX0 U57 ( .INP(in2[15]), .ZN(n14) );
  INVX0 U58 ( .INP(in2[16]), .ZN(n15) );
  INVX0 U59 ( .INP(in2[17]), .ZN(n16) );
  INVX0 U60 ( .INP(in2[18]), .ZN(n17) );
  INVX0 U61 ( .INP(in2[19]), .ZN(n18) );
  INVX0 U62 ( .INP(in2[20]), .ZN(n19) );
  INVX0 U63 ( .INP(in2[21]), .ZN(n20) );
  INVX0 U64 ( .INP(in2[22]), .ZN(n21) );
  INVX0 U65 ( .INP(in1[1]), .ZN(n22) );
  INVX0 U66 ( .INP(in1[2]), .ZN(n111) );
  INVX0 U67 ( .INP(n138), .ZN(n140) );
  NOR2X0 U68 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n25) );
  AOI21X1 U69 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n25), .QN(n27) );
  NOR2X0 U70 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U71 ( .IN1(n24), .IN2(in2[0]), .IN3(n138), .IN4(n27), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U72 ( .INP(n133), .ZN(n67) );
  NOR2X0 U73 ( .IN1(n67), .IN2(n6), .QN(n28) );
  OA21X1 U74 ( .IN1(n25), .IN2(n6), .IN3(n30), .Q(n29) );
  AO22X1 U75 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n29), .Q(n26) );
  AOI22X1 U76 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n29), .QN(n32) );
  NOR2X0 U77 ( .IN1(in2[3]), .IN2(n30), .QN(n33) );
  AO21X1 U78 ( .IN1(in2[3]), .IN2(n30), .IN3(n33), .Q(n34) );
  OA22X1 U79 ( .IN1(n6), .IN2(n130), .IN3(n140), .IN4(n34), .Q(n31) );
  OA21X1 U80 ( .IN1(n33), .IN2(n7), .IN3(n37), .Q(n38) );
  AOI22X1 U81 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n38), .QN(n36) );
  OA22X1 U82 ( .IN1(n67), .IN2(n7), .IN3(n141), .IN4(n34), .Q(n35) );
  NOR2X0 U83 ( .IN1(in2[5]), .IN2(n37), .QN(n41) );
  AO21X1 U84 ( .IN1(in2[5]), .IN2(n37), .IN3(n41), .Q(n42) );
  OA22X1 U85 ( .IN1(n7), .IN2(n130), .IN3(n140), .IN4(n42), .Q(n40) );
  AOI22X1 U86 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n38), .QN(n39) );
  OA21X1 U87 ( .IN1(n41), .IN2(n8), .IN3(n45), .Q(n46) );
  AOI22X1 U88 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n46), .QN(n44) );
  OA22X1 U89 ( .IN1(n67), .IN2(n8), .IN3(n141), .IN4(n42), .Q(n43) );
  NOR2X0 U90 ( .IN1(in2[7]), .IN2(n45), .QN(n49) );
  AO21X1 U91 ( .IN1(in2[7]), .IN2(n45), .IN3(n49), .Q(n50) );
  OA22X1 U92 ( .IN1(n8), .IN2(n130), .IN3(n140), .IN4(n50), .Q(n48) );
  AOI22X1 U93 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n46), .QN(n47) );
  OA21X1 U94 ( .IN1(n49), .IN2(n9), .IN3(n53), .Q(n54) );
  AOI22X1 U95 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n54), .QN(n52) );
  OA22X1 U96 ( .IN1(n67), .IN2(n9), .IN3(n141), .IN4(n50), .Q(n51) );
  NOR2X0 U97 ( .IN1(in2[9]), .IN2(n53), .QN(n57) );
  AO21X1 U98 ( .IN1(in2[9]), .IN2(n53), .IN3(n57), .Q(n58) );
  OA22X1 U99 ( .IN1(n9), .IN2(n130), .IN3(n140), .IN4(n58), .Q(n56) );
  AOI22X1 U100 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n54), .QN(n55) );
  OA21X1 U101 ( .IN1(n57), .IN2(n10), .IN3(n61), .Q(n62) );
  AOI22X1 U102 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n62), .QN(n60) );
  OA22X1 U103 ( .IN1(n67), .IN2(n10), .IN3(n141), .IN4(n58), .Q(n59) );
  NOR2X0 U104 ( .IN1(in2[11]), .IN2(n61), .QN(n65) );
  AO21X1 U105 ( .IN1(in2[11]), .IN2(n61), .IN3(n65), .Q(n66) );
  OA22X1 U106 ( .IN1(n10), .IN2(n130), .IN3(n140), .IN4(n66), .Q(n64) );
  AOI22X1 U107 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n62), .QN(n63) );
  OA21X1 U108 ( .IN1(n65), .IN2(n11), .IN3(n77), .Q(n70) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n70), .QN(n69) );
  OA22X1 U110 ( .IN1(n67), .IN2(n11), .IN3(n141), .IN4(n66), .Q(n68) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n12), .S(n71), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n11), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n13), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n12), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n12), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n14), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n13), .IN4(n85), .IN5(n84), 
        .Q(out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n15), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n14), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n14), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n16), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n15), .IN4(n97), .IN5(n96), 
        .Q(out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n17), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n16), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n16), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n18), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n17), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n19), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n18), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n18), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n20), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n19), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n21), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n20), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n20), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n21), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_59 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n57), .IN2(n10), .QN(n61) );
  NAND2X0 U4 ( .IN1(n33), .IN2(n7), .QN(n37) );
  NAND2X0 U5 ( .IN1(n49), .IN2(n9), .QN(n53) );
  NAND2X0 U6 ( .IN1(n41), .IN2(n8), .QN(n45) );
  NAND2X0 U7 ( .IN1(n65), .IN2(n11), .QN(n77) );
  NAND2X0 U8 ( .IN1(n81), .IN2(n13), .QN(n89) );
  NAND2X0 U9 ( .IN1(n93), .IN2(n15), .QN(n101) );
  NAND2X0 U10 ( .IN1(n105), .IN2(n17), .QN(n114) );
  NAND2X0 U11 ( .IN1(n118), .IN2(n19), .QN(n125) );
  NAND2X0 U12 ( .IN1(n25), .IN2(n6), .QN(n30) );
  NAND2X0 U13 ( .IN1(in1[2]), .IN2(n77), .QN(n71) );
  NAND2X0 U14 ( .IN1(n70), .IN2(n132), .QN(n74) );
  NAND2X0 U15 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U16 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U17 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U18 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U19 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U20 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U21 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U22 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U23 ( .IN1(n56), .IN2(n55), .QN(out1[9]) );
  NAND2X0 U24 ( .IN1(n60), .IN2(n59), .QN(out1[10]) );
  NAND2X0 U25 ( .IN1(n64), .IN2(n63), .QN(out1[11]) );
  NAND2X0 U26 ( .IN1(n69), .IN2(n68), .QN(out1[12]) );
  NAND2X0 U27 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U28 ( .IN1(n23), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U29 ( .IN1(in1[2]), .IN2(n22), .QN(n23) );
  NAND2X0 U30 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NAND2X0 U31 ( .IN1(n27), .IN2(n132), .QN(n4) );
  NAND2X0 U32 ( .IN1(n32), .IN2(n31), .QN(out1[3]) );
  NAND2X0 U33 ( .IN1(n36), .IN2(n35), .QN(out1[4]) );
  NAND2X0 U34 ( .IN1(n44), .IN2(n43), .QN(out1[6]) );
  NAND2X0 U35 ( .IN1(n40), .IN2(n39), .QN(out1[5]) );
  NAND2X0 U36 ( .IN1(n48), .IN2(n47), .QN(out1[7]) );
  NAND2X0 U37 ( .IN1(n52), .IN2(n51), .QN(out1[8]) );
  NAND2X0 U38 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U39 ( .IN1(n141), .IN2(n130), .QN(n24) );
  NOR2X0 U40 ( .IN1(n28), .IN2(n26), .QN(n3) );
  NOR2X0 U41 ( .IN1(n142), .IN2(n21), .QN(n1) );
  INVX0 U42 ( .INP(n132), .ZN(n141) );
  INVX0 U43 ( .INP(n130), .ZN(n137) );
  NAND3X0 U44 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  NOR3X0 U45 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  NOR2X0 U46 ( .IN1(n142), .IN2(n111), .QN(n138) );
  MUX21X1 U47 ( .IN1(n22), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  INVX0 U48 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U49 ( .INP(in2[2]), .ZN(n6) );
  INVX0 U50 ( .INP(in2[4]), .ZN(n7) );
  INVX0 U51 ( .INP(in2[6]), .ZN(n8) );
  INVX0 U52 ( .INP(in2[8]), .ZN(n9) );
  INVX0 U53 ( .INP(in2[10]), .ZN(n10) );
  INVX0 U54 ( .INP(in2[12]), .ZN(n11) );
  INVX0 U55 ( .INP(in2[13]), .ZN(n12) );
  INVX0 U56 ( .INP(in2[14]), .ZN(n13) );
  INVX0 U57 ( .INP(in2[15]), .ZN(n14) );
  INVX0 U58 ( .INP(in2[16]), .ZN(n15) );
  INVX0 U59 ( .INP(in2[17]), .ZN(n16) );
  INVX0 U60 ( .INP(in2[18]), .ZN(n17) );
  INVX0 U61 ( .INP(in2[19]), .ZN(n18) );
  INVX0 U62 ( .INP(in2[20]), .ZN(n19) );
  INVX0 U63 ( .INP(in2[21]), .ZN(n20) );
  INVX0 U64 ( .INP(in2[22]), .ZN(n21) );
  INVX0 U65 ( .INP(in1[1]), .ZN(n22) );
  INVX0 U66 ( .INP(in1[2]), .ZN(n111) );
  INVX0 U67 ( .INP(n138), .ZN(n140) );
  NOR2X0 U68 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n25) );
  AOI21X1 U69 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n25), .QN(n27) );
  NOR2X0 U70 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U71 ( .IN1(n24), .IN2(in2[0]), .IN3(n138), .IN4(n27), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U72 ( .INP(n133), .ZN(n67) );
  NOR2X0 U73 ( .IN1(n67), .IN2(n6), .QN(n28) );
  OA21X1 U74 ( .IN1(n25), .IN2(n6), .IN3(n30), .Q(n29) );
  AO22X1 U75 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n29), .Q(n26) );
  AOI22X1 U76 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n29), .QN(n32) );
  NOR2X0 U77 ( .IN1(in2[3]), .IN2(n30), .QN(n33) );
  AO21X1 U78 ( .IN1(in2[3]), .IN2(n30), .IN3(n33), .Q(n34) );
  OA22X1 U79 ( .IN1(n6), .IN2(n130), .IN3(n140), .IN4(n34), .Q(n31) );
  OA21X1 U80 ( .IN1(n33), .IN2(n7), .IN3(n37), .Q(n38) );
  AOI22X1 U81 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n38), .QN(n36) );
  OA22X1 U82 ( .IN1(n67), .IN2(n7), .IN3(n141), .IN4(n34), .Q(n35) );
  NOR2X0 U83 ( .IN1(in2[5]), .IN2(n37), .QN(n41) );
  AO21X1 U84 ( .IN1(in2[5]), .IN2(n37), .IN3(n41), .Q(n42) );
  OA22X1 U85 ( .IN1(n7), .IN2(n130), .IN3(n140), .IN4(n42), .Q(n40) );
  AOI22X1 U86 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n38), .QN(n39) );
  OA21X1 U87 ( .IN1(n41), .IN2(n8), .IN3(n45), .Q(n46) );
  AOI22X1 U88 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n46), .QN(n44) );
  OA22X1 U89 ( .IN1(n67), .IN2(n8), .IN3(n141), .IN4(n42), .Q(n43) );
  NOR2X0 U90 ( .IN1(in2[7]), .IN2(n45), .QN(n49) );
  AO21X1 U91 ( .IN1(in2[7]), .IN2(n45), .IN3(n49), .Q(n50) );
  OA22X1 U92 ( .IN1(n8), .IN2(n130), .IN3(n140), .IN4(n50), .Q(n48) );
  AOI22X1 U93 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n46), .QN(n47) );
  OA21X1 U94 ( .IN1(n49), .IN2(n9), .IN3(n53), .Q(n54) );
  AOI22X1 U95 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n54), .QN(n52) );
  OA22X1 U96 ( .IN1(n67), .IN2(n9), .IN3(n141), .IN4(n50), .Q(n51) );
  NOR2X0 U97 ( .IN1(in2[9]), .IN2(n53), .QN(n57) );
  AO21X1 U98 ( .IN1(in2[9]), .IN2(n53), .IN3(n57), .Q(n58) );
  OA22X1 U99 ( .IN1(n9), .IN2(n130), .IN3(n140), .IN4(n58), .Q(n56) );
  AOI22X1 U100 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n54), .QN(n55) );
  OA21X1 U101 ( .IN1(n57), .IN2(n10), .IN3(n61), .Q(n62) );
  AOI22X1 U102 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n62), .QN(n60) );
  OA22X1 U103 ( .IN1(n67), .IN2(n10), .IN3(n141), .IN4(n58), .Q(n59) );
  NOR2X0 U104 ( .IN1(in2[11]), .IN2(n61), .QN(n65) );
  AO21X1 U105 ( .IN1(in2[11]), .IN2(n61), .IN3(n65), .Q(n66) );
  OA22X1 U106 ( .IN1(n10), .IN2(n130), .IN3(n140), .IN4(n66), .Q(n64) );
  AOI22X1 U107 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n62), .QN(n63) );
  OA21X1 U108 ( .IN1(n65), .IN2(n11), .IN3(n77), .Q(n70) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n70), .QN(n69) );
  OA22X1 U110 ( .IN1(n67), .IN2(n11), .IN3(n141), .IN4(n66), .Q(n68) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n12), .S(n71), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n11), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n13), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n12), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n12), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n14), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n13), .IN4(n85), .IN5(n84), 
        .Q(out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n15), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n14), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n14), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n16), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n15), .IN4(n97), .IN5(n96), 
        .Q(out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n17), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n16), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n16), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n18), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n17), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n19), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n18), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n18), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n20), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n19), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n21), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n20), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n20), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n21), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_60 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n57), .IN2(n10), .QN(n61) );
  NAND2X0 U4 ( .IN1(n25), .IN2(n6), .QN(n30) );
  NAND2X0 U5 ( .IN1(n33), .IN2(n7), .QN(n37) );
  NAND2X0 U6 ( .IN1(n49), .IN2(n9), .QN(n53) );
  NAND2X0 U7 ( .IN1(n41), .IN2(n8), .QN(n45) );
  NAND2X0 U8 ( .IN1(n65), .IN2(n11), .QN(n77) );
  NAND2X0 U9 ( .IN1(n81), .IN2(n13), .QN(n89) );
  NAND2X0 U10 ( .IN1(n93), .IN2(n15), .QN(n101) );
  NAND2X0 U11 ( .IN1(n105), .IN2(n17), .QN(n114) );
  NAND2X0 U12 ( .IN1(in1[2]), .IN2(n77), .QN(n71) );
  NAND2X0 U13 ( .IN1(n70), .IN2(n132), .QN(n74) );
  NAND2X0 U14 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U15 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U16 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U17 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U18 ( .IN1(n118), .IN2(n19), .QN(n125) );
  NAND2X0 U19 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U20 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U21 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U22 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U23 ( .IN1(n141), .IN2(n130), .QN(n24) );
  NAND2X0 U24 ( .IN1(n27), .IN2(n132), .QN(n4) );
  NAND2X0 U25 ( .IN1(n56), .IN2(n55), .QN(out1[9]) );
  NAND2X0 U26 ( .IN1(n60), .IN2(n59), .QN(out1[10]) );
  NAND2X0 U27 ( .IN1(n64), .IN2(n63), .QN(out1[11]) );
  NAND2X0 U28 ( .IN1(n69), .IN2(n68), .QN(out1[12]) );
  NAND2X0 U29 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U30 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U31 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NAND2X0 U32 ( .IN1(n32), .IN2(n31), .QN(out1[3]) );
  NAND2X0 U33 ( .IN1(n36), .IN2(n35), .QN(out1[4]) );
  NAND2X0 U34 ( .IN1(n40), .IN2(n39), .QN(out1[5]) );
  NAND2X0 U35 ( .IN1(n44), .IN2(n43), .QN(out1[6]) );
  NAND2X0 U36 ( .IN1(n48), .IN2(n47), .QN(out1[7]) );
  NAND2X0 U37 ( .IN1(n52), .IN2(n51), .QN(out1[8]) );
  NAND2X0 U38 ( .IN1(n23), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U39 ( .IN1(in1[2]), .IN2(n22), .QN(n23) );
  NOR2X0 U40 ( .IN1(n28), .IN2(n26), .QN(n3) );
  NOR2X0 U41 ( .IN1(n142), .IN2(n21), .QN(n1) );
  INVX0 U42 ( .INP(n132), .ZN(n141) );
  INVX0 U43 ( .INP(n130), .ZN(n137) );
  NAND3X0 U44 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  NOR3X0 U45 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  NOR2X0 U46 ( .IN1(n142), .IN2(n111), .QN(n138) );
  MUX21X1 U47 ( .IN1(n22), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  INVX0 U48 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U49 ( .INP(in2[2]), .ZN(n6) );
  INVX0 U50 ( .INP(in2[4]), .ZN(n7) );
  INVX0 U51 ( .INP(in2[6]), .ZN(n8) );
  INVX0 U52 ( .INP(in2[8]), .ZN(n9) );
  INVX0 U53 ( .INP(in2[10]), .ZN(n10) );
  INVX0 U54 ( .INP(in2[12]), .ZN(n11) );
  INVX0 U55 ( .INP(in2[13]), .ZN(n12) );
  INVX0 U56 ( .INP(in2[14]), .ZN(n13) );
  INVX0 U57 ( .INP(in2[15]), .ZN(n14) );
  INVX0 U58 ( .INP(in2[16]), .ZN(n15) );
  INVX0 U59 ( .INP(in2[17]), .ZN(n16) );
  INVX0 U60 ( .INP(in2[18]), .ZN(n17) );
  INVX0 U61 ( .INP(in2[19]), .ZN(n18) );
  INVX0 U62 ( .INP(in2[20]), .ZN(n19) );
  INVX0 U63 ( .INP(in2[21]), .ZN(n20) );
  INVX0 U64 ( .INP(in2[22]), .ZN(n21) );
  INVX0 U65 ( .INP(in1[1]), .ZN(n22) );
  INVX0 U66 ( .INP(in1[2]), .ZN(n111) );
  INVX0 U67 ( .INP(n138), .ZN(n140) );
  NOR2X0 U68 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n25) );
  AOI21X1 U69 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n25), .QN(n27) );
  NOR2X0 U70 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U71 ( .IN1(n24), .IN2(in2[0]), .IN3(n138), .IN4(n27), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U72 ( .INP(n133), .ZN(n67) );
  NOR2X0 U73 ( .IN1(n67), .IN2(n6), .QN(n28) );
  OA21X1 U74 ( .IN1(n25), .IN2(n6), .IN3(n30), .Q(n29) );
  AO22X1 U75 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n29), .Q(n26) );
  AOI22X1 U76 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n29), .QN(n32) );
  NOR2X0 U77 ( .IN1(in2[3]), .IN2(n30), .QN(n33) );
  AO21X1 U78 ( .IN1(in2[3]), .IN2(n30), .IN3(n33), .Q(n34) );
  OA22X1 U79 ( .IN1(n6), .IN2(n130), .IN3(n140), .IN4(n34), .Q(n31) );
  OA21X1 U80 ( .IN1(n33), .IN2(n7), .IN3(n37), .Q(n38) );
  AOI22X1 U81 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n38), .QN(n36) );
  OA22X1 U82 ( .IN1(n67), .IN2(n7), .IN3(n141), .IN4(n34), .Q(n35) );
  NOR2X0 U83 ( .IN1(in2[5]), .IN2(n37), .QN(n41) );
  AO21X1 U84 ( .IN1(in2[5]), .IN2(n37), .IN3(n41), .Q(n42) );
  OA22X1 U85 ( .IN1(n7), .IN2(n130), .IN3(n140), .IN4(n42), .Q(n40) );
  AOI22X1 U86 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n38), .QN(n39) );
  OA21X1 U87 ( .IN1(n41), .IN2(n8), .IN3(n45), .Q(n46) );
  AOI22X1 U88 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n46), .QN(n44) );
  OA22X1 U89 ( .IN1(n67), .IN2(n8), .IN3(n141), .IN4(n42), .Q(n43) );
  NOR2X0 U90 ( .IN1(in2[7]), .IN2(n45), .QN(n49) );
  AO21X1 U91 ( .IN1(in2[7]), .IN2(n45), .IN3(n49), .Q(n50) );
  OA22X1 U92 ( .IN1(n8), .IN2(n130), .IN3(n140), .IN4(n50), .Q(n48) );
  AOI22X1 U93 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n46), .QN(n47) );
  OA21X1 U94 ( .IN1(n49), .IN2(n9), .IN3(n53), .Q(n54) );
  AOI22X1 U95 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n54), .QN(n52) );
  OA22X1 U96 ( .IN1(n67), .IN2(n9), .IN3(n141), .IN4(n50), .Q(n51) );
  NOR2X0 U97 ( .IN1(in2[9]), .IN2(n53), .QN(n57) );
  AO21X1 U98 ( .IN1(in2[9]), .IN2(n53), .IN3(n57), .Q(n58) );
  OA22X1 U99 ( .IN1(n9), .IN2(n130), .IN3(n140), .IN4(n58), .Q(n56) );
  AOI22X1 U100 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n54), .QN(n55) );
  OA21X1 U101 ( .IN1(n57), .IN2(n10), .IN3(n61), .Q(n62) );
  AOI22X1 U102 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n62), .QN(n60) );
  OA22X1 U103 ( .IN1(n67), .IN2(n10), .IN3(n141), .IN4(n58), .Q(n59) );
  NOR2X0 U104 ( .IN1(in2[11]), .IN2(n61), .QN(n65) );
  AO21X1 U105 ( .IN1(in2[11]), .IN2(n61), .IN3(n65), .Q(n66) );
  OA22X1 U106 ( .IN1(n10), .IN2(n130), .IN3(n140), .IN4(n66), .Q(n64) );
  AOI22X1 U107 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n62), .QN(n63) );
  OA21X1 U108 ( .IN1(n65), .IN2(n11), .IN3(n77), .Q(n70) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n70), .QN(n69) );
  OA22X1 U110 ( .IN1(n67), .IN2(n11), .IN3(n141), .IN4(n66), .Q(n68) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n12), .S(n71), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n11), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n13), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n12), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n12), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n14), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n13), .IN4(n85), .IN5(n84), 
        .Q(out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n15), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n14), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n14), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n16), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n15), .IN4(n97), .IN5(n96), 
        .Q(out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n17), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n16), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n16), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n18), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n17), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n19), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n18), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n18), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n20), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n19), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n21), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n20), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n20), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n21), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_61 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n25), .IN2(n6), .QN(n30) );
  NAND2X0 U4 ( .IN1(n33), .IN2(n7), .QN(n37) );
  NAND2X0 U5 ( .IN1(n41), .IN2(n8), .QN(n45) );
  NAND2X0 U6 ( .IN1(n57), .IN2(n10), .QN(n61) );
  NAND2X0 U7 ( .IN1(n49), .IN2(n9), .QN(n53) );
  NAND2X0 U8 ( .IN1(n65), .IN2(n11), .QN(n77) );
  NAND2X0 U9 ( .IN1(n81), .IN2(n13), .QN(n89) );
  NAND2X0 U10 ( .IN1(n93), .IN2(n15), .QN(n101) );
  NAND2X0 U11 ( .IN1(n105), .IN2(n17), .QN(n114) );
  NAND2X0 U12 ( .IN1(n118), .IN2(n19), .QN(n125) );
  NAND2X0 U13 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U14 ( .IN1(in1[2]), .IN2(n77), .QN(n71) );
  NAND2X0 U15 ( .IN1(n70), .IN2(n132), .QN(n74) );
  NAND2X0 U16 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U17 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U18 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U19 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U20 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U21 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U22 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U23 ( .IN1(n141), .IN2(n130), .QN(n24) );
  NAND2X0 U24 ( .IN1(n27), .IN2(n132), .QN(n4) );
  NAND2X0 U25 ( .IN1(n64), .IN2(n63), .QN(out1[11]) );
  NAND2X0 U26 ( .IN1(n69), .IN2(n68), .QN(out1[12]) );
  NAND2X0 U27 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U28 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U29 ( .IN1(n23), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U30 ( .IN1(in1[2]), .IN2(n22), .QN(n23) );
  NAND2X0 U31 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NAND2X0 U32 ( .IN1(n32), .IN2(n31), .QN(out1[3]) );
  NAND2X0 U33 ( .IN1(n36), .IN2(n35), .QN(out1[4]) );
  NAND2X0 U34 ( .IN1(n40), .IN2(n39), .QN(out1[5]) );
  NAND2X0 U35 ( .IN1(n44), .IN2(n43), .QN(out1[6]) );
  NAND2X0 U36 ( .IN1(n48), .IN2(n47), .QN(out1[7]) );
  NAND2X0 U37 ( .IN1(n52), .IN2(n51), .QN(out1[8]) );
  NAND2X0 U38 ( .IN1(n56), .IN2(n55), .QN(out1[9]) );
  NAND2X0 U39 ( .IN1(n60), .IN2(n59), .QN(out1[10]) );
  NOR2X0 U40 ( .IN1(n28), .IN2(n26), .QN(n3) );
  NOR2X0 U41 ( .IN1(n142), .IN2(n21), .QN(n1) );
  INVX0 U42 ( .INP(n132), .ZN(n141) );
  INVX0 U43 ( .INP(n130), .ZN(n137) );
  NOR2X0 U44 ( .IN1(n142), .IN2(n111), .QN(n138) );
  MUX21X1 U45 ( .IN1(n22), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  NAND3X0 U46 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  NOR3X0 U47 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  INVX0 U48 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U49 ( .INP(in2[2]), .ZN(n6) );
  INVX0 U50 ( .INP(in2[4]), .ZN(n7) );
  INVX0 U51 ( .INP(in2[6]), .ZN(n8) );
  INVX0 U52 ( .INP(in2[8]), .ZN(n9) );
  INVX0 U53 ( .INP(in2[10]), .ZN(n10) );
  INVX0 U54 ( .INP(in2[12]), .ZN(n11) );
  INVX0 U55 ( .INP(in2[13]), .ZN(n12) );
  INVX0 U56 ( .INP(in2[14]), .ZN(n13) );
  INVX0 U57 ( .INP(in2[15]), .ZN(n14) );
  INVX0 U58 ( .INP(in2[16]), .ZN(n15) );
  INVX0 U59 ( .INP(in2[17]), .ZN(n16) );
  INVX0 U60 ( .INP(in2[18]), .ZN(n17) );
  INVX0 U61 ( .INP(in2[19]), .ZN(n18) );
  INVX0 U62 ( .INP(in2[20]), .ZN(n19) );
  INVX0 U63 ( .INP(in2[21]), .ZN(n20) );
  INVX0 U64 ( .INP(in2[22]), .ZN(n21) );
  INVX0 U65 ( .INP(in1[1]), .ZN(n22) );
  INVX0 U66 ( .INP(in1[2]), .ZN(n111) );
  INVX0 U67 ( .INP(n138), .ZN(n140) );
  NOR2X0 U68 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n25) );
  AOI21X1 U69 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n25), .QN(n27) );
  NOR2X0 U70 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U71 ( .IN1(n24), .IN2(in2[0]), .IN3(n138), .IN4(n27), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U72 ( .INP(n133), .ZN(n67) );
  NOR2X0 U73 ( .IN1(n67), .IN2(n6), .QN(n28) );
  OA21X1 U74 ( .IN1(n25), .IN2(n6), .IN3(n30), .Q(n29) );
  AO22X1 U75 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n29), .Q(n26) );
  AOI22X1 U76 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n29), .QN(n32) );
  NOR2X0 U77 ( .IN1(in2[3]), .IN2(n30), .QN(n33) );
  AO21X1 U78 ( .IN1(in2[3]), .IN2(n30), .IN3(n33), .Q(n34) );
  OA22X1 U79 ( .IN1(n6), .IN2(n130), .IN3(n140), .IN4(n34), .Q(n31) );
  OA21X1 U80 ( .IN1(n33), .IN2(n7), .IN3(n37), .Q(n38) );
  AOI22X1 U81 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n38), .QN(n36) );
  OA22X1 U82 ( .IN1(n67), .IN2(n7), .IN3(n141), .IN4(n34), .Q(n35) );
  NOR2X0 U83 ( .IN1(in2[5]), .IN2(n37), .QN(n41) );
  AO21X1 U84 ( .IN1(in2[5]), .IN2(n37), .IN3(n41), .Q(n42) );
  OA22X1 U85 ( .IN1(n7), .IN2(n130), .IN3(n140), .IN4(n42), .Q(n40) );
  AOI22X1 U86 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n38), .QN(n39) );
  OA21X1 U87 ( .IN1(n41), .IN2(n8), .IN3(n45), .Q(n46) );
  AOI22X1 U88 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n46), .QN(n44) );
  OA22X1 U89 ( .IN1(n67), .IN2(n8), .IN3(n141), .IN4(n42), .Q(n43) );
  NOR2X0 U90 ( .IN1(in2[7]), .IN2(n45), .QN(n49) );
  AO21X1 U91 ( .IN1(in2[7]), .IN2(n45), .IN3(n49), .Q(n50) );
  OA22X1 U92 ( .IN1(n8), .IN2(n130), .IN3(n140), .IN4(n50), .Q(n48) );
  AOI22X1 U93 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n46), .QN(n47) );
  OA21X1 U94 ( .IN1(n49), .IN2(n9), .IN3(n53), .Q(n54) );
  AOI22X1 U95 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n54), .QN(n52) );
  OA22X1 U96 ( .IN1(n67), .IN2(n9), .IN3(n141), .IN4(n50), .Q(n51) );
  NOR2X0 U97 ( .IN1(in2[9]), .IN2(n53), .QN(n57) );
  AO21X1 U98 ( .IN1(in2[9]), .IN2(n53), .IN3(n57), .Q(n58) );
  OA22X1 U99 ( .IN1(n9), .IN2(n130), .IN3(n140), .IN4(n58), .Q(n56) );
  AOI22X1 U100 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n54), .QN(n55) );
  OA21X1 U101 ( .IN1(n57), .IN2(n10), .IN3(n61), .Q(n62) );
  AOI22X1 U102 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n62), .QN(n60) );
  OA22X1 U103 ( .IN1(n67), .IN2(n10), .IN3(n141), .IN4(n58), .Q(n59) );
  NOR2X0 U104 ( .IN1(in2[11]), .IN2(n61), .QN(n65) );
  AO21X1 U105 ( .IN1(in2[11]), .IN2(n61), .IN3(n65), .Q(n66) );
  OA22X1 U106 ( .IN1(n10), .IN2(n130), .IN3(n140), .IN4(n66), .Q(n64) );
  AOI22X1 U107 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n62), .QN(n63) );
  OA21X1 U108 ( .IN1(n65), .IN2(n11), .IN3(n77), .Q(n70) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n70), .QN(n69) );
  OA22X1 U110 ( .IN1(n67), .IN2(n11), .IN3(n141), .IN4(n66), .Q(n68) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n12), .S(n71), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n11), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n13), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n12), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n12), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n14), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n13), .IN4(n85), .IN5(n84), 
        .Q(out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n15), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n14), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n14), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n16), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n15), .IN4(n97), .IN5(n96), 
        .Q(out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n17), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n16), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n16), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n18), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n17), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n19), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n18), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n18), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n20), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n19), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n21), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n20), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n20), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n21), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_62 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n25), .IN2(n6), .QN(n30) );
  NAND2X0 U4 ( .IN1(n33), .IN2(n7), .QN(n37) );
  NAND2X0 U5 ( .IN1(n41), .IN2(n8), .QN(n45) );
  NAND2X0 U6 ( .IN1(n49), .IN2(n9), .QN(n53) );
  NAND2X0 U7 ( .IN1(n57), .IN2(n10), .QN(n61) );
  NAND2X0 U8 ( .IN1(n65), .IN2(n11), .QN(n77) );
  NAND2X0 U9 ( .IN1(n81), .IN2(n13), .QN(n89) );
  NAND2X0 U10 ( .IN1(n93), .IN2(n15), .QN(n101) );
  NAND2X0 U11 ( .IN1(n105), .IN2(n17), .QN(n114) );
  NAND2X0 U12 ( .IN1(n118), .IN2(n19), .QN(n125) );
  NAND2X0 U13 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U14 ( .IN1(in1[2]), .IN2(n77), .QN(n71) );
  NAND2X0 U15 ( .IN1(n70), .IN2(n132), .QN(n74) );
  NAND2X0 U16 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U17 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U18 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U19 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U20 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U21 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U22 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U23 ( .IN1(n23), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U24 ( .IN1(in1[2]), .IN2(n22), .QN(n23) );
  NAND2X0 U25 ( .IN1(n32), .IN2(n31), .QN(out1[3]) );
  NAND2X0 U26 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U27 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U28 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NAND2X0 U29 ( .IN1(n27), .IN2(n132), .QN(n4) );
  NAND2X0 U30 ( .IN1(n36), .IN2(n35), .QN(out1[4]) );
  NAND2X0 U31 ( .IN1(n40), .IN2(n39), .QN(out1[5]) );
  NAND2X0 U32 ( .IN1(n44), .IN2(n43), .QN(out1[6]) );
  NAND2X0 U33 ( .IN1(n48), .IN2(n47), .QN(out1[7]) );
  NAND2X0 U34 ( .IN1(n52), .IN2(n51), .QN(out1[8]) );
  NAND2X0 U35 ( .IN1(n56), .IN2(n55), .QN(out1[9]) );
  NAND2X0 U36 ( .IN1(n60), .IN2(n59), .QN(out1[10]) );
  NAND2X0 U37 ( .IN1(n64), .IN2(n63), .QN(out1[11]) );
  NAND2X0 U38 ( .IN1(n69), .IN2(n68), .QN(out1[12]) );
  NAND2X0 U39 ( .IN1(n141), .IN2(n130), .QN(n24) );
  NOR2X0 U40 ( .IN1(n28), .IN2(n26), .QN(n3) );
  INVX0 U41 ( .INP(n130), .ZN(n137) );
  NAND3X0 U42 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  NOR2X0 U43 ( .IN1(n142), .IN2(n21), .QN(n1) );
  NOR2X0 U44 ( .IN1(n142), .IN2(n111), .QN(n138) );
  MUX21X1 U45 ( .IN1(n22), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  INVX0 U46 ( .INP(n132), .ZN(n141) );
  NOR3X0 U47 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  INVX0 U48 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U49 ( .INP(in2[2]), .ZN(n6) );
  INVX0 U50 ( .INP(in2[4]), .ZN(n7) );
  INVX0 U51 ( .INP(in2[6]), .ZN(n8) );
  INVX0 U52 ( .INP(in2[8]), .ZN(n9) );
  INVX0 U53 ( .INP(in2[10]), .ZN(n10) );
  INVX0 U54 ( .INP(in2[12]), .ZN(n11) );
  INVX0 U55 ( .INP(in2[13]), .ZN(n12) );
  INVX0 U56 ( .INP(in2[14]), .ZN(n13) );
  INVX0 U57 ( .INP(in2[15]), .ZN(n14) );
  INVX0 U58 ( .INP(in2[16]), .ZN(n15) );
  INVX0 U59 ( .INP(in2[17]), .ZN(n16) );
  INVX0 U60 ( .INP(in2[18]), .ZN(n17) );
  INVX0 U61 ( .INP(in2[19]), .ZN(n18) );
  INVX0 U62 ( .INP(in2[20]), .ZN(n19) );
  INVX0 U63 ( .INP(in2[21]), .ZN(n20) );
  INVX0 U64 ( .INP(in2[22]), .ZN(n21) );
  INVX0 U65 ( .INP(in1[1]), .ZN(n22) );
  INVX0 U66 ( .INP(in1[2]), .ZN(n111) );
  INVX0 U67 ( .INP(n138), .ZN(n140) );
  NOR2X0 U68 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n25) );
  AOI21X1 U69 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n25), .QN(n27) );
  NOR2X0 U70 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U71 ( .IN1(n24), .IN2(in2[0]), .IN3(n138), .IN4(n27), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U72 ( .INP(n133), .ZN(n67) );
  NOR2X0 U73 ( .IN1(n67), .IN2(n6), .QN(n28) );
  OA21X1 U74 ( .IN1(n25), .IN2(n6), .IN3(n30), .Q(n29) );
  AO22X1 U75 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n29), .Q(n26) );
  AOI22X1 U76 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n29), .QN(n32) );
  NOR2X0 U77 ( .IN1(in2[3]), .IN2(n30), .QN(n33) );
  AO21X1 U78 ( .IN1(in2[3]), .IN2(n30), .IN3(n33), .Q(n34) );
  OA22X1 U79 ( .IN1(n6), .IN2(n130), .IN3(n140), .IN4(n34), .Q(n31) );
  OA21X1 U80 ( .IN1(n33), .IN2(n7), .IN3(n37), .Q(n38) );
  AOI22X1 U81 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n38), .QN(n36) );
  OA22X1 U82 ( .IN1(n67), .IN2(n7), .IN3(n141), .IN4(n34), .Q(n35) );
  NOR2X0 U83 ( .IN1(in2[5]), .IN2(n37), .QN(n41) );
  AO21X1 U84 ( .IN1(in2[5]), .IN2(n37), .IN3(n41), .Q(n42) );
  OA22X1 U85 ( .IN1(n7), .IN2(n130), .IN3(n140), .IN4(n42), .Q(n40) );
  AOI22X1 U86 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n38), .QN(n39) );
  OA21X1 U87 ( .IN1(n41), .IN2(n8), .IN3(n45), .Q(n46) );
  AOI22X1 U88 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n46), .QN(n44) );
  OA22X1 U89 ( .IN1(n67), .IN2(n8), .IN3(n141), .IN4(n42), .Q(n43) );
  NOR2X0 U90 ( .IN1(in2[7]), .IN2(n45), .QN(n49) );
  AO21X1 U91 ( .IN1(in2[7]), .IN2(n45), .IN3(n49), .Q(n50) );
  OA22X1 U92 ( .IN1(n8), .IN2(n130), .IN3(n140), .IN4(n50), .Q(n48) );
  AOI22X1 U93 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n46), .QN(n47) );
  OA21X1 U94 ( .IN1(n49), .IN2(n9), .IN3(n53), .Q(n54) );
  AOI22X1 U95 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n54), .QN(n52) );
  OA22X1 U96 ( .IN1(n67), .IN2(n9), .IN3(n141), .IN4(n50), .Q(n51) );
  NOR2X0 U97 ( .IN1(in2[9]), .IN2(n53), .QN(n57) );
  AO21X1 U98 ( .IN1(in2[9]), .IN2(n53), .IN3(n57), .Q(n58) );
  OA22X1 U99 ( .IN1(n9), .IN2(n130), .IN3(n140), .IN4(n58), .Q(n56) );
  AOI22X1 U100 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n54), .QN(n55) );
  OA21X1 U101 ( .IN1(n57), .IN2(n10), .IN3(n61), .Q(n62) );
  AOI22X1 U102 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n62), .QN(n60) );
  OA22X1 U103 ( .IN1(n67), .IN2(n10), .IN3(n141), .IN4(n58), .Q(n59) );
  NOR2X0 U104 ( .IN1(in2[11]), .IN2(n61), .QN(n65) );
  AO21X1 U105 ( .IN1(in2[11]), .IN2(n61), .IN3(n65), .Q(n66) );
  OA22X1 U106 ( .IN1(n10), .IN2(n130), .IN3(n140), .IN4(n66), .Q(n64) );
  AOI22X1 U107 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n62), .QN(n63) );
  OA21X1 U108 ( .IN1(n65), .IN2(n11), .IN3(n77), .Q(n70) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n70), .QN(n69) );
  OA22X1 U110 ( .IN1(n67), .IN2(n11), .IN3(n141), .IN4(n66), .Q(n68) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n12), .S(n71), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n11), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n13), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n12), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n12), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n14), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n13), .IN4(n85), .IN5(n84), 
        .Q(out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n15), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n14), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n14), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n16), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n15), .IN4(n97), .IN5(n96), 
        .Q(out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n17), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n16), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n16), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n18), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n17), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n19), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n18), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n18), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n20), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n19), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n21), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n20), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n20), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n21), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_63 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n25), .IN2(n6), .QN(n30) );
  NAND2X0 U4 ( .IN1(n33), .IN2(n7), .QN(n37) );
  NAND2X0 U5 ( .IN1(n41), .IN2(n8), .QN(n45) );
  NAND2X0 U6 ( .IN1(n49), .IN2(n9), .QN(n53) );
  NAND2X0 U7 ( .IN1(n57), .IN2(n10), .QN(n61) );
  NAND2X0 U8 ( .IN1(n65), .IN2(n11), .QN(n77) );
  NAND2X0 U9 ( .IN1(n81), .IN2(n13), .QN(n89) );
  NAND2X0 U10 ( .IN1(n105), .IN2(n17), .QN(n114) );
  NAND2X0 U11 ( .IN1(n93), .IN2(n15), .QN(n101) );
  NAND2X0 U12 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U13 ( .IN1(n118), .IN2(n19), .QN(n125) );
  NAND2X0 U14 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U15 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U16 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U17 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U18 ( .IN1(n27), .IN2(n132), .QN(n4) );
  NAND2X0 U19 ( .IN1(n141), .IN2(n130), .QN(n24) );
  NAND2X0 U20 ( .IN1(n32), .IN2(n31), .QN(out1[3]) );
  NAND2X0 U21 ( .IN1(n36), .IN2(n35), .QN(out1[4]) );
  NAND2X0 U22 ( .IN1(in1[2]), .IN2(n77), .QN(n71) );
  NAND2X0 U23 ( .IN1(n70), .IN2(n132), .QN(n74) );
  NAND2X0 U24 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U25 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U26 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U27 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U28 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NAND2X0 U29 ( .IN1(n40), .IN2(n39), .QN(out1[5]) );
  NAND2X0 U30 ( .IN1(n44), .IN2(n43), .QN(out1[6]) );
  NAND2X0 U31 ( .IN1(n48), .IN2(n47), .QN(out1[7]) );
  NAND2X0 U32 ( .IN1(n52), .IN2(n51), .QN(out1[8]) );
  NAND2X0 U33 ( .IN1(n56), .IN2(n55), .QN(out1[9]) );
  NAND2X0 U34 ( .IN1(n60), .IN2(n59), .QN(out1[10]) );
  NAND2X0 U35 ( .IN1(n64), .IN2(n63), .QN(out1[11]) );
  NAND2X0 U36 ( .IN1(n69), .IN2(n68), .QN(out1[12]) );
  NAND2X0 U37 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U38 ( .IN1(n23), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U39 ( .IN1(in1[2]), .IN2(n22), .QN(n23) );
  INVX0 U40 ( .INP(in1[2]), .ZN(n111) );
  NOR2X0 U41 ( .IN1(n28), .IN2(n26), .QN(n3) );
  NOR2X0 U42 ( .IN1(n142), .IN2(n21), .QN(n1) );
  INVX0 U43 ( .INP(n132), .ZN(n141) );
  INVX0 U44 ( .INP(n130), .ZN(n137) );
  NAND3X0 U45 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  NOR2X0 U46 ( .IN1(n142), .IN2(n111), .QN(n138) );
  MUX21X1 U47 ( .IN1(n22), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  NOR3X0 U48 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  INVX0 U49 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U50 ( .INP(in2[2]), .ZN(n6) );
  INVX0 U51 ( .INP(in2[4]), .ZN(n7) );
  INVX0 U52 ( .INP(in2[6]), .ZN(n8) );
  INVX0 U53 ( .INP(in2[8]), .ZN(n9) );
  INVX0 U54 ( .INP(in2[10]), .ZN(n10) );
  INVX0 U55 ( .INP(in2[12]), .ZN(n11) );
  INVX0 U56 ( .INP(in2[13]), .ZN(n12) );
  INVX0 U57 ( .INP(in2[14]), .ZN(n13) );
  INVX0 U58 ( .INP(in2[15]), .ZN(n14) );
  INVX0 U59 ( .INP(in2[16]), .ZN(n15) );
  INVX0 U60 ( .INP(in2[17]), .ZN(n16) );
  INVX0 U61 ( .INP(in2[18]), .ZN(n17) );
  INVX0 U62 ( .INP(in2[19]), .ZN(n18) );
  INVX0 U63 ( .INP(in2[20]), .ZN(n19) );
  INVX0 U64 ( .INP(in2[21]), .ZN(n20) );
  INVX0 U65 ( .INP(in2[22]), .ZN(n21) );
  INVX0 U66 ( .INP(in1[1]), .ZN(n22) );
  INVX0 U67 ( .INP(n138), .ZN(n140) );
  NOR2X0 U68 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n25) );
  AOI21X1 U69 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n25), .QN(n27) );
  NOR2X0 U70 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U71 ( .IN1(n24), .IN2(in2[0]), .IN3(n138), .IN4(n27), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U72 ( .INP(n133), .ZN(n67) );
  NOR2X0 U73 ( .IN1(n67), .IN2(n6), .QN(n28) );
  OA21X1 U74 ( .IN1(n25), .IN2(n6), .IN3(n30), .Q(n29) );
  AO22X1 U75 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n29), .Q(n26) );
  AOI22X1 U76 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n29), .QN(n32) );
  NOR2X0 U77 ( .IN1(in2[3]), .IN2(n30), .QN(n33) );
  AO21X1 U78 ( .IN1(in2[3]), .IN2(n30), .IN3(n33), .Q(n34) );
  OA22X1 U79 ( .IN1(n6), .IN2(n130), .IN3(n140), .IN4(n34), .Q(n31) );
  OA21X1 U80 ( .IN1(n33), .IN2(n7), .IN3(n37), .Q(n38) );
  AOI22X1 U81 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n38), .QN(n36) );
  OA22X1 U82 ( .IN1(n67), .IN2(n7), .IN3(n141), .IN4(n34), .Q(n35) );
  NOR2X0 U83 ( .IN1(in2[5]), .IN2(n37), .QN(n41) );
  AO21X1 U84 ( .IN1(in2[5]), .IN2(n37), .IN3(n41), .Q(n42) );
  OA22X1 U85 ( .IN1(n7), .IN2(n130), .IN3(n140), .IN4(n42), .Q(n40) );
  AOI22X1 U86 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n38), .QN(n39) );
  OA21X1 U87 ( .IN1(n41), .IN2(n8), .IN3(n45), .Q(n46) );
  AOI22X1 U88 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n46), .QN(n44) );
  OA22X1 U89 ( .IN1(n67), .IN2(n8), .IN3(n141), .IN4(n42), .Q(n43) );
  NOR2X0 U90 ( .IN1(in2[7]), .IN2(n45), .QN(n49) );
  AO21X1 U91 ( .IN1(in2[7]), .IN2(n45), .IN3(n49), .Q(n50) );
  OA22X1 U92 ( .IN1(n8), .IN2(n130), .IN3(n140), .IN4(n50), .Q(n48) );
  AOI22X1 U93 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n46), .QN(n47) );
  OA21X1 U94 ( .IN1(n49), .IN2(n9), .IN3(n53), .Q(n54) );
  AOI22X1 U95 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n54), .QN(n52) );
  OA22X1 U96 ( .IN1(n67), .IN2(n9), .IN3(n141), .IN4(n50), .Q(n51) );
  NOR2X0 U97 ( .IN1(in2[9]), .IN2(n53), .QN(n57) );
  AO21X1 U98 ( .IN1(in2[9]), .IN2(n53), .IN3(n57), .Q(n58) );
  OA22X1 U99 ( .IN1(n9), .IN2(n130), .IN3(n140), .IN4(n58), .Q(n56) );
  AOI22X1 U100 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n54), .QN(n55) );
  OA21X1 U101 ( .IN1(n57), .IN2(n10), .IN3(n61), .Q(n62) );
  AOI22X1 U102 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n62), .QN(n60) );
  OA22X1 U103 ( .IN1(n67), .IN2(n10), .IN3(n141), .IN4(n58), .Q(n59) );
  NOR2X0 U104 ( .IN1(in2[11]), .IN2(n61), .QN(n65) );
  AO21X1 U105 ( .IN1(in2[11]), .IN2(n61), .IN3(n65), .Q(n66) );
  OA22X1 U106 ( .IN1(n10), .IN2(n130), .IN3(n140), .IN4(n66), .Q(n64) );
  AOI22X1 U107 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n62), .QN(n63) );
  OA21X1 U108 ( .IN1(n65), .IN2(n11), .IN3(n77), .Q(n70) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n70), .QN(n69) );
  OA22X1 U110 ( .IN1(n67), .IN2(n11), .IN3(n141), .IN4(n66), .Q(n68) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n12), .S(n71), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n11), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n13), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n12), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n12), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n14), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n13), .IN4(n85), .IN5(n84), 
        .Q(out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n15), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n14), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n14), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n16), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n15), .IN4(n97), .IN5(n96), 
        .Q(out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n17), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n16), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n16), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n18), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n17), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n19), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n18), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n18), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n20), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n19), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n21), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n20), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n20), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n21), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_64 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n33), .IN2(n7), .QN(n37) );
  NAND2X0 U4 ( .IN1(n41), .IN2(n8), .QN(n45) );
  NAND2X0 U5 ( .IN1(n49), .IN2(n9), .QN(n53) );
  NAND2X0 U6 ( .IN1(n57), .IN2(n10), .QN(n61) );
  NAND2X0 U7 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U8 ( .IN1(n25), .IN2(n6), .QN(n30) );
  NAND2X0 U9 ( .IN1(n65), .IN2(n11), .QN(n77) );
  NAND2X0 U10 ( .IN1(n81), .IN2(n13), .QN(n89) );
  NAND2X0 U11 ( .IN1(n93), .IN2(n15), .QN(n101) );
  NAND2X0 U12 ( .IN1(n118), .IN2(n19), .QN(n125) );
  NAND2X0 U13 ( .IN1(n105), .IN2(n17), .QN(n114) );
  NAND2X0 U14 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U15 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U16 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U17 ( .IN1(n40), .IN2(n39), .QN(out1[5]) );
  NAND2X0 U18 ( .IN1(n44), .IN2(n43), .QN(out1[6]) );
  NAND2X0 U19 ( .IN1(in1[2]), .IN2(n77), .QN(n71) );
  NAND2X0 U20 ( .IN1(n70), .IN2(n132), .QN(n74) );
  NAND2X0 U21 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U22 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U23 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U24 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U25 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U26 ( .IN1(n23), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U27 ( .IN1(in1[2]), .IN2(n22), .QN(n23) );
  NAND2X0 U28 ( .IN1(n36), .IN2(n35), .QN(out1[4]) );
  NAND2X0 U29 ( .IN1(n32), .IN2(n31), .QN(out1[3]) );
  NAND2X0 U30 ( .IN1(n27), .IN2(n132), .QN(n4) );
  NAND2X0 U31 ( .IN1(n48), .IN2(n47), .QN(out1[7]) );
  NAND2X0 U32 ( .IN1(n52), .IN2(n51), .QN(out1[8]) );
  NAND2X0 U33 ( .IN1(n56), .IN2(n55), .QN(out1[9]) );
  NAND2X0 U34 ( .IN1(n60), .IN2(n59), .QN(out1[10]) );
  NAND2X0 U35 ( .IN1(n64), .IN2(n63), .QN(out1[11]) );
  NAND2X0 U36 ( .IN1(n69), .IN2(n68), .QN(out1[12]) );
  NAND2X0 U37 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U38 ( .IN1(n141), .IN2(n130), .QN(n24) );
  NAND2X0 U39 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NOR2X0 U40 ( .IN1(n28), .IN2(n26), .QN(n3) );
  NOR2X0 U41 ( .IN1(n142), .IN2(n21), .QN(n1) );
  INVX0 U42 ( .INP(n132), .ZN(n141) );
  INVX0 U43 ( .INP(n130), .ZN(n137) );
  NAND3X0 U44 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  NOR3X0 U45 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  NOR2X0 U46 ( .IN1(n142), .IN2(n111), .QN(n138) );
  MUX21X1 U47 ( .IN1(n22), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  INVX0 U48 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U49 ( .INP(in2[2]), .ZN(n6) );
  INVX0 U50 ( .INP(in2[4]), .ZN(n7) );
  INVX0 U51 ( .INP(in2[6]), .ZN(n8) );
  INVX0 U52 ( .INP(in2[8]), .ZN(n9) );
  INVX0 U53 ( .INP(in2[10]), .ZN(n10) );
  INVX0 U54 ( .INP(in2[12]), .ZN(n11) );
  INVX0 U55 ( .INP(in2[13]), .ZN(n12) );
  INVX0 U56 ( .INP(in2[14]), .ZN(n13) );
  INVX0 U57 ( .INP(in2[15]), .ZN(n14) );
  INVX0 U58 ( .INP(in2[16]), .ZN(n15) );
  INVX0 U59 ( .INP(in2[17]), .ZN(n16) );
  INVX0 U60 ( .INP(in2[18]), .ZN(n17) );
  INVX0 U61 ( .INP(in2[19]), .ZN(n18) );
  INVX0 U62 ( .INP(in2[20]), .ZN(n19) );
  INVX0 U63 ( .INP(in2[21]), .ZN(n20) );
  INVX0 U64 ( .INP(in2[22]), .ZN(n21) );
  INVX0 U65 ( .INP(in1[1]), .ZN(n22) );
  INVX0 U66 ( .INP(in1[2]), .ZN(n111) );
  INVX0 U67 ( .INP(n138), .ZN(n140) );
  NOR2X0 U68 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n25) );
  AOI21X1 U69 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n25), .QN(n27) );
  NOR2X0 U70 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U71 ( .IN1(n24), .IN2(in2[0]), .IN3(n138), .IN4(n27), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U72 ( .INP(n133), .ZN(n67) );
  NOR2X0 U73 ( .IN1(n67), .IN2(n6), .QN(n28) );
  OA21X1 U74 ( .IN1(n25), .IN2(n6), .IN3(n30), .Q(n29) );
  AO22X1 U75 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n29), .Q(n26) );
  AOI22X1 U76 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n29), .QN(n32) );
  NOR2X0 U77 ( .IN1(in2[3]), .IN2(n30), .QN(n33) );
  AO21X1 U78 ( .IN1(in2[3]), .IN2(n30), .IN3(n33), .Q(n34) );
  OA22X1 U79 ( .IN1(n6), .IN2(n130), .IN3(n140), .IN4(n34), .Q(n31) );
  OA21X1 U80 ( .IN1(n33), .IN2(n7), .IN3(n37), .Q(n38) );
  AOI22X1 U81 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n38), .QN(n36) );
  OA22X1 U82 ( .IN1(n67), .IN2(n7), .IN3(n141), .IN4(n34), .Q(n35) );
  NOR2X0 U83 ( .IN1(in2[5]), .IN2(n37), .QN(n41) );
  AO21X1 U84 ( .IN1(in2[5]), .IN2(n37), .IN3(n41), .Q(n42) );
  OA22X1 U85 ( .IN1(n7), .IN2(n130), .IN3(n140), .IN4(n42), .Q(n40) );
  AOI22X1 U86 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n38), .QN(n39) );
  OA21X1 U87 ( .IN1(n41), .IN2(n8), .IN3(n45), .Q(n46) );
  AOI22X1 U88 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n46), .QN(n44) );
  OA22X1 U89 ( .IN1(n67), .IN2(n8), .IN3(n141), .IN4(n42), .Q(n43) );
  NOR2X0 U90 ( .IN1(in2[7]), .IN2(n45), .QN(n49) );
  AO21X1 U91 ( .IN1(in2[7]), .IN2(n45), .IN3(n49), .Q(n50) );
  OA22X1 U92 ( .IN1(n8), .IN2(n130), .IN3(n140), .IN4(n50), .Q(n48) );
  AOI22X1 U93 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n46), .QN(n47) );
  OA21X1 U94 ( .IN1(n49), .IN2(n9), .IN3(n53), .Q(n54) );
  AOI22X1 U95 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n54), .QN(n52) );
  OA22X1 U96 ( .IN1(n67), .IN2(n9), .IN3(n141), .IN4(n50), .Q(n51) );
  NOR2X0 U97 ( .IN1(in2[9]), .IN2(n53), .QN(n57) );
  AO21X1 U98 ( .IN1(in2[9]), .IN2(n53), .IN3(n57), .Q(n58) );
  OA22X1 U99 ( .IN1(n9), .IN2(n130), .IN3(n140), .IN4(n58), .Q(n56) );
  AOI22X1 U100 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n54), .QN(n55) );
  OA21X1 U101 ( .IN1(n57), .IN2(n10), .IN3(n61), .Q(n62) );
  AOI22X1 U102 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n62), .QN(n60) );
  OA22X1 U103 ( .IN1(n67), .IN2(n10), .IN3(n141), .IN4(n58), .Q(n59) );
  NOR2X0 U104 ( .IN1(in2[11]), .IN2(n61), .QN(n65) );
  AO21X1 U105 ( .IN1(in2[11]), .IN2(n61), .IN3(n65), .Q(n66) );
  OA22X1 U106 ( .IN1(n10), .IN2(n130), .IN3(n140), .IN4(n66), .Q(n64) );
  AOI22X1 U107 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n62), .QN(n63) );
  OA21X1 U108 ( .IN1(n65), .IN2(n11), .IN3(n77), .Q(n70) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n70), .QN(n69) );
  OA22X1 U110 ( .IN1(n67), .IN2(n11), .IN3(n141), .IN4(n66), .Q(n68) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n12), .S(n71), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n11), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n13), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n12), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n12), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n14), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n13), .IN4(n85), .IN5(n84), 
        .Q(out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n15), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n14), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n14), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n16), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n15), .IN4(n97), .IN5(n96), 
        .Q(out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n17), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n16), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n16), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n18), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n17), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n19), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n18), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n18), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n20), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n19), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n21), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n20), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n20), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n21), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_65 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93;

  NAND2X0 U3 ( .IN1(n30), .IN2(n7), .QN(n32) );
  NAND2X0 U4 ( .IN1(n34), .IN2(n8), .QN(n36) );
  NAND2X0 U5 ( .IN1(n38), .IN2(n9), .QN(n40) );
  NAND2X0 U6 ( .IN1(n42), .IN2(n10), .QN(n47) );
  NAND2X0 U7 ( .IN1(n78), .IN2(n18), .QN(n82) );
  NAND2X0 U8 ( .IN1(n26), .IN2(n6), .QN(n28) );
  NAND2X0 U9 ( .IN1(in1[2]), .IN2(n47), .QN(n44) );
  NAND2X0 U10 ( .IN1(n52), .IN2(n12), .QN(n55) );
  NAND2X0 U11 ( .IN1(in1[2]), .IN2(n55), .QN(n51) );
  NAND2X0 U12 ( .IN1(n60), .IN2(n14), .QN(n63) );
  NAND2X0 U13 ( .IN1(in1[2]), .IN2(n63), .QN(n59) );
  NAND2X0 U14 ( .IN1(n68), .IN2(n16), .QN(n71) );
  NAND2X0 U15 ( .IN1(in1[2]), .IN2(n71), .QN(n67) );
  NAND2X0 U16 ( .IN1(in1[2]), .IN2(n82), .QN(n77) );
  NAND2X0 U17 ( .IN1(in2[21]), .IN2(n82), .QN(n83) );
  NAND2X0 U18 ( .IN1(n75), .IN2(in1[2]), .QN(n86) );
  NAND2X0 U19 ( .IN1(n3), .IN2(n4), .QN(n22) );
  NAND2X0 U20 ( .IN1(in2[1]), .IN2(in2[0]), .QN(n4) );
  NAND2X0 U21 ( .IN1(n23), .IN2(n22), .QN(out1[2]) );
  INVX0 U22 ( .INP(n86), .ZN(n89) );
  NOR2X0 U23 ( .IN1(n21), .IN2(n86), .QN(n3) );
  NOR2X0 U24 ( .IN1(in1[2]), .IN2(n75), .QN(n90) );
  NOR2X0 U25 ( .IN1(n75), .IN2(n72), .QN(n92) );
  NBUFFX2 U26 ( .INP(in1[2]), .Z(out1[26]) );
  NBUFFX2 U27 ( .INP(in1[2]), .Z(out1[25]) );
  INVX0 U28 ( .INP(in2[2]), .ZN(n5) );
  INVX0 U29 ( .INP(in2[4]), .ZN(n6) );
  INVX0 U30 ( .INP(in2[6]), .ZN(n7) );
  INVX0 U31 ( .INP(in2[8]), .ZN(n8) );
  INVX0 U32 ( .INP(in2[10]), .ZN(n9) );
  INVX0 U33 ( .INP(in2[12]), .ZN(n10) );
  INVX0 U34 ( .INP(in2[13]), .ZN(n11) );
  INVX0 U35 ( .INP(in2[14]), .ZN(n12) );
  INVX0 U36 ( .INP(in2[15]), .ZN(n13) );
  INVX0 U37 ( .INP(in2[16]), .ZN(n14) );
  INVX0 U38 ( .INP(in2[17]), .ZN(n15) );
  INVX0 U39 ( .INP(in2[18]), .ZN(n16) );
  INVX0 U40 ( .INP(in2[19]), .ZN(n17) );
  INVX0 U41 ( .INP(in2[20]), .ZN(n18) );
  INVX0 U42 ( .INP(in2[21]), .ZN(n19) );
  INVX0 U43 ( .INP(in2[22]), .ZN(n20) );
  INVX0 U44 ( .INP(in1[1]), .ZN(n75) );
  INVX0 U45 ( .INP(in1[2]), .ZN(n72) );
  NOR2X0 U46 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n21) );
  OR3X1 U47 ( .IN1(in2[2]), .IN2(in2[0]), .IN3(in2[1]), .Q(n24) );
  OA21X1 U48 ( .IN1(n21), .IN2(n5), .IN3(n24), .Q(n25) );
  AOI22X1 U49 ( .IN1(in2[2]), .IN2(n90), .IN3(n92), .IN4(n25), .QN(n23) );
  NOR2X0 U50 ( .IN1(in2[3]), .IN2(n24), .QN(n26) );
  AOI21X1 U51 ( .IN1(in2[3]), .IN2(n24), .IN3(n26), .QN(n27) );
  AO222X1 U52 ( .IN1(in2[3]), .IN2(n90), .IN3(n92), .IN4(n27), .IN5(n89), 
        .IN6(n25), .Q(out1[3]) );
  OA21X1 U53 ( .IN1(n26), .IN2(n6), .IN3(n28), .Q(n29) );
  AO222X1 U54 ( .IN1(in2[4]), .IN2(n90), .IN3(n92), .IN4(n29), .IN5(n89), 
        .IN6(n27), .Q(out1[4]) );
  NOR2X0 U55 ( .IN1(in2[5]), .IN2(n28), .QN(n30) );
  AOI21X1 U56 ( .IN1(in2[5]), .IN2(n28), .IN3(n30), .QN(n31) );
  AO222X1 U57 ( .IN1(in2[5]), .IN2(n90), .IN3(n92), .IN4(n31), .IN5(n89), 
        .IN6(n29), .Q(out1[5]) );
  OA21X1 U58 ( .IN1(n30), .IN2(n7), .IN3(n32), .Q(n33) );
  AO222X1 U59 ( .IN1(in2[6]), .IN2(n90), .IN3(n92), .IN4(n33), .IN5(n89), 
        .IN6(n31), .Q(out1[6]) );
  NOR2X0 U60 ( .IN1(in2[7]), .IN2(n32), .QN(n34) );
  AOI21X1 U61 ( .IN1(in2[7]), .IN2(n32), .IN3(n34), .QN(n35) );
  AO222X1 U62 ( .IN1(in2[7]), .IN2(n90), .IN3(n92), .IN4(n35), .IN5(n89), 
        .IN6(n33), .Q(out1[7]) );
  OA21X1 U63 ( .IN1(n34), .IN2(n8), .IN3(n36), .Q(n37) );
  AO222X1 U64 ( .IN1(in2[8]), .IN2(n90), .IN3(n92), .IN4(n37), .IN5(n89), 
        .IN6(n35), .Q(out1[8]) );
  NOR2X0 U65 ( .IN1(in2[9]), .IN2(n36), .QN(n38) );
  AOI21X1 U66 ( .IN1(in2[9]), .IN2(n36), .IN3(n38), .QN(n39) );
  AO222X1 U67 ( .IN1(in2[9]), .IN2(n90), .IN3(n92), .IN4(n39), .IN5(n89), 
        .IN6(n37), .Q(out1[9]) );
  OA21X1 U68 ( .IN1(n38), .IN2(n9), .IN3(n40), .Q(n41) );
  AO222X1 U69 ( .IN1(in2[10]), .IN2(n90), .IN3(n92), .IN4(n41), .IN5(n89), 
        .IN6(n39), .Q(out1[10]) );
  NOR2X0 U70 ( .IN1(in2[11]), .IN2(n40), .QN(n42) );
  AOI21X1 U71 ( .IN1(in2[11]), .IN2(n40), .IN3(n42), .QN(n43) );
  AO222X1 U72 ( .IN1(in2[11]), .IN2(n90), .IN3(n92), .IN4(n43), .IN5(n89), 
        .IN6(n41), .Q(out1[11]) );
  OA21X1 U73 ( .IN1(n42), .IN2(n10), .IN3(n47), .Q(n45) );
  AO222X1 U74 ( .IN1(in2[12]), .IN2(n90), .IN3(n92), .IN4(n45), .IN5(n89), 
        .IN6(n43), .Q(out1[12]) );
  MUX21X1 U75 ( .IN1(n11), .IN2(in2[13]), .S(n44), .Q(n46) );
  AO22X1 U76 ( .IN1(in1[1]), .IN2(n46), .IN3(n89), .IN4(n45), .Q(out1[13]) );
  NOR2X0 U77 ( .IN1(in2[13]), .IN2(n47), .QN(n52) );
  AO21X1 U78 ( .IN1(in2[13]), .IN2(n47), .IN3(n86), .Q(n50) );
  NOR2X0 U79 ( .IN1(n52), .IN2(n72), .QN(n48) );
  MUX21X1 U80 ( .IN1(n12), .IN2(in2[14]), .S(n48), .Q(n49) );
  OAI22X1 U81 ( .IN1(n52), .IN2(n50), .IN3(n75), .IN4(n49), .QN(out1[14]) );
  MUX21X1 U82 ( .IN1(n13), .IN2(in2[15]), .S(n51), .Q(n54) );
  OA21X1 U83 ( .IN1(n52), .IN2(n12), .IN3(n89), .Q(n53) );
  AO22X1 U84 ( .IN1(in1[1]), .IN2(n54), .IN3(n53), .IN4(n55), .Q(out1[15]) );
  NOR2X0 U85 ( .IN1(in2[15]), .IN2(n55), .QN(n60) );
  AO21X1 U86 ( .IN1(in2[15]), .IN2(n55), .IN3(n86), .Q(n58) );
  NOR2X0 U87 ( .IN1(n60), .IN2(n72), .QN(n56) );
  MUX21X1 U88 ( .IN1(n14), .IN2(in2[16]), .S(n56), .Q(n57) );
  OAI22X1 U89 ( .IN1(n60), .IN2(n58), .IN3(n75), .IN4(n57), .QN(out1[16]) );
  MUX21X1 U90 ( .IN1(n15), .IN2(in2[17]), .S(n59), .Q(n62) );
  OA21X1 U91 ( .IN1(n60), .IN2(n14), .IN3(n89), .Q(n61) );
  AO22X1 U92 ( .IN1(in1[1]), .IN2(n62), .IN3(n61), .IN4(n63), .Q(out1[17]) );
  NOR2X0 U93 ( .IN1(in2[17]), .IN2(n63), .QN(n68) );
  AO21X1 U94 ( .IN1(in2[17]), .IN2(n63), .IN3(n86), .Q(n66) );
  NOR2X0 U95 ( .IN1(n68), .IN2(n72), .QN(n64) );
  MUX21X1 U96 ( .IN1(n16), .IN2(in2[18]), .S(n64), .Q(n65) );
  OAI22X1 U97 ( .IN1(n68), .IN2(n66), .IN3(n75), .IN4(n65), .QN(out1[18]) );
  MUX21X1 U98 ( .IN1(n17), .IN2(in2[19]), .S(n67), .Q(n70) );
  OA21X1 U99 ( .IN1(n68), .IN2(n16), .IN3(n89), .Q(n69) );
  AO22X1 U100 ( .IN1(in1[1]), .IN2(n70), .IN3(n69), .IN4(n71), .Q(out1[19]) );
  NOR2X0 U101 ( .IN1(in2[19]), .IN2(n71), .QN(n78) );
  AO21X1 U102 ( .IN1(in2[19]), .IN2(n71), .IN3(n86), .Q(n76) );
  NOR2X0 U103 ( .IN1(n78), .IN2(n72), .QN(n73) );
  MUX21X1 U104 ( .IN1(n18), .IN2(in2[20]), .S(n73), .Q(n74) );
  OAI22X1 U105 ( .IN1(n78), .IN2(n76), .IN3(n75), .IN4(n74), .QN(out1[20]) );
  MUX21X1 U106 ( .IN1(n19), .IN2(in2[21]), .S(n77), .Q(n80) );
  MUX21X1 U107 ( .IN1(n18), .IN2(in2[20]), .S(n78), .Q(n79) );
  AO22X1 U108 ( .IN1(in1[1]), .IN2(n80), .IN3(n89), .IN4(n79), .Q(out1[21]) );
  INVX0 U109 ( .INP(n92), .ZN(n81) );
  OR2X1 U110 ( .IN1(n82), .IN2(in2[21]), .Q(n88) );
  NOR2X0 U111 ( .IN1(n81), .IN2(n88), .QN(n87) );
  NOR2X0 U112 ( .IN1(in2[22]), .IN2(n81), .QN(n84) );
  OA221X1 U113 ( .IN1(n84), .IN2(n89), .IN3(n84), .IN4(n83), .IN5(n88), .Q(n85) );
  AO221X1 U114 ( .IN1(in2[22]), .IN2(n87), .IN3(in2[22]), .IN4(n90), .IN5(n85), 
        .Q(out1[22]) );
  NOR2X0 U115 ( .IN1(n86), .IN2(n88), .QN(n93) );
  AO21X1 U116 ( .IN1(n89), .IN2(n88), .IN3(n87), .Q(n91) );
  AO221X1 U117 ( .IN1(in2[22]), .IN2(n93), .IN3(n20), .IN4(n91), .IN5(n90), 
        .Q(out1[23]) );
  AO21X1 U118 ( .IN1(n93), .IN2(n20), .IN3(n92), .Q(out1[24]) );
endmodule


module mul26_5 ( clk, rst_n, in1, in2, en, mulout );
  input [25:0] in1;
  input [25:0] in2;
  output [50:0] mulout;
  input clk, rst_n, en;
  wire   N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24,
         N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38,
         N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N62, N63,
         N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77,
         N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91,
         N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n131, n132, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22,
         SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24,
         SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26,
         SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28,
         SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30,
         SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32,
         SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34,
         SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36,
         SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38,
         SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40,
         SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42,
         SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44,
         SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46,
         SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48,
         SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50,
         SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52,
         SYNOPSYS_UNCONNECTED_53, SYNOPSYS_UNCONNECTED_54,
         SYNOPSYS_UNCONNECTED_55, SYNOPSYS_UNCONNECTED_56,
         SYNOPSYS_UNCONNECTED_57, SYNOPSYS_UNCONNECTED_58,
         SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_60,
         SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_62,
         SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_64,
         SYNOPSYS_UNCONNECTED_65, SYNOPSYS_UNCONNECTED_66,
         SYNOPSYS_UNCONNECTED_67, SYNOPSYS_UNCONNECTED_68,
         SYNOPSYS_UNCONNECTED_69, SYNOPSYS_UNCONNECTED_70,
         SYNOPSYS_UNCONNECTED_71, SYNOPSYS_UNCONNECTED_72,
         SYNOPSYS_UNCONNECTED_73, SYNOPSYS_UNCONNECTED_74,
         SYNOPSYS_UNCONNECTED_75, SYNOPSYS_UNCONNECTED_76,
         SYNOPSYS_UNCONNECTED_77, SYNOPSYS_UNCONNECTED_78,
         SYNOPSYS_UNCONNECTED_79, SYNOPSYS_UNCONNECTED_80,
         SYNOPSYS_UNCONNECTED_81, SYNOPSYS_UNCONNECTED_82,
         SYNOPSYS_UNCONNECTED_83, SYNOPSYS_UNCONNECTED_84,
         SYNOPSYS_UNCONNECTED_85, SYNOPSYS_UNCONNECTED_86,
         SYNOPSYS_UNCONNECTED_87, SYNOPSYS_UNCONNECTED_88,
         SYNOPSYS_UNCONNECTED_89, SYNOPSYS_UNCONNECTED_90,
         SYNOPSYS_UNCONNECTED_91, SYNOPSYS_UNCONNECTED_92,
         SYNOPSYS_UNCONNECTED_93, SYNOPSYS_UNCONNECTED_94,
         SYNOPSYS_UNCONNECTED_95, SYNOPSYS_UNCONNECTED_96,
         SYNOPSYS_UNCONNECTED_97, SYNOPSYS_UNCONNECTED_98,
         SYNOPSYS_UNCONNECTED_99, SYNOPSYS_UNCONNECTED_100,
         SYNOPSYS_UNCONNECTED_101, SYNOPSYS_UNCONNECTED_102,
         SYNOPSYS_UNCONNECTED_103, SYNOPSYS_UNCONNECTED_104,
         SYNOPSYS_UNCONNECTED_105, SYNOPSYS_UNCONNECTED_106,
         SYNOPSYS_UNCONNECTED_107, SYNOPSYS_UNCONNECTED_108,
         SYNOPSYS_UNCONNECTED_109, SYNOPSYS_UNCONNECTED_110,
         SYNOPSYS_UNCONNECTED_111, SYNOPSYS_UNCONNECTED_112,
         SYNOPSYS_UNCONNECTED_113, SYNOPSYS_UNCONNECTED_114,
         SYNOPSYS_UNCONNECTED_115, SYNOPSYS_UNCONNECTED_116,
         SYNOPSYS_UNCONNECTED_117, SYNOPSYS_UNCONNECTED_118,
         SYNOPSYS_UNCONNECTED_119, SYNOPSYS_UNCONNECTED_120,
         SYNOPSYS_UNCONNECTED_121, SYNOPSYS_UNCONNECTED_122,
         SYNOPSYS_UNCONNECTED_123, SYNOPSYS_UNCONNECTED_124,
         SYNOPSYS_UNCONNECTED_125, SYNOPSYS_UNCONNECTED_126,
         SYNOPSYS_UNCONNECTED_127, SYNOPSYS_UNCONNECTED_128,
         SYNOPSYS_UNCONNECTED_129, SYNOPSYS_UNCONNECTED_130,
         SYNOPSYS_UNCONNECTED_131, SYNOPSYS_UNCONNECTED_132,
         SYNOPSYS_UNCONNECTED_133, SYNOPSYS_UNCONNECTED_134,
         SYNOPSYS_UNCONNECTED_135, SYNOPSYS_UNCONNECTED_136,
         SYNOPSYS_UNCONNECTED_137, SYNOPSYS_UNCONNECTED_138,
         SYNOPSYS_UNCONNECTED_139, SYNOPSYS_UNCONNECTED_140,
         SYNOPSYS_UNCONNECTED_141, SYNOPSYS_UNCONNECTED_142,
         SYNOPSYS_UNCONNECTED_143, SYNOPSYS_UNCONNECTED_144,
         SYNOPSYS_UNCONNECTED_145, SYNOPSYS_UNCONNECTED_146,
         SYNOPSYS_UNCONNECTED_147, SYNOPSYS_UNCONNECTED_148,
         SYNOPSYS_UNCONNECTED_149, SYNOPSYS_UNCONNECTED_150,
         SYNOPSYS_UNCONNECTED_151, SYNOPSYS_UNCONNECTED_152,
         SYNOPSYS_UNCONNECTED_153, SYNOPSYS_UNCONNECTED_154,
         SYNOPSYS_UNCONNECTED_155, SYNOPSYS_UNCONNECTED_156,
         SYNOPSYS_UNCONNECTED_157, SYNOPSYS_UNCONNECTED_158,
         SYNOPSYS_UNCONNECTED_159, SYNOPSYS_UNCONNECTED_160,
         SYNOPSYS_UNCONNECTED_161, SYNOPSYS_UNCONNECTED_162,
         SYNOPSYS_UNCONNECTED_163, SYNOPSYS_UNCONNECTED_164,
         SYNOPSYS_UNCONNECTED_165, SYNOPSYS_UNCONNECTED_166,
         SYNOPSYS_UNCONNECTED_167, SYNOPSYS_UNCONNECTED_168,
         SYNOPSYS_UNCONNECTED_169, SYNOPSYS_UNCONNECTED_170,
         SYNOPSYS_UNCONNECTED_171, SYNOPSYS_UNCONNECTED_172,
         SYNOPSYS_UNCONNECTED_173, SYNOPSYS_UNCONNECTED_174,
         SYNOPSYS_UNCONNECTED_175, SYNOPSYS_UNCONNECTED_176,
         SYNOPSYS_UNCONNECTED_177, SYNOPSYS_UNCONNECTED_178,
         SYNOPSYS_UNCONNECTED_179, SYNOPSYS_UNCONNECTED_180,
         SYNOPSYS_UNCONNECTED_181, SYNOPSYS_UNCONNECTED_182,
         SYNOPSYS_UNCONNECTED_183, SYNOPSYS_UNCONNECTED_184,
         SYNOPSYS_UNCONNECTED_185, SYNOPSYS_UNCONNECTED_186,
         SYNOPSYS_UNCONNECTED_187, SYNOPSYS_UNCONNECTED_188,
         SYNOPSYS_UNCONNECTED_189, SYNOPSYS_UNCONNECTED_190,
         SYNOPSYS_UNCONNECTED_191, SYNOPSYS_UNCONNECTED_192,
         SYNOPSYS_UNCONNECTED_193, SYNOPSYS_UNCONNECTED_194,
         SYNOPSYS_UNCONNECTED_195, SYNOPSYS_UNCONNECTED_196,
         SYNOPSYS_UNCONNECTED_197, SYNOPSYS_UNCONNECTED_198,
         SYNOPSYS_UNCONNECTED_199, SYNOPSYS_UNCONNECTED_200,
         SYNOPSYS_UNCONNECTED_201, SYNOPSYS_UNCONNECTED_202,
         SYNOPSYS_UNCONNECTED_203, SYNOPSYS_UNCONNECTED_204,
         SYNOPSYS_UNCONNECTED_205, SYNOPSYS_UNCONNECTED_206,
         SYNOPSYS_UNCONNECTED_207, SYNOPSYS_UNCONNECTED_208,
         SYNOPSYS_UNCONNECTED_209, SYNOPSYS_UNCONNECTED_210,
         SYNOPSYS_UNCONNECTED_211, SYNOPSYS_UNCONNECTED_212,
         SYNOPSYS_UNCONNECTED_213, SYNOPSYS_UNCONNECTED_214,
         SYNOPSYS_UNCONNECTED_215, SYNOPSYS_UNCONNECTED_216,
         SYNOPSYS_UNCONNECTED_217, SYNOPSYS_UNCONNECTED_218,
         SYNOPSYS_UNCONNECTED_219, SYNOPSYS_UNCONNECTED_220,
         SYNOPSYS_UNCONNECTED_221, SYNOPSYS_UNCONNECTED_222,
         SYNOPSYS_UNCONNECTED_223, SYNOPSYS_UNCONNECTED_224,
         SYNOPSYS_UNCONNECTED_225, SYNOPSYS_UNCONNECTED_226,
         SYNOPSYS_UNCONNECTED_227, SYNOPSYS_UNCONNECTED_228,
         SYNOPSYS_UNCONNECTED_229, SYNOPSYS_UNCONNECTED_230,
         SYNOPSYS_UNCONNECTED_231, SYNOPSYS_UNCONNECTED_232,
         SYNOPSYS_UNCONNECTED_233, SYNOPSYS_UNCONNECTED_234,
         SYNOPSYS_UNCONNECTED_235, SYNOPSYS_UNCONNECTED_236,
         SYNOPSYS_UNCONNECTED_237, SYNOPSYS_UNCONNECTED_238,
         SYNOPSYS_UNCONNECTED_239, SYNOPSYS_UNCONNECTED_240,
         SYNOPSYS_UNCONNECTED_241, SYNOPSYS_UNCONNECTED_242,
         SYNOPSYS_UNCONNECTED_243, SYNOPSYS_UNCONNECTED_244,
         SYNOPSYS_UNCONNECTED_245, SYNOPSYS_UNCONNECTED_246,
         SYNOPSYS_UNCONNECTED_247, SYNOPSYS_UNCONNECTED_248,
         SYNOPSYS_UNCONNECTED_249, SYNOPSYS_UNCONNECTED_250,
         SYNOPSYS_UNCONNECTED_251, SYNOPSYS_UNCONNECTED_252,
         SYNOPSYS_UNCONNECTED_253, SYNOPSYS_UNCONNECTED_254,
         SYNOPSYS_UNCONNECTED_255, SYNOPSYS_UNCONNECTED_256,
         SYNOPSYS_UNCONNECTED_257, SYNOPSYS_UNCONNECTED_258,
         SYNOPSYS_UNCONNECTED_259, SYNOPSYS_UNCONNECTED_260,
         SYNOPSYS_UNCONNECTED_261, SYNOPSYS_UNCONNECTED_262,
         SYNOPSYS_UNCONNECTED_263, SYNOPSYS_UNCONNECTED_264,
         SYNOPSYS_UNCONNECTED_265, SYNOPSYS_UNCONNECTED_266,
         SYNOPSYS_UNCONNECTED_267, SYNOPSYS_UNCONNECTED_268,
         SYNOPSYS_UNCONNECTED_269, SYNOPSYS_UNCONNECTED_270,
         SYNOPSYS_UNCONNECTED_271, SYNOPSYS_UNCONNECTED_272,
         SYNOPSYS_UNCONNECTED_273, SYNOPSYS_UNCONNECTED_274,
         SYNOPSYS_UNCONNECTED_275, SYNOPSYS_UNCONNECTED_276,
         SYNOPSYS_UNCONNECTED_277, SYNOPSYS_UNCONNECTED_278,
         SYNOPSYS_UNCONNECTED_279, SYNOPSYS_UNCONNECTED_280,
         SYNOPSYS_UNCONNECTED_281, SYNOPSYS_UNCONNECTED_282,
         SYNOPSYS_UNCONNECTED_283, SYNOPSYS_UNCONNECTED_284,
         SYNOPSYS_UNCONNECTED_285, SYNOPSYS_UNCONNECTED_286,
         SYNOPSYS_UNCONNECTED_287, SYNOPSYS_UNCONNECTED_288,
         SYNOPSYS_UNCONNECTED_289, SYNOPSYS_UNCONNECTED_290,
         SYNOPSYS_UNCONNECTED_291, SYNOPSYS_UNCONNECTED_292,
         SYNOPSYS_UNCONNECTED_293, SYNOPSYS_UNCONNECTED_294,
         SYNOPSYS_UNCONNECTED_295, SYNOPSYS_UNCONNECTED_296,
         SYNOPSYS_UNCONNECTED_297, SYNOPSYS_UNCONNECTED_298,
         SYNOPSYS_UNCONNECTED_299, SYNOPSYS_UNCONNECTED_300,
         SYNOPSYS_UNCONNECTED_301, SYNOPSYS_UNCONNECTED_302,
         SYNOPSYS_UNCONNECTED_303, SYNOPSYS_UNCONNECTED_304,
         SYNOPSYS_UNCONNECTED_305, SYNOPSYS_UNCONNECTED_306,
         SYNOPSYS_UNCONNECTED_307, SYNOPSYS_UNCONNECTED_308,
         SYNOPSYS_UNCONNECTED_309, SYNOPSYS_UNCONNECTED_310,
         SYNOPSYS_UNCONNECTED_311, SYNOPSYS_UNCONNECTED_312,
         SYNOPSYS_UNCONNECTED_313, SYNOPSYS_UNCONNECTED_314,
         SYNOPSYS_UNCONNECTED_315, SYNOPSYS_UNCONNECTED_316,
         SYNOPSYS_UNCONNECTED_317, SYNOPSYS_UNCONNECTED_318,
         SYNOPSYS_UNCONNECTED_319, SYNOPSYS_UNCONNECTED_320,
         SYNOPSYS_UNCONNECTED_321, SYNOPSYS_UNCONNECTED_322,
         SYNOPSYS_UNCONNECTED_323, SYNOPSYS_UNCONNECTED_324,
         SYNOPSYS_UNCONNECTED_325, SYNOPSYS_UNCONNECTED_326,
         SYNOPSYS_UNCONNECTED_327, SYNOPSYS_UNCONNECTED_328,
         SYNOPSYS_UNCONNECTED_329, SYNOPSYS_UNCONNECTED_330,
         SYNOPSYS_UNCONNECTED_331, SYNOPSYS_UNCONNECTED_332,
         SYNOPSYS_UNCONNECTED_333, SYNOPSYS_UNCONNECTED_334,
         SYNOPSYS_UNCONNECTED_335, SYNOPSYS_UNCONNECTED_336,
         SYNOPSYS_UNCONNECTED_337, SYNOPSYS_UNCONNECTED_338,
         SYNOPSYS_UNCONNECTED_339, SYNOPSYS_UNCONNECTED_340,
         SYNOPSYS_UNCONNECTED_341, SYNOPSYS_UNCONNECTED_342,
         SYNOPSYS_UNCONNECTED_343, SYNOPSYS_UNCONNECTED_344,
         SYNOPSYS_UNCONNECTED_345, SYNOPSYS_UNCONNECTED_346,
         SYNOPSYS_UNCONNECTED_347, SYNOPSYS_UNCONNECTED_348,
         SYNOPSYS_UNCONNECTED_349, SYNOPSYS_UNCONNECTED_350,
         SYNOPSYS_UNCONNECTED_351, SYNOPSYS_UNCONNECTED_352,
         SYNOPSYS_UNCONNECTED_353, SYNOPSYS_UNCONNECTED_354,
         SYNOPSYS_UNCONNECTED_355, SYNOPSYS_UNCONNECTED_356,
         SYNOPSYS_UNCONNECTED_357, SYNOPSYS_UNCONNECTED_358,
         SYNOPSYS_UNCONNECTED_359, SYNOPSYS_UNCONNECTED_360,
         SYNOPSYS_UNCONNECTED_361, SYNOPSYS_UNCONNECTED_362,
         SYNOPSYS_UNCONNECTED_363, SYNOPSYS_UNCONNECTED_364,
         SYNOPSYS_UNCONNECTED_365, SYNOPSYS_UNCONNECTED_366,
         SYNOPSYS_UNCONNECTED_367, SYNOPSYS_UNCONNECTED_368,
         SYNOPSYS_UNCONNECTED_369, SYNOPSYS_UNCONNECTED_370,
         SYNOPSYS_UNCONNECTED_371, SYNOPSYS_UNCONNECTED_372,
         SYNOPSYS_UNCONNECTED_373, SYNOPSYS_UNCONNECTED_374,
         SYNOPSYS_UNCONNECTED_375, SYNOPSYS_UNCONNECTED_376,
         SYNOPSYS_UNCONNECTED_377, SYNOPSYS_UNCONNECTED_378,
         SYNOPSYS_UNCONNECTED_379, SYNOPSYS_UNCONNECTED_380,
         SYNOPSYS_UNCONNECTED_381, SYNOPSYS_UNCONNECTED_382,
         SYNOPSYS_UNCONNECTED_383, SYNOPSYS_UNCONNECTED_384,
         SYNOPSYS_UNCONNECTED_385, SYNOPSYS_UNCONNECTED_386,
         SYNOPSYS_UNCONNECTED_387, SYNOPSYS_UNCONNECTED_388,
         SYNOPSYS_UNCONNECTED_389, SYNOPSYS_UNCONNECTED_390,
         SYNOPSYS_UNCONNECTED_391, SYNOPSYS_UNCONNECTED_392,
         SYNOPSYS_UNCONNECTED_393, SYNOPSYS_UNCONNECTED_394,
         SYNOPSYS_UNCONNECTED_395, SYNOPSYS_UNCONNECTED_396,
         SYNOPSYS_UNCONNECTED_397, SYNOPSYS_UNCONNECTED_398,
         SYNOPSYS_UNCONNECTED_399, SYNOPSYS_UNCONNECTED_400,
         SYNOPSYS_UNCONNECTED_401, SYNOPSYS_UNCONNECTED_402,
         SYNOPSYS_UNCONNECTED_403, SYNOPSYS_UNCONNECTED_404,
         SYNOPSYS_UNCONNECTED_405, SYNOPSYS_UNCONNECTED_406,
         SYNOPSYS_UNCONNECTED_407, SYNOPSYS_UNCONNECTED_408,
         SYNOPSYS_UNCONNECTED_409, SYNOPSYS_UNCONNECTED_410,
         SYNOPSYS_UNCONNECTED_411, SYNOPSYS_UNCONNECTED_412;
  wire   [26:2] boothout1;
  wire   [26:0] boothout2;
  wire   [26:0] boothout3;
  wire   [26:0] boothout4;
  wire   [26:0] boothout5;
  wire   [26:0] boothout6;
  wire   [26:0] boothout7;
  wire   [26:0] boothout8;
  wire   [26:0] boothout9;
  wire   [26:0] boothout10;
  wire   [26:0] boothout11;
  wire   [25:0] boothout12;
  wire   [22:0] boothout13;
  wire   [29:2] cout1;
  wire   [31:3] mulout1;
  wire   [35:8] cout2;
  wire   [37:6] mulout2;
  wire   [41:14] cout3;
  wire   [42:12] mulout3;
  wire   [46:20] cout4;
  wire   [47:18] mulout4;
  wire   [31:3] cout5;
  wire   [46:4] mulout5;
  wire   [37:9] cout6;
  wire   [42:6] mulout6;
  wire   [46:18] cout7;
  wire   [47:12] mulout7;
  wire   [38:4] cout8;
  wire   [46:5] mulout8;
  wire   [46:12] cout9;
  wire   [47:6] mulout9;
  wire   [46:5] cout10;
  wire   [47:6] mulout10;
  wire   [46:6] cout11;
  wire   [47:7] mulout11;
  wire   [47:0] a;
  wire   [47:8] b;

  booth27_65 booth1 ( .out1({boothout1, SYNOPSYS_UNCONNECTED_1, 
        SYNOPSYS_UNCONNECTED_2}), .in1({in1[1:0], 1'b0}), .in2({1'b0, 1'b0, 
        1'b1, n34, n33, n32, n31, n30, n29, n28, n27, n26, n25, in2[12], n24, 
        in2[10], n23, in2[8], n21, in2[6], n20, in2[4], n19, in2[2], n18, n17}) );
  booth27_64 booth2 ( .out1(boothout2), .in1(in1[3:1]), .in2({1'b0, 1'b0, 1'b1, 
        n34, n33, n32, n31, n30, n29, n28, n27, n26, n25, in2[12], n24, 
        in2[10], n23, in2[8], n21, in2[6], n20, in2[4], n19, in2[2], n18, n17}) );
  booth27_63 booth3 ( .out1(boothout3), .in1(in1[5:3]), .in2({1'b0, 1'b0, 1'b1, 
        n34, n33, n32, n31, n30, n29, n28, n27, n26, n25, in2[12], n24, 
        in2[10], n23, in2[8], n21, in2[6], n20, in2[4], n19, in2[2], n18, n17}) );
  booth27_62 booth4 ( .out1(boothout4), .in1(in1[7:5]), .in2({1'b0, 1'b0, 1'b1, 
        n34, n33, n32, n31, n30, n29, n28, n27, n26, n25, in2[12], n24, 
        in2[10], n23, in2[8], n21, in2[6], n20, in2[4], n19, in2[2], n18, n17}) );
  booth27_61 booth5 ( .out1(boothout5), .in1(in1[9:7]), .in2({1'b0, 1'b0, 1'b1, 
        n34, n33, n32, n31, n30, n29, n28, n27, n26, n25, in2[12], n24, 
        in2[10], n23, in2[8], n21, in2[6], n20, in2[4], n19, in2[2], n18, n17}) );
  booth27_60 booth6 ( .out1(boothout6), .in1(in1[11:9]), .in2({1'b0, 1'b0, 
        1'b1, n34, n33, n32, n31, n30, n29, n28, n27, n26, n25, in2[12], n24, 
        in2[10], n23, in2[8], n21, in2[6], n20, in2[4], n19, in2[2], n18, n17}) );
  booth27_59 booth7 ( .out1(boothout7), .in1(in1[13:11]), .in2({1'b0, 1'b0, 
        1'b1, n34, n33, n32, n31, n30, n29, n28, n27, n26, n25, in2[12], n24, 
        in2[10], n23, in2[8], n21, in2[6], n20, in2[4], n19, in2[2], n18, n17}) );
  booth27_58 booth8 ( .out1(boothout8), .in1(in1[15:13]), .in2({1'b0, 1'b0, 
        1'b1, n34, n33, n32, n31, n30, n29, n28, n27, n26, n25, in2[12], n24, 
        in2[10], n23, in2[8], n21, in2[6], n20, in2[4], n19, in2[2], n18, n17}) );
  booth27_57 booth9 ( .out1(boothout9), .in1(in1[17:15]), .in2({1'b0, 1'b0, 
        1'b1, n34, n33, n32, n31, n30, n29, n28, n27, n26, n25, in2[12], n24, 
        in2[10], n23, in2[8], n21, in2[6], n20, in2[4], n19, in2[2], n18, n17}) );
  booth27_56 booth10 ( .out1(boothout10), .in1(in1[19:17]), .in2({1'b0, 1'b0, 
        1'b1, n34, n33, n32, n31, n30, n29, n28, n27, n26, n25, in2[12], n24, 
        in2[10], n23, in2[8], n21, in2[6], n20, in2[4], n19, in2[2], n18, n17}) );
  booth27_55 booth11 ( .out1(boothout11), .in1(in1[21:19]), .in2({1'b0, 1'b0, 
        1'b1, n34, n33, n32, n31, n30, n29, n28, n27, n26, n25, in2[12], n24, 
        in2[10], n23, in2[8], n21, in2[6], n20, in2[4], n19, in2[2], n18, n17}) );
  booth27_54 booth12 ( .out1({SYNOPSYS_UNCONNECTED_3, boothout12}), .in1({1'b1, 
        in1[22:21]}), .in2({1'b0, 1'b0, 1'b1, n34, n33, n32, n31, n30, n29, 
        n28, n27, n26, n25, in2[12], n24, in2[10], n23, in2[8], n21, in2[6], 
        n20, in2[4], n19, in2[2], n18, n17}) );
  booth27_53 booth13 ( .out1({SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, 
        SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, boothout13}), .in1({
        1'b0, 1'b0, 1'b1}), .in2({1'b0, 1'b0, 1'b1, n34, n33, n32, n31, n30, 
        n29, n28, n27, n26, n25, in2[12], n24, in2[10], n23, in2[8], n21, 
        in2[6], n20, in2[4], n19, in2[2], n18, n17}) );
  csa51squ_60 csa51squ1 ( .cout({SYNOPSYS_UNCONNECTED_8, 
        SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10, 
        SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12, 
        SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14, 
        SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16, 
        SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18, 
        SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20, 
        SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22, 
        SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24, 
        SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26, 
        SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28, cout1, 
        SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30}), .sumout({
        SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32, 
        SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34, 
        SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36, 
        SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38, 
        SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40, 
        SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42, 
        SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44, 
        SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46, 
        SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48, 
        SYNOPSYS_UNCONNECTED_49, mulout1[31], SYNOPSYS_UNCONNECTED_50, 
        mulout1[29:3], SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52, 
        SYNOPSYS_UNCONNECTED_53}), .in1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, boothout1, 1'b0, 1'b0}), .in2({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, boothout2, 
        1'b0, 1'b0}), .in3({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n132, 
        1'b0, boothout3[25:0], 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_59 csa51squ2 ( .cout({SYNOPSYS_UNCONNECTED_54, 
        SYNOPSYS_UNCONNECTED_55, SYNOPSYS_UNCONNECTED_56, 
        SYNOPSYS_UNCONNECTED_57, SYNOPSYS_UNCONNECTED_58, 
        SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_60, 
        SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_62, 
        SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_64, 
        SYNOPSYS_UNCONNECTED_65, SYNOPSYS_UNCONNECTED_66, 
        SYNOPSYS_UNCONNECTED_67, SYNOPSYS_UNCONNECTED_68, cout2, 
        SYNOPSYS_UNCONNECTED_69, SYNOPSYS_UNCONNECTED_70, 
        SYNOPSYS_UNCONNECTED_71, SYNOPSYS_UNCONNECTED_72, 
        SYNOPSYS_UNCONNECTED_73, SYNOPSYS_UNCONNECTED_74, 
        SYNOPSYS_UNCONNECTED_75, SYNOPSYS_UNCONNECTED_76}), .sumout({
        SYNOPSYS_UNCONNECTED_77, SYNOPSYS_UNCONNECTED_78, 
        SYNOPSYS_UNCONNECTED_79, SYNOPSYS_UNCONNECTED_80, 
        SYNOPSYS_UNCONNECTED_81, SYNOPSYS_UNCONNECTED_82, 
        SYNOPSYS_UNCONNECTED_83, SYNOPSYS_UNCONNECTED_84, 
        SYNOPSYS_UNCONNECTED_85, SYNOPSYS_UNCONNECTED_86, 
        SYNOPSYS_UNCONNECTED_87, SYNOPSYS_UNCONNECTED_88, 
        SYNOPSYS_UNCONNECTED_89, mulout2[37], SYNOPSYS_UNCONNECTED_90, 
        mulout2[35:6], SYNOPSYS_UNCONNECTED_91, SYNOPSYS_UNCONNECTED_92, 
        SYNOPSYS_UNCONNECTED_93, SYNOPSYS_UNCONNECTED_94, 
        SYNOPSYS_UNCONNECTED_95, SYNOPSYS_UNCONNECTED_96}), .in1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, boothout4, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, boothout5, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .in3({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n131, 1'b0, boothout6[25:0], 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_58 csa51squ3 ( .cout({SYNOPSYS_UNCONNECTED_97, 
        SYNOPSYS_UNCONNECTED_98, SYNOPSYS_UNCONNECTED_99, 
        SYNOPSYS_UNCONNECTED_100, SYNOPSYS_UNCONNECTED_101, 
        SYNOPSYS_UNCONNECTED_102, SYNOPSYS_UNCONNECTED_103, 
        SYNOPSYS_UNCONNECTED_104, SYNOPSYS_UNCONNECTED_105, cout3, 
        SYNOPSYS_UNCONNECTED_106, SYNOPSYS_UNCONNECTED_107, 
        SYNOPSYS_UNCONNECTED_108, SYNOPSYS_UNCONNECTED_109, 
        SYNOPSYS_UNCONNECTED_110, SYNOPSYS_UNCONNECTED_111, 
        SYNOPSYS_UNCONNECTED_112, SYNOPSYS_UNCONNECTED_113, 
        SYNOPSYS_UNCONNECTED_114, SYNOPSYS_UNCONNECTED_115, 
        SYNOPSYS_UNCONNECTED_116, SYNOPSYS_UNCONNECTED_117, 
        SYNOPSYS_UNCONNECTED_118, SYNOPSYS_UNCONNECTED_119}), .sumout({
        SYNOPSYS_UNCONNECTED_120, SYNOPSYS_UNCONNECTED_121, 
        SYNOPSYS_UNCONNECTED_122, SYNOPSYS_UNCONNECTED_123, 
        SYNOPSYS_UNCONNECTED_124, SYNOPSYS_UNCONNECTED_125, 
        SYNOPSYS_UNCONNECTED_126, SYNOPSYS_UNCONNECTED_127, mulout3, 
        SYNOPSYS_UNCONNECTED_128, SYNOPSYS_UNCONNECTED_129, 
        SYNOPSYS_UNCONNECTED_130, SYNOPSYS_UNCONNECTED_131, 
        SYNOPSYS_UNCONNECTED_132, SYNOPSYS_UNCONNECTED_133, 
        SYNOPSYS_UNCONNECTED_134, SYNOPSYS_UNCONNECTED_135, 
        SYNOPSYS_UNCONNECTED_136, SYNOPSYS_UNCONNECTED_137, 
        SYNOPSYS_UNCONNECTED_138, SYNOPSYS_UNCONNECTED_139}), .in1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, boothout7, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, boothout8, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .in3({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        boothout9, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_57 csa51squ4 ( .cout({SYNOPSYS_UNCONNECTED_140, 
        SYNOPSYS_UNCONNECTED_141, SYNOPSYS_UNCONNECTED_142, 
        SYNOPSYS_UNCONNECTED_143, cout4, SYNOPSYS_UNCONNECTED_144, 
        SYNOPSYS_UNCONNECTED_145, SYNOPSYS_UNCONNECTED_146, 
        SYNOPSYS_UNCONNECTED_147, SYNOPSYS_UNCONNECTED_148, 
        SYNOPSYS_UNCONNECTED_149, SYNOPSYS_UNCONNECTED_150, 
        SYNOPSYS_UNCONNECTED_151, SYNOPSYS_UNCONNECTED_152, 
        SYNOPSYS_UNCONNECTED_153, SYNOPSYS_UNCONNECTED_154, 
        SYNOPSYS_UNCONNECTED_155, SYNOPSYS_UNCONNECTED_156, 
        SYNOPSYS_UNCONNECTED_157, SYNOPSYS_UNCONNECTED_158, 
        SYNOPSYS_UNCONNECTED_159, SYNOPSYS_UNCONNECTED_160, 
        SYNOPSYS_UNCONNECTED_161, SYNOPSYS_UNCONNECTED_162, 
        SYNOPSYS_UNCONNECTED_163}), .sumout({SYNOPSYS_UNCONNECTED_164, 
        SYNOPSYS_UNCONNECTED_165, SYNOPSYS_UNCONNECTED_166, mulout4, 
        SYNOPSYS_UNCONNECTED_167, SYNOPSYS_UNCONNECTED_168, 
        SYNOPSYS_UNCONNECTED_169, SYNOPSYS_UNCONNECTED_170, 
        SYNOPSYS_UNCONNECTED_171, SYNOPSYS_UNCONNECTED_172, 
        SYNOPSYS_UNCONNECTED_173, SYNOPSYS_UNCONNECTED_174, 
        SYNOPSYS_UNCONNECTED_175, SYNOPSYS_UNCONNECTED_176, 
        SYNOPSYS_UNCONNECTED_177, SYNOPSYS_UNCONNECTED_178, 
        SYNOPSYS_UNCONNECTED_179, SYNOPSYS_UNCONNECTED_180, 
        SYNOPSYS_UNCONNECTED_181, SYNOPSYS_UNCONNECTED_182, 
        SYNOPSYS_UNCONNECTED_183, SYNOPSYS_UNCONNECTED_184}), .in1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, boothout10, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 1'b0, 1'b0, 1'b0, boothout11, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .in3({1'b0, 1'b0, 1'b0, boothout12, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_56 csa51squ5 ( .cout({SYNOPSYS_UNCONNECTED_185, 
        SYNOPSYS_UNCONNECTED_186, SYNOPSYS_UNCONNECTED_187, 
        SYNOPSYS_UNCONNECTED_188, SYNOPSYS_UNCONNECTED_189, 
        SYNOPSYS_UNCONNECTED_190, SYNOPSYS_UNCONNECTED_191, 
        SYNOPSYS_UNCONNECTED_192, SYNOPSYS_UNCONNECTED_193, 
        SYNOPSYS_UNCONNECTED_194, SYNOPSYS_UNCONNECTED_195, 
        SYNOPSYS_UNCONNECTED_196, SYNOPSYS_UNCONNECTED_197, 
        SYNOPSYS_UNCONNECTED_198, SYNOPSYS_UNCONNECTED_199, 
        SYNOPSYS_UNCONNECTED_200, SYNOPSYS_UNCONNECTED_201, 
        SYNOPSYS_UNCONNECTED_202, SYNOPSYS_UNCONNECTED_203, cout5, 
        SYNOPSYS_UNCONNECTED_204, SYNOPSYS_UNCONNECTED_205, 
        SYNOPSYS_UNCONNECTED_206}), .sumout({SYNOPSYS_UNCONNECTED_207, 
        SYNOPSYS_UNCONNECTED_208, SYNOPSYS_UNCONNECTED_209, 
        SYNOPSYS_UNCONNECTED_210, mulout5, SYNOPSYS_UNCONNECTED_211, 
        SYNOPSYS_UNCONNECTED_212, SYNOPSYS_UNCONNECTED_213, 
        SYNOPSYS_UNCONNECTED_214}), .in1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, cout1, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, mulout1[31], 1'b0, mulout1[29:3], 1'b0, 1'b0, 1'b0}), 
        .in3({1'b0, 1'b0, 1'b0, 1'b1, boothout13, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_55 csa51squ6 ( .cout({SYNOPSYS_UNCONNECTED_215, 
        SYNOPSYS_UNCONNECTED_216, SYNOPSYS_UNCONNECTED_217, 
        SYNOPSYS_UNCONNECTED_218, SYNOPSYS_UNCONNECTED_219, 
        SYNOPSYS_UNCONNECTED_220, SYNOPSYS_UNCONNECTED_221, 
        SYNOPSYS_UNCONNECTED_222, SYNOPSYS_UNCONNECTED_223, 
        SYNOPSYS_UNCONNECTED_224, SYNOPSYS_UNCONNECTED_225, 
        SYNOPSYS_UNCONNECTED_226, SYNOPSYS_UNCONNECTED_227, cout6, 
        SYNOPSYS_UNCONNECTED_228, SYNOPSYS_UNCONNECTED_229, 
        SYNOPSYS_UNCONNECTED_230, SYNOPSYS_UNCONNECTED_231, 
        SYNOPSYS_UNCONNECTED_232, SYNOPSYS_UNCONNECTED_233, 
        SYNOPSYS_UNCONNECTED_234, SYNOPSYS_UNCONNECTED_235, 
        SYNOPSYS_UNCONNECTED_236}), .sumout({SYNOPSYS_UNCONNECTED_237, 
        SYNOPSYS_UNCONNECTED_238, SYNOPSYS_UNCONNECTED_239, 
        SYNOPSYS_UNCONNECTED_240, SYNOPSYS_UNCONNECTED_241, 
        SYNOPSYS_UNCONNECTED_242, SYNOPSYS_UNCONNECTED_243, 
        SYNOPSYS_UNCONNECTED_244, mulout6, SYNOPSYS_UNCONNECTED_245, 
        SYNOPSYS_UNCONNECTED_246, SYNOPSYS_UNCONNECTED_247, 
        SYNOPSYS_UNCONNECTED_248, SYNOPSYS_UNCONNECTED_249, 
        SYNOPSYS_UNCONNECTED_250}), .in1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, cout2, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        mulout2[37], 1'b0, mulout2[35:6], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .in3({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, cout3, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  csa51squ_54 csa51squ7 ( .cout({SYNOPSYS_UNCONNECTED_251, 
        SYNOPSYS_UNCONNECTED_252, SYNOPSYS_UNCONNECTED_253, 
        SYNOPSYS_UNCONNECTED_254, cout7, SYNOPSYS_UNCONNECTED_255, 
        SYNOPSYS_UNCONNECTED_256, SYNOPSYS_UNCONNECTED_257, 
        SYNOPSYS_UNCONNECTED_258, SYNOPSYS_UNCONNECTED_259, 
        SYNOPSYS_UNCONNECTED_260, SYNOPSYS_UNCONNECTED_261, 
        SYNOPSYS_UNCONNECTED_262, SYNOPSYS_UNCONNECTED_263, 
        SYNOPSYS_UNCONNECTED_264, SYNOPSYS_UNCONNECTED_265, 
        SYNOPSYS_UNCONNECTED_266, SYNOPSYS_UNCONNECTED_267, 
        SYNOPSYS_UNCONNECTED_268, SYNOPSYS_UNCONNECTED_269, 
        SYNOPSYS_UNCONNECTED_270, SYNOPSYS_UNCONNECTED_271, 
        SYNOPSYS_UNCONNECTED_272}), .sumout({SYNOPSYS_UNCONNECTED_273, 
        SYNOPSYS_UNCONNECTED_274, SYNOPSYS_UNCONNECTED_275, mulout7, 
        SYNOPSYS_UNCONNECTED_276, SYNOPSYS_UNCONNECTED_277, 
        SYNOPSYS_UNCONNECTED_278, SYNOPSYS_UNCONNECTED_279, 
        SYNOPSYS_UNCONNECTED_280, SYNOPSYS_UNCONNECTED_281, 
        SYNOPSYS_UNCONNECTED_282, SYNOPSYS_UNCONNECTED_283, 
        SYNOPSYS_UNCONNECTED_284, SYNOPSYS_UNCONNECTED_285, 
        SYNOPSYS_UNCONNECTED_286, SYNOPSYS_UNCONNECTED_287}), .in1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mulout3, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 1'b0, 
        1'b0, cout4, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in3({1'b0, 1'b0, 1'b0, mulout4, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_53 csa51squ8 ( .cout({SYNOPSYS_UNCONNECTED_288, 
        SYNOPSYS_UNCONNECTED_289, SYNOPSYS_UNCONNECTED_290, 
        SYNOPSYS_UNCONNECTED_291, SYNOPSYS_UNCONNECTED_292, 
        SYNOPSYS_UNCONNECTED_293, SYNOPSYS_UNCONNECTED_294, 
        SYNOPSYS_UNCONNECTED_295, SYNOPSYS_UNCONNECTED_296, 
        SYNOPSYS_UNCONNECTED_297, SYNOPSYS_UNCONNECTED_298, 
        SYNOPSYS_UNCONNECTED_299, cout8, SYNOPSYS_UNCONNECTED_300, 
        SYNOPSYS_UNCONNECTED_301, SYNOPSYS_UNCONNECTED_302, 
        SYNOPSYS_UNCONNECTED_303}), .sumout({SYNOPSYS_UNCONNECTED_304, 
        SYNOPSYS_UNCONNECTED_305, SYNOPSYS_UNCONNECTED_306, 
        SYNOPSYS_UNCONNECTED_307, mulout8, SYNOPSYS_UNCONNECTED_308, 
        SYNOPSYS_UNCONNECTED_309, SYNOPSYS_UNCONNECTED_310, 
        SYNOPSYS_UNCONNECTED_311, SYNOPSYS_UNCONNECTED_312}), .in1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, cout5, 1'b0, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 
        1'b0, 1'b0, 1'b1, mulout5, 1'b0, 1'b0, 1'b0, 1'b0}), .in3({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, cout6, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_52 csa51squ9 ( .cout({SYNOPSYS_UNCONNECTED_313, 
        SYNOPSYS_UNCONNECTED_314, SYNOPSYS_UNCONNECTED_315, 
        SYNOPSYS_UNCONNECTED_316, cout9, SYNOPSYS_UNCONNECTED_317, 
        SYNOPSYS_UNCONNECTED_318, SYNOPSYS_UNCONNECTED_319, 
        SYNOPSYS_UNCONNECTED_320, SYNOPSYS_UNCONNECTED_321, 
        SYNOPSYS_UNCONNECTED_322, SYNOPSYS_UNCONNECTED_323, 
        SYNOPSYS_UNCONNECTED_324, SYNOPSYS_UNCONNECTED_325, 
        SYNOPSYS_UNCONNECTED_326, SYNOPSYS_UNCONNECTED_327, 
        SYNOPSYS_UNCONNECTED_328}), .sumout({SYNOPSYS_UNCONNECTED_329, 
        SYNOPSYS_UNCONNECTED_330, SYNOPSYS_UNCONNECTED_331, mulout9, 
        SYNOPSYS_UNCONNECTED_332, SYNOPSYS_UNCONNECTED_333, 
        SYNOPSYS_UNCONNECTED_334, SYNOPSYS_UNCONNECTED_335, 
        SYNOPSYS_UNCONNECTED_336, SYNOPSYS_UNCONNECTED_337}), .in1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mulout6, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .in2({1'b0, 1'b0, 1'b0, cout7, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .in3({1'b0, 1'b0, 1'b0, mulout7, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_51 csa51squ10 ( .cout({SYNOPSYS_UNCONNECTED_338, 
        SYNOPSYS_UNCONNECTED_339, SYNOPSYS_UNCONNECTED_340, 
        SYNOPSYS_UNCONNECTED_341, cout10, SYNOPSYS_UNCONNECTED_342, 
        SYNOPSYS_UNCONNECTED_343, SYNOPSYS_UNCONNECTED_344, 
        SYNOPSYS_UNCONNECTED_345, SYNOPSYS_UNCONNECTED_346}), .sumout({
        SYNOPSYS_UNCONNECTED_347, SYNOPSYS_UNCONNECTED_348, 
        SYNOPSYS_UNCONNECTED_349, mulout10, SYNOPSYS_UNCONNECTED_350, 
        SYNOPSYS_UNCONNECTED_351, SYNOPSYS_UNCONNECTED_352, 
        SYNOPSYS_UNCONNECTED_353, SYNOPSYS_UNCONNECTED_354, 
        SYNOPSYS_UNCONNECTED_355}), .in1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, cout8, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .in2({1'b0, 1'b0, 1'b0, 1'b1, mulout8, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .in3({1'b0, 1'b0, 1'b0, cout9, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_50 csa51squ11 ( .cout({SYNOPSYS_UNCONNECTED_356, 
        SYNOPSYS_UNCONNECTED_357, SYNOPSYS_UNCONNECTED_358, 
        SYNOPSYS_UNCONNECTED_359, cout11, SYNOPSYS_UNCONNECTED_360, 
        SYNOPSYS_UNCONNECTED_361, SYNOPSYS_UNCONNECTED_362, 
        SYNOPSYS_UNCONNECTED_363, SYNOPSYS_UNCONNECTED_364, 
        SYNOPSYS_UNCONNECTED_365}), .sumout({SYNOPSYS_UNCONNECTED_366, 
        SYNOPSYS_UNCONNECTED_367, SYNOPSYS_UNCONNECTED_368, mulout11, 
        SYNOPSYS_UNCONNECTED_369, SYNOPSYS_UNCONNECTED_370, 
        SYNOPSYS_UNCONNECTED_371, SYNOPSYS_UNCONNECTED_372, 
        SYNOPSYS_UNCONNECTED_373, SYNOPSYS_UNCONNECTED_374, 
        SYNOPSYS_UNCONNECTED_375}), .in1({1'b0, 1'b0, 1'b0, mulout9, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 1'b0, 1'b0, cout10, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in3({1'b0, 1'b0, 1'b0, mulout10, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_49 csa51squ12 ( .sumout({SYNOPSYS_UNCONNECTED_376, 
        SYNOPSYS_UNCONNECTED_377, SYNOPSYS_UNCONNECTED_378, N101, N100, N99, 
        N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, 
        N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, 
        N70, N69, N68, N67, N66, N65, N64, N63, N62, SYNOPSYS_UNCONNECTED_379, 
        SYNOPSYS_UNCONNECTED_380, SYNOPSYS_UNCONNECTED_381, 
        SYNOPSYS_UNCONNECTED_382, SYNOPSYS_UNCONNECTED_383, 
        SYNOPSYS_UNCONNECTED_384, SYNOPSYS_UNCONNECTED_385, 
        SYNOPSYS_UNCONNECTED_386}), .in1({1'b0, 1'b0, 1'b0, mulout11, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 1'b0, 1'b0, cout11, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in3({1'b1, 1'b0, 1'b1, 
        1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 
        1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .cout_46_(N50), .cout_44_(N48), .cout_42_(N46), .cout_40_(N44), .cout_38_(
        N42), .cout_36_(N40), .cout_34_(N38), .cout_32_(N36), .cout_30_(N34), 
        .cout_28_(N32), .cout_27_(N31), .cout_7__BAR(N11), .cout_8__BAR(N12), 
        .cout_9__BAR(N13), .cout_10__BAR(N14), .cout_11__BAR(N15), 
        .cout_12__BAR(N16), .cout_13__BAR(N17), .cout_14__BAR(N18), 
        .cout_15__BAR(N19), .cout_16__BAR(N20), .cout_17__BAR(N21), 
        .cout_18__BAR(N22), .cout_19__BAR(N23), .cout_20__BAR(N24), 
        .cout_21__BAR(N25), .cout_22__BAR(N26), .cout_23__BAR(N27), 
        .cout_24__BAR(N28), .cout_25__BAR(N29), .cout_26__BAR(N30), 
        .cout_29__BAR(N33), .cout_31__BAR(N35), .cout_33__BAR(N37), 
        .cout_35__BAR(N39), .cout_37__BAR(N41), .cout_39__BAR(N43), 
        .cout_41__BAR(N45), .cout_43__BAR(N47), .cout_45__BAR(N49) );
  cla51squ_5 cla51squ ( .out({SYNOPSYS_UNCONNECTED_387, 
        SYNOPSYS_UNCONNECTED_388, SYNOPSYS_UNCONNECTED_389, mulout[47:23], 
        SYNOPSYS_UNCONNECTED_390, SYNOPSYS_UNCONNECTED_391, 
        SYNOPSYS_UNCONNECTED_392, SYNOPSYS_UNCONNECTED_393, 
        SYNOPSYS_UNCONNECTED_394, SYNOPSYS_UNCONNECTED_395, 
        SYNOPSYS_UNCONNECTED_396, SYNOPSYS_UNCONNECTED_397, 
        SYNOPSYS_UNCONNECTED_398, SYNOPSYS_UNCONNECTED_399, 
        SYNOPSYS_UNCONNECTED_400, SYNOPSYS_UNCONNECTED_401, 
        SYNOPSYS_UNCONNECTED_402, SYNOPSYS_UNCONNECTED_403, 
        SYNOPSYS_UNCONNECTED_404, SYNOPSYS_UNCONNECTED_405, 
        SYNOPSYS_UNCONNECTED_406, SYNOPSYS_UNCONNECTED_407, 
        SYNOPSYS_UNCONNECTED_408, SYNOPSYS_UNCONNECTED_409, 
        SYNOPSYS_UNCONNECTED_410, SYNOPSYS_UNCONNECTED_411, 
        SYNOPSYS_UNCONNECTED_412}), .a({1'b0, 1'b0, 1'b0, a[47:8], 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({1'b0, 1'b0, 1'b0, b, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  DFFARX1 b_reg_47_ ( .D(N101), .CLK(clk), .RSTB(rst_n), .Q(b[47]) );
  DFFARX1 b_reg_46_ ( .D(N100), .CLK(clk), .RSTB(rst_n), .Q(b[46]) );
  DFFARX1 b_reg_45_ ( .D(N99), .CLK(clk), .RSTB(rst_n), .Q(b[45]) );
  DFFARX1 b_reg_44_ ( .D(N98), .CLK(clk), .RSTB(rst_n), .Q(b[44]) );
  DFFARX1 b_reg_43_ ( .D(N97), .CLK(clk), .RSTB(rst_n), .Q(b[43]) );
  DFFARX1 b_reg_42_ ( .D(N96), .CLK(clk), .RSTB(rst_n), .Q(b[42]) );
  DFFARX1 b_reg_41_ ( .D(N95), .CLK(clk), .RSTB(rst_n), .Q(b[41]) );
  DFFARX1 b_reg_40_ ( .D(N94), .CLK(clk), .RSTB(rst_n), .Q(b[40]) );
  DFFARX1 b_reg_39_ ( .D(N93), .CLK(clk), .RSTB(rst_n), .Q(b[39]) );
  DFFARX1 b_reg_38_ ( .D(N92), .CLK(clk), .RSTB(rst_n), .Q(b[38]) );
  DFFARX1 b_reg_37_ ( .D(N91), .CLK(clk), .RSTB(rst_n), .Q(b[37]) );
  DFFARX1 b_reg_36_ ( .D(N90), .CLK(clk), .RSTB(rst_n), .Q(b[36]) );
  DFFARX1 b_reg_35_ ( .D(N89), .CLK(clk), .RSTB(rst_n), .Q(b[35]) );
  DFFARX1 b_reg_34_ ( .D(N88), .CLK(clk), .RSTB(rst_n), .Q(b[34]) );
  DFFARX1 b_reg_33_ ( .D(N87), .CLK(clk), .RSTB(rst_n), .Q(b[33]) );
  DFFARX1 b_reg_32_ ( .D(N86), .CLK(clk), .RSTB(rst_n), .Q(b[32]) );
  DFFARX1 b_reg_31_ ( .D(N85), .CLK(clk), .RSTB(rst_n), .Q(b[31]) );
  DFFARX1 b_reg_30_ ( .D(N84), .CLK(clk), .RSTB(rst_n), .Q(b[30]) );
  DFFARX1 b_reg_29_ ( .D(N83), .CLK(clk), .RSTB(rst_n), .Q(b[29]) );
  DFFARX1 b_reg_28_ ( .D(N82), .CLK(clk), .RSTB(rst_n), .Q(b[28]) );
  DFFARX1 b_reg_27_ ( .D(N81), .CLK(clk), .RSTB(rst_n), .Q(b[27]) );
  DFFARX1 b_reg_26_ ( .D(N80), .CLK(clk), .RSTB(rst_n), .Q(b[26]) );
  DFFARX1 b_reg_25_ ( .D(N79), .CLK(clk), .RSTB(rst_n), .Q(b[25]) );
  DFFARX1 b_reg_24_ ( .D(N78), .CLK(clk), .RSTB(rst_n), .Q(b[24]) );
  DFFARX1 b_reg_23_ ( .D(N77), .CLK(clk), .RSTB(rst_n), .Q(b[23]) );
  DFFARX1 b_reg_22_ ( .D(N76), .CLK(clk), .RSTB(rst_n), .Q(b[22]) );
  DFFARX1 b_reg_21_ ( .D(N75), .CLK(clk), .RSTB(rst_n), .Q(b[21]) );
  DFFARX1 b_reg_20_ ( .D(N74), .CLK(clk), .RSTB(rst_n), .Q(b[20]) );
  DFFARX1 b_reg_19_ ( .D(N73), .CLK(clk), .RSTB(rst_n), .Q(b[19]) );
  DFFARX1 b_reg_18_ ( .D(N72), .CLK(clk), .RSTB(rst_n), .Q(b[18]) );
  DFFARX1 b_reg_17_ ( .D(N71), .CLK(clk), .RSTB(rst_n), .Q(b[17]) );
  DFFARX1 b_reg_16_ ( .D(N70), .CLK(clk), .RSTB(rst_n), .Q(b[16]) );
  DFFARX1 b_reg_15_ ( .D(N69), .CLK(clk), .RSTB(rst_n), .Q(b[15]) );
  DFFARX1 b_reg_14_ ( .D(N68), .CLK(clk), .RSTB(rst_n), .Q(b[14]) );
  DFFARX1 b_reg_13_ ( .D(N67), .CLK(clk), .RSTB(rst_n), .Q(b[13]) );
  DFFARX1 b_reg_12_ ( .D(N66), .CLK(clk), .RSTB(rst_n), .Q(b[12]) );
  DFFARX1 b_reg_11_ ( .D(N65), .CLK(clk), .RSTB(rst_n), .Q(b[11]) );
  DFFARX1 b_reg_10_ ( .D(N64), .CLK(clk), .RSTB(rst_n), .Q(b[10]) );
  DFFARX1 b_reg_9_ ( .D(N63), .CLK(clk), .RSTB(rst_n), .Q(b[9]) );
  DFFARX1 b_reg_8_ ( .D(N62), .CLK(clk), .RSTB(rst_n), .Q(b[8]) );
  DFFARX1 a_reg_47_ ( .D(N50), .CLK(clk), .RSTB(rst_n), .Q(a[47]) );
  DFFARX1 a_reg_46_ ( .D(n63), .CLK(clk), .RSTB(rst_n), .Q(a[46]) );
  DFFARX1 a_reg_45_ ( .D(N48), .CLK(clk), .RSTB(rst_n), .Q(a[45]) );
  DFFARX1 a_reg_44_ ( .D(n64), .CLK(clk), .RSTB(rst_n), .Q(a[44]) );
  DFFARX1 a_reg_43_ ( .D(N46), .CLK(clk), .RSTB(rst_n), .Q(a[43]) );
  DFFARX1 a_reg_42_ ( .D(n65), .CLK(clk), .RSTB(rst_n), .Q(a[42]) );
  DFFARX1 a_reg_41_ ( .D(N44), .CLK(clk), .RSTB(rst_n), .Q(a[41]) );
  DFFARX1 a_reg_40_ ( .D(n66), .CLK(clk), .RSTB(rst_n), .Q(a[40]) );
  DFFARX1 a_reg_39_ ( .D(N42), .CLK(clk), .RSTB(rst_n), .Q(a[39]) );
  DFFARX1 a_reg_38_ ( .D(n67), .CLK(clk), .RSTB(rst_n), .Q(a[38]) );
  DFFARX1 a_reg_37_ ( .D(N40), .CLK(clk), .RSTB(rst_n), .Q(a[37]) );
  DFFARX1 a_reg_36_ ( .D(n68), .CLK(clk), .RSTB(rst_n), .Q(a[36]) );
  DFFARX1 a_reg_35_ ( .D(N38), .CLK(clk), .RSTB(rst_n), .Q(a[35]) );
  DFFARX1 a_reg_34_ ( .D(n69), .CLK(clk), .RSTB(rst_n), .Q(a[34]) );
  DFFARX1 a_reg_33_ ( .D(N36), .CLK(clk), .RSTB(rst_n), .Q(a[33]) );
  DFFARX1 a_reg_32_ ( .D(n70), .CLK(clk), .RSTB(rst_n), .Q(a[32]) );
  DFFARX1 a_reg_31_ ( .D(N34), .CLK(clk), .RSTB(rst_n), .Q(a[31]) );
  DFFARX1 a_reg_30_ ( .D(n71), .CLK(clk), .RSTB(rst_n), .Q(a[30]) );
  DFFARX1 a_reg_29_ ( .D(N32), .CLK(clk), .RSTB(rst_n), .Q(a[29]) );
  DFFARX1 a_reg_28_ ( .D(N31), .CLK(clk), .RSTB(rst_n), .Q(a[28]) );
  DFFARX1 a_reg_27_ ( .D(n72), .CLK(clk), .RSTB(rst_n), .Q(a[27]) );
  DFFARX1 a_reg_26_ ( .D(n73), .CLK(clk), .RSTB(rst_n), .Q(a[26]) );
  DFFARX1 a_reg_25_ ( .D(n74), .CLK(clk), .RSTB(rst_n), .Q(a[25]) );
  DFFARX1 a_reg_24_ ( .D(n75), .CLK(clk), .RSTB(rst_n), .Q(a[24]) );
  DFFARX1 a_reg_23_ ( .D(n76), .CLK(clk), .RSTB(rst_n), .Q(a[23]) );
  DFFARX1 a_reg_22_ ( .D(n77), .CLK(clk), .RSTB(rst_n), .Q(a[22]) );
  DFFARX1 a_reg_21_ ( .D(n78), .CLK(clk), .RSTB(rst_n), .Q(a[21]) );
  DFFARX1 a_reg_20_ ( .D(n79), .CLK(clk), .RSTB(rst_n), .Q(a[20]) );
  DFFARX1 a_reg_19_ ( .D(n80), .CLK(clk), .RSTB(rst_n), .Q(a[19]) );
  DFFARX1 a_reg_18_ ( .D(n81), .CLK(clk), .RSTB(rst_n), .Q(a[18]) );
  DFFARX1 a_reg_17_ ( .D(n82), .CLK(clk), .RSTB(rst_n), .Q(a[17]) );
  DFFARX1 a_reg_16_ ( .D(n83), .CLK(clk), .RSTB(rst_n), .Q(a[16]) );
  DFFARX1 a_reg_15_ ( .D(n84), .CLK(clk), .RSTB(rst_n), .Q(a[15]) );
  DFFARX1 a_reg_14_ ( .D(n85), .CLK(clk), .RSTB(rst_n), .Q(a[14]) );
  DFFARX1 a_reg_13_ ( .D(n86), .CLK(clk), .RSTB(rst_n), .Q(a[13]) );
  DFFARX1 a_reg_12_ ( .D(n87), .CLK(clk), .RSTB(rst_n), .Q(a[12]) );
  DFFARX1 a_reg_11_ ( .D(n88), .CLK(clk), .RSTB(rst_n), .Q(a[11]) );
  DFFARX1 a_reg_10_ ( .D(n89), .CLK(clk), .RSTB(rst_n), .Q(a[10]) );
  DFFARX1 a_reg_9_ ( .D(n90), .CLK(clk), .RSTB(rst_n), .Q(a[9]) );
  DFFARX1 a_reg_8_ ( .D(n91), .CLK(clk), .RSTB(rst_n), .Q(a[8]) );
  INVX0 U5 ( .INP(boothout3[26]), .ZN(n132) );
  INVX0 U8 ( .INP(boothout6[26]), .ZN(n131) );
  NBUFFX8 U3 ( .INP(in2[15]), .Z(n27) );
  NBUFFX8 U4 ( .INP(in2[21]), .Z(n33) );
  NBUFFX8 U6 ( .INP(in2[22]), .Z(n34) );
  NBUFFX8 U7 ( .INP(in2[18]), .Z(n30) );
  NBUFFX8 U9 ( .INP(in2[14]), .Z(n26) );
  NBUFFX8 U10 ( .INP(in2[16]), .Z(n28) );
  NBUFFX8 U11 ( .INP(in2[20]), .Z(n32) );
  NBUFFX8 U12 ( .INP(in2[19]), .Z(n31) );
  NBUFFX8 U13 ( .INP(in2[17]), .Z(n29) );
  NBUFFX8 U14 ( .INP(in2[13]), .Z(n25) );
  NBUFFX8 U15 ( .INP(in2[3]), .Z(n19) );
  NBUFFX8 U16 ( .INP(in2[5]), .Z(n20) );
  NBUFFX8 U17 ( .INP(in2[9]), .Z(n23) );
  NBUFFX8 U18 ( .INP(in2[11]), .Z(n24) );
  INVX0 U19 ( .INP(n22), .ZN(n21) );
  NBUFFX8 U20 ( .INP(in2[1]), .Z(n18) );
  NBUFFX8 U21 ( .INP(in2[0]), .Z(n17) );
  INVX0 U36 ( .INP(in2[7]), .ZN(n22) );
  INVX0 U72 ( .INP(N49), .ZN(n63) );
  INVX0 U73 ( .INP(N47), .ZN(n64) );
  INVX0 U74 ( .INP(N45), .ZN(n65) );
  INVX0 U75 ( .INP(N43), .ZN(n66) );
  INVX0 U76 ( .INP(N41), .ZN(n67) );
  INVX0 U77 ( .INP(N39), .ZN(n68) );
  INVX0 U78 ( .INP(N37), .ZN(n69) );
  INVX0 U79 ( .INP(N35), .ZN(n70) );
  INVX0 U80 ( .INP(N33), .ZN(n71) );
  INVX0 U81 ( .INP(N30), .ZN(n72) );
  INVX0 U82 ( .INP(N29), .ZN(n73) );
  INVX0 U83 ( .INP(N28), .ZN(n74) );
  INVX0 U84 ( .INP(N27), .ZN(n75) );
  INVX0 U85 ( .INP(N26), .ZN(n76) );
  INVX0 U86 ( .INP(N25), .ZN(n77) );
  INVX0 U87 ( .INP(N24), .ZN(n78) );
  INVX0 U88 ( .INP(N23), .ZN(n79) );
  INVX0 U89 ( .INP(N22), .ZN(n80) );
  INVX0 U90 ( .INP(N21), .ZN(n81) );
  INVX0 U91 ( .INP(N20), .ZN(n82) );
  INVX0 U92 ( .INP(N19), .ZN(n83) );
  INVX0 U93 ( .INP(N18), .ZN(n84) );
  INVX0 U94 ( .INP(N17), .ZN(n85) );
  INVX0 U95 ( .INP(N16), .ZN(n86) );
  INVX0 U96 ( .INP(N15), .ZN(n87) );
  INVX0 U97 ( .INP(N14), .ZN(n88) );
  INVX0 U98 ( .INP(N13), .ZN(n89) );
  INVX0 U99 ( .INP(N12), .ZN(n90) );
  INVX0 U100 ( .INP(N11), .ZN(n91) );
endmodule


module add_545 ( s, a, b, co, ci_BAR );
  input a, b, ci_BAR;
  output s, co;


  XOR2X1 U1 ( .IN1(a), .IN2(ci_BAR), .Q(s) );
endmodule


module add_546 ( s, a, b, ci, co_BAR );
  input a, b, ci;
  output s, co_BAR;


  NAND2X0 U1 ( .IN1(ci), .IN2(a), .QN(co_BAR) );
  OA21X1 U2 ( .IN1(ci), .IN2(a), .IN3(co_BAR), .Q(s) );
endmodule


module add_547 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_548 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_549 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_550 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_551 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  INVX0 U1 ( .INP(a), .ZN(s) );
  NBUFFX2 U2 ( .INP(a), .Z(co) );
endmodule


module add_552 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  NBUFFX2 U1 ( .INP(a), .Z(s) );
endmodule


module adder8_39 ( out, a, b, cin );
  output [7:0] out;
  input [7:0] a;
  input [7:0] b;
  input cin;

  wire   [6:1] c;

  add_552 add_01 ( .s(out[0]), .a(a[0]), .b(1'b1), .ci(1'b1) );
  add_551 add_02 ( .s(out[1]), .a(a[1]), .b(1'b0), .ci(1'b1), .co(c[1]) );
  add_550 add_03 ( .s(out[2]), .a(a[2]), .b(1'b0), .ci(c[1]), .co(c[2]) );
  add_549 add_04 ( .s(out[3]), .a(a[3]), .b(1'b0), .ci(c[2]), .co(c[3]) );
  add_548 add_05 ( .s(out[4]), .a(a[4]), .b(1'b0), .ci(c[3]), .co(c[4]) );
  add_547 add_06 ( .s(out[5]), .a(a[5]), .b(1'b0), .ci(c[4]), .co(c[5]) );
  add_546 add_07 ( .s(out[6]), .a(a[6]), .b(1'b0), .ci(c[5]), .co_BAR(c[6]) );
  add_545 add_08 ( .s(out[7]), .a(a[7]), .b(1'b1), .ci_BAR(c[6]) );
endmodule


module add_553 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  XOR3X1 U1 ( .IN1(b), .IN2(ci), .IN3(a), .Q(s) );
endmodule


module add_554 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_555 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_556 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_557 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_558 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_559 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_560 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(b), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(b), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module adder8_40 ( out, a, b, cin );
  output [7:0] out;
  input [7:0] a;
  input [7:0] b;
  input cin;

  wire   [6:0] c;

  add_560 add_01 ( .s(out[0]), .a(a[0]), .b(b[0]), .ci(1'b0), .co(c[0]) );
  add_559 add_02 ( .s(out[1]), .a(a[1]), .b(b[1]), .ci(c[0]), .co(c[1]) );
  add_558 add_03 ( .s(out[2]), .a(a[2]), .b(b[2]), .ci(c[1]), .co(c[2]) );
  add_557 add_04 ( .s(out[3]), .a(a[3]), .b(b[3]), .ci(c[2]), .co(c[3]) );
  add_556 add_05 ( .s(out[4]), .a(a[4]), .b(b[4]), .ci(c[3]), .co(c[4]) );
  add_555 add_06 ( .s(out[5]), .a(a[5]), .b(b[5]), .ci(c[4]), .co(c[5]) );
  add_554 add_07 ( .s(out[6]), .a(a[6]), .b(b[6]), .ci(c[5]), .co(c[6]) );
  add_553 add_08 ( .s(out[7]), .a(a[7]), .b(b[7]), .ci(c[6]) );
endmodule


module floating_point_multiple_5 ( clk, rst_n, input_factor_01, 
        input_factor_02, output_multiply );
  input [31:0] input_factor_01;
  input [31:0] input_factor_02;
  output [31:0] output_multiply;
  input clk, rst_n;
  wire   N5, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22,
         N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N48, N49, N50, N51,
         N52, N53, N54, N55, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22,
         SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24,
         SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26;
  wire   [47:23] base_multiply_result;
  wire   [47:23] mulout;
  wire   [7:0] exponent_factor_12;
  wire   [7:0] pre_mul_output_exponent;

  mul26_5 mul26_01 ( .clk(clk), .rst_n(rst_n), .in1({1'b0, 1'b0, 1'b1, 
        input_factor_01[22:0]}), .in2({1'b0, 1'b0, 1'b1, input_factor_02[22:0]}), .en(1'b1), .mulout({SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, 
        SYNOPSYS_UNCONNECTED_3, mulout, SYNOPSYS_UNCONNECTED_4, 
        SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, 
        SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, 
        SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11, 
        SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13, 
        SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, 
        SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17, 
        SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19, 
        SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21, 
        SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_23, 
        SYNOPSYS_UNCONNECTED_24, SYNOPSYS_UNCONNECTED_25, 
        SYNOPSYS_UNCONNECTED_26}) );
  adder8_40 adder8_01 ( .out(exponent_factor_12), .a(input_factor_01[30:23]), 
        .b(input_factor_02[30:23]), .cin(1'b0) );
  adder8_39 adder8_02 ( .out(pre_mul_output_exponent), .a(exponent_factor_12), 
        .b({1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0}), .cin(1'b1) );
  DFFARX1 mul_output_sign_reg ( .D(N5), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[31]) );
  DFFARX1 base_multiply_result_reg_47_ ( .D(mulout[47]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[47]) );
  DFFARX1 base_multiply_result_reg_46_ ( .D(mulout[46]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[46]) );
  DFFARX1 base_multiply_result_reg_45_ ( .D(mulout[45]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[45]) );
  DFFARX1 base_multiply_result_reg_44_ ( .D(mulout[44]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[44]) );
  DFFARX1 base_multiply_result_reg_43_ ( .D(mulout[43]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[43]) );
  DFFARX1 base_multiply_result_reg_42_ ( .D(mulout[42]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[42]) );
  DFFARX1 base_multiply_result_reg_41_ ( .D(mulout[41]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[41]) );
  DFFARX1 base_multiply_result_reg_40_ ( .D(mulout[40]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[40]) );
  DFFARX1 base_multiply_result_reg_39_ ( .D(mulout[39]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[39]) );
  DFFARX1 base_multiply_result_reg_38_ ( .D(mulout[38]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[38]) );
  DFFARX1 base_multiply_result_reg_37_ ( .D(mulout[37]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[37]) );
  DFFARX1 base_multiply_result_reg_36_ ( .D(mulout[36]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[36]) );
  DFFARX1 base_multiply_result_reg_35_ ( .D(mulout[35]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[35]) );
  DFFARX1 base_multiply_result_reg_34_ ( .D(mulout[34]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[34]) );
  DFFARX1 base_multiply_result_reg_33_ ( .D(mulout[33]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[33]) );
  DFFARX1 base_multiply_result_reg_32_ ( .D(mulout[32]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[32]) );
  DFFARX1 base_multiply_result_reg_31_ ( .D(mulout[31]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[31]) );
  DFFARX1 base_multiply_result_reg_30_ ( .D(mulout[30]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[30]) );
  DFFARX1 base_multiply_result_reg_29_ ( .D(mulout[29]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[29]) );
  DFFARX1 base_multiply_result_reg_28_ ( .D(mulout[28]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[28]) );
  DFFARX1 base_multiply_result_reg_27_ ( .D(mulout[27]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[27]) );
  DFFARX1 base_multiply_result_reg_26_ ( .D(mulout[26]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[26]) );
  DFFARX1 base_multiply_result_reg_25_ ( .D(mulout[25]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[25]) );
  DFFARX1 base_multiply_result_reg_24_ ( .D(mulout[24]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[24]) );
  DFFARX1 base_multiply_result_reg_23_ ( .D(mulout[23]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[23]) );
  DFFARX1 mul_output_significand_reg_22_ ( .D(N32), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[22]) );
  DFFARX1 mul_output_significand_reg_21_ ( .D(N31), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[21]) );
  DFFARX1 mul_output_significand_reg_20_ ( .D(N30), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[20]) );
  DFFARX1 mul_output_significand_reg_19_ ( .D(N29), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[19]) );
  DFFARX1 mul_output_significand_reg_18_ ( .D(N28), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[18]) );
  DFFARX1 mul_output_significand_reg_17_ ( .D(N27), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[17]) );
  DFFARX1 mul_output_significand_reg_16_ ( .D(N26), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[16]) );
  DFFARX1 mul_output_significand_reg_15_ ( .D(N25), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[15]) );
  DFFARX1 mul_output_significand_reg_14_ ( .D(N24), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[14]) );
  DFFARX1 mul_output_significand_reg_13_ ( .D(N23), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[13]) );
  DFFARX1 mul_output_significand_reg_12_ ( .D(N22), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[12]) );
  DFFARX1 mul_output_significand_reg_11_ ( .D(N21), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[11]) );
  DFFARX1 mul_output_significand_reg_10_ ( .D(N20), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[10]) );
  DFFARX1 mul_output_significand_reg_9_ ( .D(N19), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[9]) );
  DFFARX1 mul_output_significand_reg_8_ ( .D(N18), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[8]) );
  DFFARX1 mul_output_significand_reg_7_ ( .D(N17), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[7]) );
  DFFARX1 mul_output_significand_reg_6_ ( .D(N16), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[6]) );
  DFFARX1 mul_output_significand_reg_5_ ( .D(N15), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[5]) );
  DFFARX1 mul_output_significand_reg_4_ ( .D(N14), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[4]) );
  DFFARX1 mul_output_significand_reg_3_ ( .D(N13), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[3]) );
  DFFARX1 mul_output_significand_reg_2_ ( .D(N12), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[2]) );
  DFFARX1 mul_output_significand_reg_1_ ( .D(N11), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[1]) );
  DFFARX1 mul_output_significand_reg_0_ ( .D(N10), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[0]) );
  DFFARX1 mul_output_exponent_reg_7_ ( .D(N55), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[30]) );
  DFFARX1 mul_output_exponent_reg_6_ ( .D(N54), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[29]) );
  DFFARX1 mul_output_exponent_reg_5_ ( .D(N53), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[28]) );
  DFFARX1 mul_output_exponent_reg_4_ ( .D(N52), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[27]) );
  DFFARX1 mul_output_exponent_reg_3_ ( .D(N51), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[26]) );
  DFFARX1 mul_output_exponent_reg_2_ ( .D(N50), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[25]) );
  DFFARX1 mul_output_exponent_reg_1_ ( .D(N49), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[24]) );
  DFFARX1 mul_output_exponent_reg_0_ ( .D(N48), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[23]) );
  AND2X1 U3 ( .IN1(base_multiply_result[47]), .IN2(n35), .Q(n32) );
  INVX0 U4 ( .INP(n1), .ZN(n2) );
  OR2X1 U5 ( .IN1(base_multiply_result[47]), .IN2(n24), .Q(n1) );
  INVX0 U6 ( .INP(input_factor_02[31]), .ZN(n3) );
  NOR4X0 U7 ( .IN1(input_factor_01[0]), .IN2(input_factor_01[10]), .IN3(
        input_factor_01[11]), .IN4(input_factor_01[12]), .QN(n7) );
  NOR4X0 U8 ( .IN1(input_factor_01[13]), .IN2(input_factor_01[14]), .IN3(
        input_factor_01[15]), .IN4(input_factor_01[16]), .QN(n6) );
  NOR4X0 U9 ( .IN1(input_factor_01[17]), .IN2(input_factor_01[18]), .IN3(
        input_factor_01[19]), .IN4(input_factor_01[1]), .QN(n5) );
  NOR4X0 U10 ( .IN1(input_factor_01[20]), .IN2(input_factor_01[21]), .IN3(
        input_factor_01[22]), .IN4(input_factor_01[23]), .QN(n4) );
  NAND4X0 U11 ( .IN1(n7), .IN2(n6), .IN3(n5), .IN4(n4), .QN(n23) );
  NOR4X0 U12 ( .IN1(input_factor_01[24]), .IN2(input_factor_01[25]), .IN3(
        input_factor_01[26]), .IN4(input_factor_01[27]), .QN(n11) );
  NOR4X0 U13 ( .IN1(input_factor_01[28]), .IN2(input_factor_01[29]), .IN3(
        input_factor_01[2]), .IN4(input_factor_01[30]), .QN(n10) );
  NOR4X0 U14 ( .IN1(input_factor_01[31]), .IN2(input_factor_01[3]), .IN3(
        input_factor_01[4]), .IN4(input_factor_01[5]), .QN(n9) );
  NOR4X0 U15 ( .IN1(input_factor_01[6]), .IN2(input_factor_01[7]), .IN3(
        input_factor_01[8]), .IN4(input_factor_01[9]), .QN(n8) );
  NAND4X0 U16 ( .IN1(n11), .IN2(n10), .IN3(n9), .IN4(n8), .QN(n22) );
  NOR4X0 U17 ( .IN1(input_factor_02[0]), .IN2(input_factor_02[10]), .IN3(
        input_factor_02[11]), .IN4(input_factor_02[12]), .QN(n15) );
  NOR4X0 U18 ( .IN1(input_factor_02[13]), .IN2(input_factor_02[14]), .IN3(
        input_factor_02[15]), .IN4(input_factor_02[16]), .QN(n14) );
  NOR4X0 U19 ( .IN1(input_factor_02[17]), .IN2(input_factor_02[18]), .IN3(
        input_factor_02[19]), .IN4(input_factor_02[1]), .QN(n13) );
  NOR4X0 U20 ( .IN1(input_factor_02[20]), .IN2(input_factor_02[21]), .IN3(
        input_factor_02[22]), .IN4(input_factor_02[23]), .QN(n12) );
  NAND4X0 U21 ( .IN1(n15), .IN2(n14), .IN3(n13), .IN4(n12), .QN(n21) );
  NOR4X0 U22 ( .IN1(input_factor_02[24]), .IN2(input_factor_02[25]), .IN3(
        input_factor_02[26]), .IN4(input_factor_02[27]), .QN(n19) );
  NOR4X0 U23 ( .IN1(input_factor_02[28]), .IN2(input_factor_02[29]), .IN3(
        input_factor_02[2]), .IN4(input_factor_02[30]), .QN(n18) );
  NOR4X0 U24 ( .IN1(input_factor_02[31]), .IN2(input_factor_02[3]), .IN3(
        input_factor_02[4]), .IN4(input_factor_02[5]), .QN(n17) );
  NOR4X0 U25 ( .IN1(input_factor_02[6]), .IN2(input_factor_02[7]), .IN3(
        input_factor_02[8]), .IN4(input_factor_02[9]), .QN(n16) );
  NAND4X0 U26 ( .IN1(n19), .IN2(n18), .IN3(n17), .IN4(n16), .QN(n20) );
  OA22X1 U27 ( .IN1(n23), .IN2(n22), .IN3(n21), .IN4(n20), .Q(n35) );
  INVX0 U28 ( .INP(n35), .ZN(n24) );
  AO22X1 U29 ( .IN1(n2), .IN2(base_multiply_result[23]), .IN3(n32), .IN4(
        base_multiply_result[24]), .Q(N10) );
  AO22X1 U30 ( .IN1(n2), .IN2(base_multiply_result[24]), .IN3(n32), .IN4(
        base_multiply_result[25]), .Q(N11) );
  AO22X1 U31 ( .IN1(n2), .IN2(base_multiply_result[25]), .IN3(n32), .IN4(
        base_multiply_result[26]), .Q(N12) );
  AO22X1 U32 ( .IN1(n2), .IN2(base_multiply_result[26]), .IN3(n32), .IN4(
        base_multiply_result[27]), .Q(N13) );
  AO22X1 U33 ( .IN1(n2), .IN2(base_multiply_result[27]), .IN3(n32), .IN4(
        base_multiply_result[28]), .Q(N14) );
  AO22X1 U34 ( .IN1(n2), .IN2(base_multiply_result[28]), .IN3(n32), .IN4(
        base_multiply_result[29]), .Q(N15) );
  AO22X1 U35 ( .IN1(n2), .IN2(base_multiply_result[29]), .IN3(n32), .IN4(
        base_multiply_result[30]), .Q(N16) );
  AO22X1 U36 ( .IN1(n2), .IN2(base_multiply_result[30]), .IN3(n32), .IN4(
        base_multiply_result[31]), .Q(N17) );
  AO22X1 U37 ( .IN1(n2), .IN2(base_multiply_result[31]), .IN3(n32), .IN4(
        base_multiply_result[32]), .Q(N18) );
  AO22X1 U38 ( .IN1(n2), .IN2(base_multiply_result[32]), .IN3(n32), .IN4(
        base_multiply_result[33]), .Q(N19) );
  AO22X1 U39 ( .IN1(n2), .IN2(base_multiply_result[33]), .IN3(n32), .IN4(
        base_multiply_result[34]), .Q(N20) );
  AO22X1 U40 ( .IN1(n2), .IN2(base_multiply_result[34]), .IN3(n32), .IN4(
        base_multiply_result[35]), .Q(N21) );
  AO22X1 U41 ( .IN1(n2), .IN2(base_multiply_result[35]), .IN3(n32), .IN4(
        base_multiply_result[36]), .Q(N22) );
  AO22X1 U42 ( .IN1(n2), .IN2(base_multiply_result[36]), .IN3(n32), .IN4(
        base_multiply_result[37]), .Q(N23) );
  AO22X1 U43 ( .IN1(n2), .IN2(base_multiply_result[37]), .IN3(n32), .IN4(
        base_multiply_result[38]), .Q(N24) );
  AO22X1 U44 ( .IN1(n2), .IN2(base_multiply_result[38]), .IN3(n32), .IN4(
        base_multiply_result[39]), .Q(N25) );
  AO22X1 U45 ( .IN1(n2), .IN2(base_multiply_result[39]), .IN3(n32), .IN4(
        base_multiply_result[40]), .Q(N26) );
  AO22X1 U46 ( .IN1(n2), .IN2(base_multiply_result[40]), .IN3(n32), .IN4(
        base_multiply_result[41]), .Q(N27) );
  AO22X1 U47 ( .IN1(n2), .IN2(base_multiply_result[41]), .IN3(n32), .IN4(
        base_multiply_result[42]), .Q(N28) );
  AO22X1 U48 ( .IN1(n2), .IN2(base_multiply_result[42]), .IN3(n32), .IN4(
        base_multiply_result[43]), .Q(N29) );
  AO22X1 U49 ( .IN1(n2), .IN2(base_multiply_result[43]), .IN3(n32), .IN4(
        base_multiply_result[44]), .Q(N30) );
  AO22X1 U50 ( .IN1(n2), .IN2(base_multiply_result[44]), .IN3(n32), .IN4(
        base_multiply_result[45]), .Q(N31) );
  AO22X1 U51 ( .IN1(n2), .IN2(base_multiply_result[45]), .IN3(n32), .IN4(
        base_multiply_result[46]), .Q(N32) );
  MUX21X1 U52 ( .IN1(n2), .IN2(n32), .S(pre_mul_output_exponent[0]), .Q(N48)
         );
  AO21X1 U53 ( .IN1(pre_mul_output_exponent[0]), .IN2(n2), .IN3(n32), .Q(n25)
         );
  NOR3X0 U54 ( .IN1(pre_mul_output_exponent[1]), .IN2(
        pre_mul_output_exponent[0]), .IN3(n1), .QN(n27) );
  AO21X1 U55 ( .IN1(pre_mul_output_exponent[1]), .IN2(n25), .IN3(n27), .Q(N49)
         );
  INVX0 U56 ( .INP(input_factor_01[31]), .ZN(n26) );
  OA221X1 U57 ( .IN1(input_factor_01[31]), .IN2(input_factor_02[31]), .IN3(n26), .IN4(n3), .IN5(n35), .Q(N5) );
  AO221X1 U58 ( .IN1(n2), .IN2(pre_mul_output_exponent[1]), .IN3(n2), .IN4(
        pre_mul_output_exponent[0]), .IN5(n32), .Q(n28) );
  MUX21X1 U59 ( .IN1(n27), .IN2(n28), .S(pre_mul_output_exponent[2]), .Q(N50)
         );
  AND2X1 U60 ( .IN1(n2), .IN2(pre_mul_output_exponent[2]), .Q(n29) );
  OR4X1 U61 ( .IN1(pre_mul_output_exponent[1]), .IN2(
        pre_mul_output_exponent[0]), .IN3(pre_mul_output_exponent[3]), .IN4(
        pre_mul_output_exponent[2]), .Q(n34) );
  NOR2X0 U62 ( .IN1(n1), .IN2(n34), .QN(n31) );
  AO221X1 U63 ( .IN1(pre_mul_output_exponent[3]), .IN2(n29), .IN3(
        pre_mul_output_exponent[3]), .IN4(n28), .IN5(n31), .Q(N51) );
  OA21X1 U64 ( .IN1(base_multiply_result[47]), .IN2(n34), .IN3(n35), .Q(n30)
         );
  MUX21X1 U65 ( .IN1(n31), .IN2(n30), .S(pre_mul_output_exponent[4]), .Q(N52)
         );
  AO221X1 U66 ( .IN1(n2), .IN2(pre_mul_output_exponent[4]), .IN3(n2), .IN4(n34), .IN5(n32), .Q(n33) );
  NOR4X0 U67 ( .IN1(pre_mul_output_exponent[5]), .IN2(
        pre_mul_output_exponent[4]), .IN3(n34), .IN4(n1), .QN(n37) );
  AO21X1 U68 ( .IN1(pre_mul_output_exponent[5]), .IN2(n33), .IN3(n37), .Q(N53)
         );
  OR3X1 U69 ( .IN1(pre_mul_output_exponent[5]), .IN2(
        pre_mul_output_exponent[4]), .IN3(n34), .Q(n36) );
  OA21X1 U70 ( .IN1(base_multiply_result[47]), .IN2(n36), .IN3(n35), .Q(n39)
         );
  INVX0 U71 ( .INP(n37), .ZN(n38) );
  NOR2X0 U72 ( .IN1(pre_mul_output_exponent[6]), .IN2(n38), .QN(n41) );
  AO21X1 U73 ( .IN1(pre_mul_output_exponent[6]), .IN2(n39), .IN3(n41), .Q(N54)
         );
  AO21X1 U74 ( .IN1(n2), .IN2(pre_mul_output_exponent[6]), .IN3(n39), .Q(n40)
         );
  MUX21X1 U75 ( .IN1(n41), .IN2(n40), .S(pre_mul_output_exponent[7]), .Q(N55)
         );
endmodule


module cla51squ_6 ( out, a, b );
  output [50:0] out;
  input [50:0] a;
  input [50:0] b;
  wire   intadd_6_CI, intadd_6_n24, intadd_6_n23, intadd_6_n22, intadd_6_n21,
         intadd_6_n20, intadd_6_n19, intadd_6_n18, intadd_6_n17, intadd_6_n16,
         intadd_6_n15, intadd_6_n14, intadd_6_n13, intadd_6_n12, intadd_6_n11,
         intadd_6_n10, intadd_6_n9, intadd_6_n8, intadd_6_n7, intadd_6_n6,
         intadd_6_n5, intadd_6_n4, intadd_6_n3, intadd_6_n2, intadd_6_n1, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14;

  FADDX1 intadd_6_U25 ( .A(b[23]), .B(a[23]), .CI(intadd_6_CI), .CO(
        intadd_6_n24), .S(out[23]) );
  FADDX1 intadd_6_U24 ( .A(b[24]), .B(a[24]), .CI(intadd_6_n24), .CO(
        intadd_6_n23), .S(out[24]) );
  FADDX1 intadd_6_U23 ( .A(b[25]), .B(a[25]), .CI(intadd_6_n23), .CO(
        intadd_6_n22), .S(out[25]) );
  FADDX1 intadd_6_U22 ( .A(b[26]), .B(a[26]), .CI(intadd_6_n22), .CO(
        intadd_6_n21), .S(out[26]) );
  FADDX1 intadd_6_U21 ( .A(b[27]), .B(a[27]), .CI(intadd_6_n21), .CO(
        intadd_6_n20), .S(out[27]) );
  FADDX1 intadd_6_U20 ( .A(b[28]), .B(a[28]), .CI(intadd_6_n20), .CO(
        intadd_6_n19), .S(out[28]) );
  FADDX1 intadd_6_U19 ( .A(b[29]), .B(a[29]), .CI(intadd_6_n19), .CO(
        intadd_6_n18), .S(out[29]) );
  FADDX1 intadd_6_U18 ( .A(b[30]), .B(a[30]), .CI(intadd_6_n18), .CO(
        intadd_6_n17), .S(out[30]) );
  FADDX1 intadd_6_U17 ( .A(b[31]), .B(a[31]), .CI(intadd_6_n17), .CO(
        intadd_6_n16), .S(out[31]) );
  FADDX1 intadd_6_U16 ( .A(b[32]), .B(a[32]), .CI(intadd_6_n16), .CO(
        intadd_6_n15), .S(out[32]) );
  FADDX1 intadd_6_U15 ( .A(b[33]), .B(a[33]), .CI(intadd_6_n15), .CO(
        intadd_6_n14), .S(out[33]) );
  FADDX1 intadd_6_U14 ( .A(b[34]), .B(a[34]), .CI(intadd_6_n14), .CO(
        intadd_6_n13), .S(out[34]) );
  FADDX1 intadd_6_U13 ( .A(b[35]), .B(a[35]), .CI(intadd_6_n13), .CO(
        intadd_6_n12), .S(out[35]) );
  FADDX1 intadd_6_U12 ( .A(b[36]), .B(a[36]), .CI(intadd_6_n12), .CO(
        intadd_6_n11), .S(out[36]) );
  FADDX1 intadd_6_U11 ( .A(b[37]), .B(a[37]), .CI(intadd_6_n11), .CO(
        intadd_6_n10), .S(out[37]) );
  FADDX1 intadd_6_U10 ( .A(b[38]), .B(a[38]), .CI(intadd_6_n10), .CO(
        intadd_6_n9), .S(out[38]) );
  FADDX1 intadd_6_U9 ( .A(b[39]), .B(a[39]), .CI(intadd_6_n9), .CO(intadd_6_n8), .S(out[39]) );
  FADDX1 intadd_6_U8 ( .A(b[40]), .B(a[40]), .CI(intadd_6_n8), .CO(intadd_6_n7), .S(out[40]) );
  FADDX1 intadd_6_U7 ( .A(b[41]), .B(a[41]), .CI(intadd_6_n7), .CO(intadd_6_n6), .S(out[41]) );
  FADDX1 intadd_6_U6 ( .A(b[42]), .B(a[42]), .CI(intadd_6_n6), .CO(intadd_6_n5), .S(out[42]) );
  FADDX1 intadd_6_U5 ( .A(b[43]), .B(a[43]), .CI(intadd_6_n5), .CO(intadd_6_n4), .S(out[43]) );
  FADDX1 intadd_6_U4 ( .A(b[44]), .B(a[44]), .CI(intadd_6_n4), .CO(intadd_6_n3), .S(out[44]) );
  FADDX1 intadd_6_U3 ( .A(b[45]), .B(a[45]), .CI(intadd_6_n3), .CO(intadd_6_n2), .S(out[45]) );
  FADDX1 intadd_6_U2 ( .A(b[46]), .B(a[46]), .CI(intadd_6_n2), .CO(intadd_6_n1), .S(out[46]) );
  OA21X1 U2 ( .IN1(b[9]), .IN2(a[9]), .IN3(a[8]), .Q(n1) );
  AO22X1 U3 ( .IN1(b[9]), .IN2(a[9]), .IN3(b[8]), .IN4(n1), .Q(n2) );
  AO222X1 U4 ( .IN1(b[10]), .IN2(a[10]), .IN3(b[10]), .IN4(n2), .IN5(a[10]), 
        .IN6(n2), .Q(n3) );
  AO222X1 U5 ( .IN1(b[11]), .IN2(a[11]), .IN3(b[11]), .IN4(n3), .IN5(a[11]), 
        .IN6(n3), .Q(n4) );
  AO222X1 U6 ( .IN1(b[12]), .IN2(a[12]), .IN3(b[12]), .IN4(n4), .IN5(a[12]), 
        .IN6(n4), .Q(n5) );
  AO222X1 U7 ( .IN1(b[13]), .IN2(a[13]), .IN3(b[13]), .IN4(n5), .IN5(a[13]), 
        .IN6(n5), .Q(n6) );
  AO222X1 U8 ( .IN1(b[14]), .IN2(a[14]), .IN3(b[14]), .IN4(n6), .IN5(a[14]), 
        .IN6(n6), .Q(n7) );
  AO222X1 U9 ( .IN1(b[15]), .IN2(a[15]), .IN3(b[15]), .IN4(n7), .IN5(a[15]), 
        .IN6(n7), .Q(n8) );
  AO222X1 U10 ( .IN1(b[16]), .IN2(a[16]), .IN3(b[16]), .IN4(n8), .IN5(a[16]), 
        .IN6(n8), .Q(n9) );
  AO222X1 U11 ( .IN1(b[17]), .IN2(a[17]), .IN3(b[17]), .IN4(n9), .IN5(a[17]), 
        .IN6(n9), .Q(n10) );
  AO222X1 U12 ( .IN1(b[18]), .IN2(a[18]), .IN3(b[18]), .IN4(n10), .IN5(a[18]), 
        .IN6(n10), .Q(n11) );
  AO222X1 U13 ( .IN1(b[19]), .IN2(a[19]), .IN3(b[19]), .IN4(n11), .IN5(a[19]), 
        .IN6(n11), .Q(n12) );
  AO222X1 U14 ( .IN1(b[20]), .IN2(a[20]), .IN3(b[20]), .IN4(n12), .IN5(a[20]), 
        .IN6(n12), .Q(n13) );
  AO222X1 U15 ( .IN1(b[21]), .IN2(a[21]), .IN3(b[21]), .IN4(n13), .IN5(a[21]), 
        .IN6(n13), .Q(n14) );
  AO222X1 U16 ( .IN1(b[22]), .IN2(a[22]), .IN3(b[22]), .IN4(n14), .IN5(a[22]), 
        .IN6(n14), .Q(intadd_6_CI) );
  XOR3X1 U17 ( .IN1(intadd_6_n1), .IN2(a[47]), .IN3(b[47]), .Q(out[47]) );
endmodule


module csa51squ_61 ( sumout, in1, in2, in3, cout_50_, cout_49_, cout_48_, 
        cout_47_, cout_46_, cout_44_, cout_42_, cout_40_, cout_38_, cout_36_, 
        cout_34_, cout_32_, cout_30_, cout_28_, cout_27_, cout_7__BAR, cout_6_, 
        cout_5_, cout_4_, cout_3_, cout_2_, cout_1_, cout_0_, cout_8__BAR, 
        cout_9__BAR, cout_10__BAR, cout_11__BAR, cout_12__BAR, cout_13__BAR, 
        cout_14__BAR, cout_15__BAR, cout_16__BAR, cout_17__BAR, cout_18__BAR, 
        cout_19__BAR, cout_20__BAR, cout_21__BAR, cout_22__BAR, cout_23__BAR, 
        cout_24__BAR, cout_25__BAR, cout_26__BAR, cout_29__BAR, cout_31__BAR, 
        cout_33__BAR, cout_35__BAR, cout_37__BAR, cout_39__BAR, cout_41__BAR, 
        cout_43__BAR, cout_45__BAR );
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  output cout_50_, cout_49_, cout_48_, cout_47_, cout_46_, cout_44_, cout_42_,
         cout_40_, cout_38_, cout_36_, cout_34_, cout_32_, cout_30_, cout_28_,
         cout_27_, cout_7__BAR, cout_6_, cout_5_, cout_4_, cout_3_, cout_2_,
         cout_1_, cout_0_, cout_8__BAR, cout_9__BAR, cout_10__BAR,
         cout_11__BAR, cout_12__BAR, cout_13__BAR, cout_14__BAR, cout_15__BAR,
         cout_16__BAR, cout_17__BAR, cout_18__BAR, cout_19__BAR, cout_20__BAR,
         cout_21__BAR, cout_22__BAR, cout_23__BAR, cout_24__BAR, cout_25__BAR,
         cout_26__BAR, cout_29__BAR, cout_31__BAR, cout_33__BAR, cout_35__BAR,
         cout_37__BAR, cout_39__BAR, cout_41__BAR, cout_43__BAR, cout_45__BAR;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11;

  NAND2X0 U1 ( .IN1(in2[8]), .IN2(in1[8]), .QN(cout_8__BAR) );
  NAND2X0 U2 ( .IN1(in2[9]), .IN2(in1[9]), .QN(cout_9__BAR) );
  NAND2X0 U3 ( .IN1(in2[10]), .IN2(in1[10]), .QN(cout_10__BAR) );
  NAND2X0 U4 ( .IN1(in2[11]), .IN2(in1[11]), .QN(cout_11__BAR) );
  NAND2X0 U5 ( .IN1(in2[12]), .IN2(in1[12]), .QN(cout_12__BAR) );
  NAND2X0 U6 ( .IN1(in2[13]), .IN2(in1[13]), .QN(cout_13__BAR) );
  NAND2X0 U7 ( .IN1(in2[14]), .IN2(in1[14]), .QN(cout_14__BAR) );
  NAND2X0 U8 ( .IN1(in2[15]), .IN2(in1[15]), .QN(cout_15__BAR) );
  NAND2X0 U9 ( .IN1(in2[16]), .IN2(in1[16]), .QN(cout_16__BAR) );
  NAND2X0 U10 ( .IN1(in2[17]), .IN2(in1[17]), .QN(cout_17__BAR) );
  NAND2X0 U11 ( .IN1(in2[18]), .IN2(in1[18]), .QN(cout_18__BAR) );
  NAND2X0 U12 ( .IN1(in2[19]), .IN2(in1[19]), .QN(cout_19__BAR) );
  NAND2X0 U13 ( .IN1(in2[20]), .IN2(in1[20]), .QN(cout_20__BAR) );
  NAND2X0 U14 ( .IN1(in2[21]), .IN2(in1[21]), .QN(cout_21__BAR) );
  NAND2X0 U15 ( .IN1(in2[22]), .IN2(in1[22]), .QN(cout_22__BAR) );
  NAND2X0 U16 ( .IN1(in2[23]), .IN2(in1[23]), .QN(cout_23__BAR) );
  NAND2X0 U17 ( .IN1(in2[24]), .IN2(in1[24]), .QN(cout_24__BAR) );
  NAND2X0 U18 ( .IN1(in2[25]), .IN2(in1[25]), .QN(cout_25__BAR) );
  NAND2X0 U19 ( .IN1(in2[26]), .IN2(in1[26]), .QN(cout_26__BAR) );
  NAND2X0 U20 ( .IN1(in2[29]), .IN2(in1[29]), .QN(cout_29__BAR) );
  NAND2X0 U21 ( .IN1(in2[31]), .IN2(in1[31]), .QN(cout_31__BAR) );
  NAND2X0 U22 ( .IN1(in2[33]), .IN2(in1[33]), .QN(cout_33__BAR) );
  NAND2X0 U23 ( .IN1(in2[35]), .IN2(in1[35]), .QN(cout_35__BAR) );
  NAND2X0 U24 ( .IN1(in2[37]), .IN2(in1[37]), .QN(cout_37__BAR) );
  NAND2X0 U25 ( .IN1(in2[39]), .IN2(in1[39]), .QN(cout_39__BAR) );
  NAND2X0 U26 ( .IN1(in2[41]), .IN2(in1[41]), .QN(cout_41__BAR) );
  NAND2X0 U27 ( .IN1(in2[43]), .IN2(in1[43]), .QN(cout_43__BAR) );
  NAND2X0 U28 ( .IN1(in2[45]), .IN2(in1[45]), .QN(cout_45__BAR) );
  NAND2X0 U29 ( .IN1(in2[7]), .IN2(in1[7]), .QN(cout_7__BAR) );
  NAND2X0 U30 ( .IN1(n1), .IN2(cout_27_), .QN(sumout[27]) );
  NAND2X0 U31 ( .IN1(in1[27]), .IN2(in2[27]), .QN(n1) );
  NAND2X0 U32 ( .IN1(n2), .IN2(cout_28_), .QN(sumout[28]) );
  NAND2X0 U33 ( .IN1(in1[28]), .IN2(in2[28]), .QN(n2) );
  NAND2X0 U34 ( .IN1(n3), .IN2(cout_30_), .QN(sumout[30]) );
  NAND2X0 U35 ( .IN1(in1[30]), .IN2(in2[30]), .QN(n3) );
  NAND2X0 U36 ( .IN1(n4), .IN2(cout_32_), .QN(sumout[32]) );
  NAND2X0 U37 ( .IN1(in1[32]), .IN2(in2[32]), .QN(n4) );
  NAND2X0 U38 ( .IN1(n5), .IN2(cout_34_), .QN(sumout[34]) );
  NAND2X0 U39 ( .IN1(in1[34]), .IN2(in2[34]), .QN(n5) );
  NAND2X0 U40 ( .IN1(n6), .IN2(cout_36_), .QN(sumout[36]) );
  NAND2X0 U41 ( .IN1(in1[36]), .IN2(in2[36]), .QN(n6) );
  NAND2X0 U42 ( .IN1(n7), .IN2(cout_38_), .QN(sumout[38]) );
  NAND2X0 U43 ( .IN1(in1[38]), .IN2(in2[38]), .QN(n7) );
  NAND2X0 U44 ( .IN1(n8), .IN2(cout_40_), .QN(sumout[40]) );
  NAND2X0 U45 ( .IN1(in1[40]), .IN2(in2[40]), .QN(n8) );
  NAND2X0 U46 ( .IN1(n9), .IN2(cout_42_), .QN(sumout[42]) );
  NAND2X0 U47 ( .IN1(in1[42]), .IN2(in2[42]), .QN(n9) );
  NAND2X0 U48 ( .IN1(n10), .IN2(cout_44_), .QN(sumout[44]) );
  NAND2X0 U49 ( .IN1(in1[44]), .IN2(in2[44]), .QN(n10) );
  NAND2X0 U50 ( .IN1(n11), .IN2(cout_46_), .QN(sumout[46]) );
  NAND2X0 U51 ( .IN1(in1[46]), .IN2(in2[46]), .QN(n11) );
  OR2X1 U52 ( .IN1(in2[27]), .IN2(in1[27]), .Q(cout_27_) );
  OR2X1 U53 ( .IN1(in2[28]), .IN2(in1[28]), .Q(cout_28_) );
  OR2X1 U54 ( .IN1(in2[30]), .IN2(in1[30]), .Q(cout_30_) );
  OR2X1 U55 ( .IN1(in2[32]), .IN2(in1[32]), .Q(cout_32_) );
  OR2X1 U56 ( .IN1(in2[34]), .IN2(in1[34]), .Q(cout_34_) );
  OR2X1 U57 ( .IN1(in2[36]), .IN2(in1[36]), .Q(cout_36_) );
  OR2X1 U58 ( .IN1(in2[38]), .IN2(in1[38]), .Q(cout_38_) );
  OR2X1 U59 ( .IN1(in2[40]), .IN2(in1[40]), .Q(cout_40_) );
  OR2X1 U60 ( .IN1(in2[42]), .IN2(in1[42]), .Q(cout_42_) );
  OR2X1 U61 ( .IN1(in2[44]), .IN2(in1[44]), .Q(cout_44_) );
  OR2X1 U62 ( .IN1(in2[46]), .IN2(in1[46]), .Q(cout_46_) );
  OA21X1 U63 ( .IN1(in2[8]), .IN2(in1[8]), .IN3(cout_8__BAR), .Q(sumout[8]) );
  OA21X1 U64 ( .IN1(in2[9]), .IN2(in1[9]), .IN3(cout_9__BAR), .Q(sumout[9]) );
  OA21X1 U65 ( .IN1(in2[10]), .IN2(in1[10]), .IN3(cout_10__BAR), .Q(sumout[10]) );
  OA21X1 U66 ( .IN1(in2[11]), .IN2(in1[11]), .IN3(cout_11__BAR), .Q(sumout[11]) );
  OA21X1 U67 ( .IN1(in2[12]), .IN2(in1[12]), .IN3(cout_12__BAR), .Q(sumout[12]) );
  OA21X1 U68 ( .IN1(in2[13]), .IN2(in1[13]), .IN3(cout_13__BAR), .Q(sumout[13]) );
  OA21X1 U69 ( .IN1(in2[14]), .IN2(in1[14]), .IN3(cout_14__BAR), .Q(sumout[14]) );
  OA21X1 U70 ( .IN1(in2[15]), .IN2(in1[15]), .IN3(cout_15__BAR), .Q(sumout[15]) );
  OA21X1 U71 ( .IN1(in2[16]), .IN2(in1[16]), .IN3(cout_16__BAR), .Q(sumout[16]) );
  OA21X1 U72 ( .IN1(in2[17]), .IN2(in1[17]), .IN3(cout_17__BAR), .Q(sumout[17]) );
  OA21X1 U73 ( .IN1(in2[18]), .IN2(in1[18]), .IN3(cout_18__BAR), .Q(sumout[18]) );
  OA21X1 U74 ( .IN1(in2[19]), .IN2(in1[19]), .IN3(cout_19__BAR), .Q(sumout[19]) );
  OA21X1 U75 ( .IN1(in2[20]), .IN2(in1[20]), .IN3(cout_20__BAR), .Q(sumout[20]) );
  OA21X1 U76 ( .IN1(in2[21]), .IN2(in1[21]), .IN3(cout_21__BAR), .Q(sumout[21]) );
  OA21X1 U77 ( .IN1(in2[22]), .IN2(in1[22]), .IN3(cout_22__BAR), .Q(sumout[22]) );
  OA21X1 U78 ( .IN1(in2[23]), .IN2(in1[23]), .IN3(cout_23__BAR), .Q(sumout[23]) );
  OA21X1 U79 ( .IN1(in2[24]), .IN2(in1[24]), .IN3(cout_24__BAR), .Q(sumout[24]) );
  OA21X1 U80 ( .IN1(in2[25]), .IN2(in1[25]), .IN3(cout_25__BAR), .Q(sumout[25]) );
  OA21X1 U81 ( .IN1(in2[26]), .IN2(in1[26]), .IN3(cout_26__BAR), .Q(sumout[26]) );
  OA21X1 U82 ( .IN1(in2[29]), .IN2(in1[29]), .IN3(cout_29__BAR), .Q(sumout[29]) );
  OA21X1 U83 ( .IN1(in2[31]), .IN2(in1[31]), .IN3(cout_31__BAR), .Q(sumout[31]) );
  OA21X1 U84 ( .IN1(in2[33]), .IN2(in1[33]), .IN3(cout_33__BAR), .Q(sumout[33]) );
  OA21X1 U85 ( .IN1(in2[35]), .IN2(in1[35]), .IN3(cout_35__BAR), .Q(sumout[35]) );
  OA21X1 U86 ( .IN1(in2[37]), .IN2(in1[37]), .IN3(cout_37__BAR), .Q(sumout[37]) );
  OA21X1 U87 ( .IN1(in2[39]), .IN2(in1[39]), .IN3(cout_39__BAR), .Q(sumout[39]) );
  OA21X1 U88 ( .IN1(in2[41]), .IN2(in1[41]), .IN3(cout_41__BAR), .Q(sumout[41]) );
  OA21X1 U89 ( .IN1(in2[43]), .IN2(in1[43]), .IN3(cout_43__BAR), .Q(sumout[43]) );
  OA21X1 U90 ( .IN1(in2[45]), .IN2(in1[45]), .IN3(cout_45__BAR), .Q(sumout[45]) );
  XOR2X1 U91 ( .IN1(in1[47]), .IN2(in2[47]), .Q(sumout[47]) );
endmodule


module csa51squ_62 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;


  AO222X1 U1 ( .IN1(in2[6]), .IN2(in3[6]), .IN3(in2[6]), .IN4(in1[6]), .IN5(
        in3[6]), .IN6(in1[6]), .Q(cout[6]) );
  FADDX1 U2 ( .A(in1[10]), .B(in2[10]), .CI(in3[10]), .CO(cout[10]), .S(
        sumout[10]) );
  FADDX1 U3 ( .A(in1[11]), .B(in2[11]), .CI(in3[11]), .CO(cout[11]), .S(
        sumout[11]) );
  FADDX1 U4 ( .A(in1[12]), .B(in2[12]), .CI(in3[12]), .CO(cout[12]), .S(
        sumout[12]) );
  FADDX1 U5 ( .A(in1[13]), .B(in2[13]), .CI(in3[13]), .CO(cout[13]), .S(
        sumout[13]) );
  FADDX1 U6 ( .A(in1[14]), .B(in2[14]), .CI(in3[14]), .CO(cout[14]), .S(
        sumout[14]) );
  FADDX1 U7 ( .A(in1[15]), .B(in2[15]), .CI(in3[15]), .CO(cout[15]), .S(
        sumout[15]) );
  FADDX1 U8 ( .A(in1[16]), .B(in2[16]), .CI(in3[16]), .CO(cout[16]), .S(
        sumout[16]) );
  FADDX1 U9 ( .A(in1[17]), .B(in2[17]), .CI(in3[17]), .CO(cout[17]), .S(
        sumout[17]) );
  FADDX1 U10 ( .A(in1[18]), .B(in2[18]), .CI(in3[18]), .CO(cout[18]), .S(
        sumout[18]) );
  FADDX1 U11 ( .A(in1[19]), .B(in2[19]), .CI(in3[19]), .CO(cout[19]), .S(
        sumout[19]) );
  FADDX1 U12 ( .A(in1[20]), .B(in2[20]), .CI(in3[20]), .CO(cout[20]), .S(
        sumout[20]) );
  FADDX1 U13 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U14 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U15 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U16 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U17 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U18 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U19 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U20 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U21 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U22 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U23 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U24 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
  FADDX1 U25 ( .A(in1[33]), .B(in2[33]), .CI(in3[33]), .CO(cout[33]), .S(
        sumout[33]) );
  FADDX1 U26 ( .A(in1[34]), .B(in2[34]), .CI(in3[34]), .CO(cout[34]), .S(
        sumout[34]) );
  FADDX1 U27 ( .A(in1[35]), .B(in2[35]), .CI(in3[35]), .CO(cout[35]), .S(
        sumout[35]) );
  FADDX1 U28 ( .A(in1[36]), .B(in2[36]), .CI(in3[36]), .CO(cout[36]), .S(
        sumout[36]) );
  FADDX1 U29 ( .A(in1[37]), .B(in2[37]), .CI(in3[37]), .CO(cout[37]), .S(
        sumout[37]) );
  FADDX1 U30 ( .A(in1[38]), .B(in2[38]), .CI(in3[38]), .CO(cout[38]), .S(
        sumout[38]) );
  FADDX1 U31 ( .A(in1[39]), .B(in2[39]), .CI(in3[39]), .CO(cout[39]), .S(
        sumout[39]) );
  FADDX1 U32 ( .A(in1[40]), .B(in2[40]), .CI(in3[40]), .CO(cout[40]), .S(
        sumout[40]) );
  FADDX1 U33 ( .A(in1[41]), .B(in2[41]), .CI(in3[41]), .CO(cout[41]), .S(
        sumout[41]) );
  FADDX1 U34 ( .A(in1[42]), .B(in2[42]), .CI(in3[42]), .CO(cout[42]), .S(
        sumout[42]) );
  FADDX1 U35 ( .A(in1[43]), .B(in2[43]), .CI(in3[43]), .CO(cout[43]), .S(
        sumout[43]) );
  FADDX1 U36 ( .A(in1[44]), .B(in2[44]), .CI(in3[44]), .CO(cout[44]), .S(
        sumout[44]) );
  FADDX1 U37 ( .A(in1[45]), .B(in2[45]), .CI(in3[45]), .CO(cout[45]), .S(
        sumout[45]) );
  FADDX1 U38 ( .A(in1[46]), .B(in2[46]), .CI(in3[46]), .CO(cout[46]), .S(
        sumout[46]) );
  XOR3X1 U39 ( .IN1(in2[47]), .IN2(in3[47]), .IN3(in1[47]), .Q(sumout[47]) );
  FADDX1 U40 ( .A(in1[7]), .B(in2[7]), .CI(in3[7]), .CO(cout[7]), .S(sumout[7]) );
  FADDX1 U41 ( .A(in1[8]), .B(in2[8]), .CI(in3[8]), .CO(cout[8]), .S(sumout[8]) );
  FADDX1 U42 ( .A(in1[9]), .B(in2[9]), .CI(in3[9]), .CO(cout[9]), .S(sumout[9]) );
endmodule


module csa51squ_63 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14;

  AND2X1 U1 ( .IN1(in2[7]), .IN2(in1[7]), .Q(cout[7]) );
  NOR2X0 U2 ( .IN1(in2[7]), .IN2(in1[7]), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(cout[7]), .QN(sumout[7]) );
  AND2X1 U4 ( .IN1(in2[8]), .IN2(in1[8]), .Q(cout[8]) );
  NOR2X0 U5 ( .IN1(in2[8]), .IN2(in1[8]), .QN(n2) );
  NOR2X0 U6 ( .IN1(n2), .IN2(cout[8]), .QN(sumout[8]) );
  AND2X1 U7 ( .IN1(in2[9]), .IN2(in1[9]), .Q(cout[9]) );
  NOR2X0 U8 ( .IN1(in2[9]), .IN2(in1[9]), .QN(n3) );
  NOR2X0 U9 ( .IN1(n3), .IN2(cout[9]), .QN(sumout[9]) );
  AND2X1 U10 ( .IN1(in2[10]), .IN2(in1[10]), .Q(cout[10]) );
  NOR2X0 U11 ( .IN1(in2[10]), .IN2(in1[10]), .QN(n4) );
  NOR2X0 U12 ( .IN1(n4), .IN2(cout[10]), .QN(sumout[10]) );
  AND2X1 U13 ( .IN1(in2[11]), .IN2(in1[11]), .Q(cout[11]) );
  NOR2X0 U14 ( .IN1(in2[11]), .IN2(in1[11]), .QN(n5) );
  NOR2X0 U15 ( .IN1(n5), .IN2(cout[11]), .QN(sumout[11]) );
  AND2X1 U16 ( .IN1(in2[12]), .IN2(in1[12]), .Q(cout[12]) );
  NOR2X0 U17 ( .IN1(in2[12]), .IN2(in1[12]), .QN(n6) );
  NOR2X0 U18 ( .IN1(n6), .IN2(cout[12]), .QN(sumout[12]) );
  AND2X1 U19 ( .IN1(in3[40]), .IN2(in2[40]), .Q(cout[40]) );
  NOR2X0 U20 ( .IN1(in3[40]), .IN2(in2[40]), .QN(n7) );
  NOR2X0 U21 ( .IN1(n7), .IN2(cout[40]), .QN(sumout[40]) );
  AND2X1 U22 ( .IN1(in3[41]), .IN2(in2[41]), .Q(cout[41]) );
  NOR2X0 U23 ( .IN1(in3[41]), .IN2(in2[41]), .QN(n8) );
  NOR2X0 U24 ( .IN1(n8), .IN2(cout[41]), .QN(sumout[41]) );
  AND2X1 U25 ( .IN1(in3[42]), .IN2(in2[42]), .Q(cout[42]) );
  NOR2X0 U26 ( .IN1(in3[42]), .IN2(in2[42]), .QN(n9) );
  NOR2X0 U27 ( .IN1(n9), .IN2(cout[42]), .QN(sumout[42]) );
  AND2X1 U28 ( .IN1(in3[43]), .IN2(in2[43]), .Q(cout[43]) );
  NOR2X0 U29 ( .IN1(in3[43]), .IN2(in2[43]), .QN(n10) );
  NOR2X0 U30 ( .IN1(n10), .IN2(cout[43]), .QN(sumout[43]) );
  AND2X1 U31 ( .IN1(in3[44]), .IN2(in2[44]), .Q(cout[44]) );
  NOR2X0 U32 ( .IN1(in3[44]), .IN2(in2[44]), .QN(n11) );
  NOR2X0 U33 ( .IN1(n11), .IN2(cout[44]), .QN(sumout[44]) );
  AND2X1 U34 ( .IN1(in3[45]), .IN2(in2[45]), .Q(cout[45]) );
  NOR2X0 U35 ( .IN1(in3[45]), .IN2(in2[45]), .QN(n12) );
  NOR2X0 U36 ( .IN1(n12), .IN2(cout[45]), .QN(sumout[45]) );
  AND2X1 U37 ( .IN1(in3[46]), .IN2(in2[46]), .Q(cout[46]) );
  NOR2X0 U38 ( .IN1(in3[46]), .IN2(in2[46]), .QN(n13) );
  NOR2X0 U39 ( .IN1(n13), .IN2(cout[46]), .QN(sumout[46]) );
  INVX0 U40 ( .INP(in3[47]), .ZN(sumout[47]) );
  AND2X1 U41 ( .IN1(in2[5]), .IN2(in1[5]), .Q(cout[5]) );
  AND2X1 U42 ( .IN1(in2[6]), .IN2(in1[6]), .Q(cout[6]) );
  NOR2X0 U43 ( .IN1(in2[6]), .IN2(in1[6]), .QN(n14) );
  NOR2X0 U44 ( .IN1(n14), .IN2(cout[6]), .QN(sumout[6]) );
  FADDX1 U45 ( .A(in1[13]), .B(in2[13]), .CI(in3[13]), .CO(cout[13]), .S(
        sumout[13]) );
  FADDX1 U46 ( .A(in1[14]), .B(in2[14]), .CI(in3[14]), .CO(cout[14]), .S(
        sumout[14]) );
  FADDX1 U47 ( .A(in1[15]), .B(in2[15]), .CI(in3[15]), .CO(cout[15]), .S(
        sumout[15]) );
  FADDX1 U48 ( .A(in1[16]), .B(in2[16]), .CI(in3[16]), .CO(cout[16]), .S(
        sumout[16]) );
  FADDX1 U49 ( .A(in1[17]), .B(in2[17]), .CI(in3[17]), .CO(cout[17]), .S(
        sumout[17]) );
  FADDX1 U50 ( .A(in1[18]), .B(in2[18]), .CI(in3[18]), .CO(cout[18]), .S(
        sumout[18]) );
  FADDX1 U51 ( .A(in1[19]), .B(in2[19]), .CI(in3[19]), .CO(cout[19]), .S(
        sumout[19]) );
  FADDX1 U52 ( .A(in1[20]), .B(in2[20]), .CI(in3[20]), .CO(cout[20]), .S(
        sumout[20]) );
  FADDX1 U53 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U54 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U55 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U56 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U57 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U58 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U59 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U60 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U61 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U62 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U63 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U64 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
  FADDX1 U65 ( .A(in1[33]), .B(in2[33]), .CI(in3[33]), .CO(cout[33]), .S(
        sumout[33]) );
  FADDX1 U66 ( .A(in1[34]), .B(in2[34]), .CI(in3[34]), .CO(cout[34]), .S(
        sumout[34]) );
  FADDX1 U67 ( .A(in1[35]), .B(in2[35]), .CI(in3[35]), .CO(cout[35]), .S(
        sumout[35]) );
  FADDX1 U68 ( .A(in1[36]), .B(in2[36]), .CI(in3[36]), .CO(cout[36]), .S(
        sumout[36]) );
  FADDX1 U69 ( .A(in1[37]), .B(in2[37]), .CI(in3[37]), .CO(cout[37]), .S(
        sumout[37]) );
  FADDX1 U70 ( .A(in1[38]), .B(in2[38]), .CI(in3[38]), .CO(cout[38]), .S(
        sumout[38]) );
  FADDX1 U71 ( .A(in1[39]), .B(in2[39]), .CI(in3[39]), .CO(cout[39]), .S(
        sumout[39]) );
endmodule


module csa51squ_64 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17;

  NBUFFX2 U1 ( .INP(in1[6]), .Z(sumout[6]) );
  NBUFFX2 U2 ( .INP(in1[7]), .Z(sumout[7]) );
  NBUFFX2 U3 ( .INP(in1[8]), .Z(sumout[8]) );
  NBUFFX2 U4 ( .INP(in1[9]), .Z(sumout[9]) );
  NBUFFX2 U5 ( .INP(in1[10]), .Z(sumout[10]) );
  NBUFFX2 U6 ( .INP(in1[11]), .Z(sumout[11]) );
  AND2X1 U7 ( .IN1(in3[13]), .IN2(in1[13]), .Q(cout[13]) );
  NOR2X0 U8 ( .IN1(in3[13]), .IN2(in1[13]), .QN(n7) );
  NOR2X0 U9 ( .IN1(n7), .IN2(cout[13]), .QN(sumout[13]) );
  AND2X1 U10 ( .IN1(in3[15]), .IN2(in1[15]), .Q(cout[15]) );
  NOR2X0 U11 ( .IN1(in3[15]), .IN2(in1[15]), .QN(n8) );
  NOR2X0 U12 ( .IN1(n8), .IN2(cout[15]), .QN(sumout[15]) );
  AND2X1 U13 ( .IN1(in3[17]), .IN2(in1[17]), .Q(cout[17]) );
  NOR2X0 U14 ( .IN1(in3[17]), .IN2(in1[17]), .QN(n9) );
  NOR2X0 U15 ( .IN1(n9), .IN2(cout[17]), .QN(sumout[17]) );
  AND2X1 U16 ( .IN1(in3[43]), .IN2(in2[43]), .Q(cout[43]) );
  NOR2X0 U17 ( .IN1(in3[43]), .IN2(in2[43]), .QN(n10) );
  NOR2X0 U18 ( .IN1(n10), .IN2(cout[43]), .QN(sumout[43]) );
  AND2X1 U19 ( .IN1(in3[44]), .IN2(in2[44]), .Q(cout[44]) );
  NOR2X0 U20 ( .IN1(in3[44]), .IN2(in2[44]), .QN(n11) );
  NOR2X0 U21 ( .IN1(n11), .IN2(cout[44]), .QN(sumout[44]) );
  AND2X1 U22 ( .IN1(in3[45]), .IN2(in2[45]), .Q(cout[45]) );
  NOR2X0 U23 ( .IN1(in3[45]), .IN2(in2[45]), .QN(n12) );
  NOR2X0 U24 ( .IN1(n12), .IN2(cout[45]), .QN(sumout[45]) );
  AND2X1 U25 ( .IN1(in3[46]), .IN2(in2[46]), .Q(cout[46]) );
  NOR2X0 U26 ( .IN1(in3[46]), .IN2(in2[46]), .QN(n13) );
  NOR2X0 U27 ( .IN1(n13), .IN2(cout[46]), .QN(sumout[46]) );
  XOR2X1 U28 ( .IN1(in3[47]), .IN2(in2[47]), .Q(sumout[47]) );
  AND2X1 U29 ( .IN1(in3[12]), .IN2(in1[12]), .Q(cout[12]) );
  NOR2X0 U30 ( .IN1(in3[12]), .IN2(in1[12]), .QN(n14) );
  NOR2X0 U31 ( .IN1(n14), .IN2(cout[12]), .QN(sumout[12]) );
  AND2X1 U32 ( .IN1(in3[14]), .IN2(in1[14]), .Q(cout[14]) );
  NOR2X0 U33 ( .IN1(in3[14]), .IN2(in1[14]), .QN(n15) );
  NOR2X0 U34 ( .IN1(n15), .IN2(cout[14]), .QN(sumout[14]) );
  AND2X1 U35 ( .IN1(in3[16]), .IN2(in1[16]), .Q(cout[16]) );
  NOR2X0 U36 ( .IN1(in3[16]), .IN2(in1[16]), .QN(n16) );
  NOR2X0 U37 ( .IN1(n16), .IN2(cout[16]), .QN(sumout[16]) );
  AND2X1 U38 ( .IN1(in3[18]), .IN2(in1[18]), .Q(cout[18]) );
  NOR2X0 U39 ( .IN1(in3[18]), .IN2(in1[18]), .QN(n17) );
  NOR2X0 U40 ( .IN1(n17), .IN2(cout[18]), .QN(sumout[18]) );
  FADDX1 U41 ( .A(in1[19]), .B(in2[19]), .CI(in3[19]), .CO(cout[19]), .S(
        sumout[19]) );
  FADDX1 U42 ( .A(in1[20]), .B(in2[20]), .CI(in3[20]), .CO(cout[20]), .S(
        sumout[20]) );
  FADDX1 U43 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U44 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U45 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U46 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U47 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U48 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U49 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U50 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U51 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U52 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U53 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U54 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
  FADDX1 U55 ( .A(in1[33]), .B(in2[33]), .CI(in3[33]), .CO(cout[33]), .S(
        sumout[33]) );
  FADDX1 U56 ( .A(in1[34]), .B(in2[34]), .CI(in3[34]), .CO(cout[34]), .S(
        sumout[34]) );
  FADDX1 U57 ( .A(in1[35]), .B(in2[35]), .CI(in3[35]), .CO(cout[35]), .S(
        sumout[35]) );
  FADDX1 U58 ( .A(in1[36]), .B(in2[36]), .CI(in3[36]), .CO(cout[36]), .S(
        sumout[36]) );
  FADDX1 U59 ( .A(in1[37]), .B(in2[37]), .CI(in3[37]), .CO(cout[37]), .S(
        sumout[37]) );
  FADDX1 U60 ( .A(in1[38]), .B(in2[38]), .CI(in3[38]), .CO(cout[38]), .S(
        sumout[38]) );
  FADDX1 U61 ( .A(in1[39]), .B(in2[39]), .CI(in3[39]), .CO(cout[39]), .S(
        sumout[39]) );
  FADDX1 U62 ( .A(in1[40]), .B(in2[40]), .CI(in3[40]), .CO(cout[40]), .S(
        sumout[40]) );
  FADDX1 U63 ( .A(in1[41]), .B(in2[41]), .CI(in3[41]), .CO(cout[41]), .S(
        sumout[41]) );
  FADDX1 U64 ( .A(in1[42]), .B(in2[42]), .CI(in3[42]), .CO(cout[42]), .S(
        sumout[42]) );
endmodule


module csa51squ_65 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19;

  NBUFFX2 U1 ( .INP(in2[46]), .Z(sumout[46]) );
  NBUFFX2 U2 ( .INP(in2[45]), .Z(sumout[45]) );
  NBUFFX2 U3 ( .INP(in2[44]), .Z(sumout[44]) );
  NBUFFX2 U4 ( .INP(in2[43]), .Z(sumout[43]) );
  NBUFFX2 U5 ( .INP(in2[42]), .Z(sumout[42]) );
  NBUFFX2 U6 ( .INP(in2[41]), .Z(sumout[41]) );
  NBUFFX2 U7 ( .INP(in2[40]), .Z(sumout[40]) );
  NBUFFX2 U8 ( .INP(in2[39]), .Z(sumout[39]) );
  AND2X1 U9 ( .IN1(in2[7]), .IN2(in1[7]), .Q(cout[7]) );
  NOR2X0 U10 ( .IN1(in2[7]), .IN2(in1[7]), .QN(n9) );
  NOR2X0 U11 ( .IN1(n9), .IN2(cout[7]), .QN(sumout[7]) );
  AND2X1 U12 ( .IN1(in2[8]), .IN2(in1[8]), .Q(cout[8]) );
  NOR2X0 U13 ( .IN1(in2[8]), .IN2(in1[8]), .QN(n10) );
  NOR2X0 U14 ( .IN1(n10), .IN2(cout[8]), .QN(sumout[8]) );
  AND2X1 U15 ( .IN1(in2[9]), .IN2(in1[9]), .Q(cout[9]) );
  NOR2X0 U16 ( .IN1(in2[9]), .IN2(in1[9]), .QN(n11) );
  NOR2X0 U17 ( .IN1(n11), .IN2(cout[9]), .QN(sumout[9]) );
  AND2X1 U18 ( .IN1(in3[33]), .IN2(in2[33]), .Q(cout[33]) );
  NOR2X0 U19 ( .IN1(in3[33]), .IN2(in2[33]), .QN(n12) );
  NOR2X0 U20 ( .IN1(n12), .IN2(cout[33]), .QN(sumout[33]) );
  AND2X1 U21 ( .IN1(in3[34]), .IN2(in2[34]), .Q(cout[34]) );
  NOR2X0 U22 ( .IN1(in3[34]), .IN2(in2[34]), .QN(n13) );
  NOR2X0 U23 ( .IN1(n13), .IN2(cout[34]), .QN(sumout[34]) );
  AND2X1 U24 ( .IN1(in3[35]), .IN2(in2[35]), .Q(cout[35]) );
  NOR2X0 U25 ( .IN1(in3[35]), .IN2(in2[35]), .QN(n14) );
  NOR2X0 U26 ( .IN1(n14), .IN2(cout[35]), .QN(sumout[35]) );
  AND2X1 U27 ( .IN1(in3[36]), .IN2(in2[36]), .Q(cout[36]) );
  NOR2X0 U28 ( .IN1(in3[36]), .IN2(in2[36]), .QN(n15) );
  NOR2X0 U29 ( .IN1(n15), .IN2(cout[36]), .QN(sumout[36]) );
  AND2X1 U30 ( .IN1(in3[37]), .IN2(in2[37]), .Q(cout[37]) );
  NOR2X0 U31 ( .IN1(in3[37]), .IN2(in2[37]), .QN(n16) );
  NOR2X0 U32 ( .IN1(n16), .IN2(cout[37]), .QN(sumout[37]) );
  AND2X1 U33 ( .IN1(in3[38]), .IN2(in2[38]), .Q(cout[38]) );
  NOR2X0 U34 ( .IN1(in3[38]), .IN2(in2[38]), .QN(n17) );
  NOR2X0 U35 ( .IN1(n17), .IN2(cout[38]), .QN(sumout[38]) );
  AND2X1 U36 ( .IN1(in2[4]), .IN2(in1[4]), .Q(cout[4]) );
  AND2X1 U37 ( .IN1(in2[5]), .IN2(in1[5]), .Q(cout[5]) );
  NOR2X0 U38 ( .IN1(in2[5]), .IN2(in1[5]), .QN(n18) );
  NOR2X0 U39 ( .IN1(n18), .IN2(cout[5]), .QN(sumout[5]) );
  AND2X1 U40 ( .IN1(in2[6]), .IN2(in1[6]), .Q(cout[6]) );
  NOR2X0 U41 ( .IN1(in2[6]), .IN2(in1[6]), .QN(n19) );
  NOR2X0 U42 ( .IN1(n19), .IN2(cout[6]), .QN(sumout[6]) );
  FADDX1 U43 ( .A(in1[10]), .B(in2[10]), .CI(in3[10]), .CO(cout[10]), .S(
        sumout[10]) );
  FADDX1 U44 ( .A(in1[11]), .B(in2[11]), .CI(in3[11]), .CO(cout[11]), .S(
        sumout[11]) );
  FADDX1 U45 ( .A(in1[12]), .B(in2[12]), .CI(in3[12]), .CO(cout[12]), .S(
        sumout[12]) );
  FADDX1 U46 ( .A(in1[13]), .B(in2[13]), .CI(in3[13]), .CO(cout[13]), .S(
        sumout[13]) );
  FADDX1 U47 ( .A(in1[14]), .B(in2[14]), .CI(in3[14]), .CO(cout[14]), .S(
        sumout[14]) );
  FADDX1 U48 ( .A(in1[15]), .B(in2[15]), .CI(in3[15]), .CO(cout[15]), .S(
        sumout[15]) );
  FADDX1 U49 ( .A(in1[16]), .B(in2[16]), .CI(in3[16]), .CO(cout[16]), .S(
        sumout[16]) );
  FADDX1 U50 ( .A(in1[17]), .B(in2[17]), .CI(in3[17]), .CO(cout[17]), .S(
        sumout[17]) );
  FADDX1 U51 ( .A(in1[18]), .B(in2[18]), .CI(in3[18]), .CO(cout[18]), .S(
        sumout[18]) );
  FADDX1 U52 ( .A(in1[19]), .B(in2[19]), .CI(in3[19]), .CO(cout[19]), .S(
        sumout[19]) );
  FADDX1 U53 ( .A(in1[20]), .B(in2[20]), .CI(in3[20]), .CO(cout[20]), .S(
        sumout[20]) );
  FADDX1 U54 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U55 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U56 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U57 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U58 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U59 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U60 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U61 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U62 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U63 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U64 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U65 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
endmodule


module csa51squ_66 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n7, n8, n9, n10, n11, n12, n13;

  NBUFFX2 U1 ( .INP(in1[12]), .Z(sumout[12]) );
  NBUFFX2 U2 ( .INP(in1[13]), .Z(sumout[13]) );
  NBUFFX2 U3 ( .INP(in1[14]), .Z(sumout[14]) );
  NBUFFX2 U4 ( .INP(in1[15]), .Z(sumout[15]) );
  NBUFFX2 U5 ( .INP(in1[16]), .Z(sumout[16]) );
  NBUFFX2 U6 ( .INP(in1[17]), .Z(sumout[17]) );
  AND2X1 U7 ( .IN1(in3[19]), .IN2(in1[19]), .Q(cout[19]) );
  NOR2X0 U8 ( .IN1(in3[19]), .IN2(in1[19]), .QN(n7) );
  NOR2X0 U9 ( .IN1(n7), .IN2(cout[19]), .QN(sumout[19]) );
  AND2X1 U10 ( .IN1(in3[44]), .IN2(in2[44]), .Q(cout[44]) );
  NOR2X0 U11 ( .IN1(in3[44]), .IN2(in2[44]), .QN(n8) );
  NOR2X0 U12 ( .IN1(n8), .IN2(cout[44]), .QN(sumout[44]) );
  AND2X1 U13 ( .IN1(in3[45]), .IN2(in2[45]), .Q(cout[45]) );
  NOR2X0 U14 ( .IN1(in3[45]), .IN2(in2[45]), .QN(n9) );
  NOR2X0 U15 ( .IN1(n9), .IN2(cout[45]), .QN(sumout[45]) );
  AND2X1 U16 ( .IN1(in3[46]), .IN2(in2[46]), .Q(cout[46]) );
  NOR2X0 U17 ( .IN1(in3[46]), .IN2(in2[46]), .QN(n10) );
  NOR2X0 U18 ( .IN1(n10), .IN2(cout[46]), .QN(sumout[46]) );
  XOR2X1 U19 ( .IN1(in3[47]), .IN2(in2[47]), .Q(sumout[47]) );
  AND2X1 U20 ( .IN1(in3[18]), .IN2(in1[18]), .Q(cout[18]) );
  NOR2X0 U21 ( .IN1(in3[18]), .IN2(in1[18]), .QN(n11) );
  NOR2X0 U22 ( .IN1(n11), .IN2(cout[18]), .QN(sumout[18]) );
  AND2X1 U23 ( .IN1(in3[20]), .IN2(in1[20]), .Q(cout[20]) );
  NOR2X0 U24 ( .IN1(in3[20]), .IN2(in1[20]), .QN(n12) );
  NOR2X0 U25 ( .IN1(n12), .IN2(cout[20]), .QN(sumout[20]) );
  INVX0 U26 ( .INP(in1[42]), .ZN(n13) );
  FADDX1 U27 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U28 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U29 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U30 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U31 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U32 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U33 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U34 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U35 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U36 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U37 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U38 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
  FADDX1 U39 ( .A(in1[33]), .B(in2[33]), .CI(in3[33]), .CO(cout[33]), .S(
        sumout[33]) );
  FADDX1 U40 ( .A(in1[34]), .B(in2[34]), .CI(in3[34]), .CO(cout[34]), .S(
        sumout[34]) );
  FADDX1 U41 ( .A(in1[35]), .B(in2[35]), .CI(in3[35]), .CO(cout[35]), .S(
        sumout[35]) );
  FADDX1 U42 ( .A(in1[36]), .B(in2[36]), .CI(in3[36]), .CO(cout[36]), .S(
        sumout[36]) );
  FADDX1 U43 ( .A(in1[37]), .B(in2[37]), .CI(in3[37]), .CO(cout[37]), .S(
        sumout[37]) );
  FADDX1 U44 ( .A(in1[38]), .B(in2[38]), .CI(in3[38]), .CO(cout[38]), .S(
        sumout[38]) );
  FADDX1 U45 ( .A(in1[39]), .B(in2[39]), .CI(in3[39]), .CO(cout[39]), .S(
        sumout[39]) );
  FADDX1 U46 ( .A(in1[40]), .B(in2[40]), .CI(in3[40]), .CO(cout[40]), .S(
        sumout[40]) );
  FADDX1 U47 ( .A(in1[41]), .B(in2[41]), .CI(in3[41]), .CO(cout[41]), .S(
        sumout[41]) );
  FADDX1 U48 ( .A(in1[42]), .B(in2[42]), .CI(in3[42]), .CO(cout[42]), .S(
        sumout[42]) );
  FADDX1 U49 ( .A(in2[43]), .B(in3[43]), .CI(n13), .CO(cout[43]), .S(
        sumout[43]) );
endmodule


module csa51squ_67 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n9, n10, n11, n12, n13, n14, n15;

  NBUFFX2 U1 ( .INP(in2[6]), .Z(sumout[6]) );
  NBUFFX2 U2 ( .INP(in2[7]), .Z(sumout[7]) );
  NBUFFX2 U3 ( .INP(in2[8]), .Z(sumout[8]) );
  NBUFFX2 U4 ( .INP(in3[42]), .Z(sumout[42]) );
  NBUFFX2 U5 ( .INP(in3[41]), .Z(sumout[41]) );
  NBUFFX2 U6 ( .INP(in3[39]), .Z(sumout[39]) );
  NBUFFX2 U7 ( .INP(in3[38]), .Z(sumout[38]) );
  NBUFFX2 U8 ( .INP(in3[40]), .Z(sumout[40]) );
  AND2X1 U9 ( .IN1(in2[13]), .IN2(in1[13]), .Q(cout[13]) );
  NOR2X0 U10 ( .IN1(in2[13]), .IN2(in1[13]), .QN(n9) );
  NOR2X0 U11 ( .IN1(n9), .IN2(cout[13]), .QN(sumout[13]) );
  AND2X1 U12 ( .IN1(in2[37]), .IN2(in3[37]), .Q(cout[37]) );
  INVX0 U13 ( .INP(in2[37]), .ZN(n15) );
  MUX21X1 U14 ( .IN1(in2[37]), .IN2(n15), .S(in3[37]), .Q(sumout[37]) );
  AND2X1 U15 ( .IN1(in2[9]), .IN2(in1[9]), .Q(cout[9]) );
  NOR2X0 U16 ( .IN1(in2[9]), .IN2(in1[9]), .QN(n10) );
  NOR2X0 U17 ( .IN1(n10), .IN2(cout[9]), .QN(sumout[9]) );
  AND2X1 U18 ( .IN1(in2[10]), .IN2(in1[10]), .Q(cout[10]) );
  NOR2X0 U19 ( .IN1(in2[10]), .IN2(in1[10]), .QN(n11) );
  NOR2X0 U20 ( .IN1(n11), .IN2(cout[10]), .QN(sumout[10]) );
  AND2X1 U21 ( .IN1(in2[11]), .IN2(in1[11]), .Q(cout[11]) );
  NOR2X0 U22 ( .IN1(in2[11]), .IN2(in1[11]), .QN(n12) );
  NOR2X0 U23 ( .IN1(n12), .IN2(cout[11]), .QN(sumout[11]) );
  AND2X1 U24 ( .IN1(in2[12]), .IN2(in1[12]), .Q(cout[12]) );
  NOR2X0 U25 ( .IN1(in2[12]), .IN2(in1[12]), .QN(n13) );
  NOR2X0 U26 ( .IN1(n13), .IN2(cout[12]), .QN(sumout[12]) );
  AND2X1 U27 ( .IN1(in2[14]), .IN2(in1[14]), .Q(cout[14]) );
  NOR2X0 U28 ( .IN1(in2[14]), .IN2(in1[14]), .QN(n14) );
  NOR2X0 U29 ( .IN1(n14), .IN2(cout[14]), .QN(sumout[14]) );
  FADDX1 U30 ( .A(in1[15]), .B(in2[15]), .CI(in3[15]), .CO(cout[15]), .S(
        sumout[15]) );
  FADDX1 U31 ( .A(in1[16]), .B(in2[16]), .CI(in3[16]), .CO(cout[16]), .S(
        sumout[16]) );
  FADDX1 U32 ( .A(in1[17]), .B(in2[17]), .CI(in3[17]), .CO(cout[17]), .S(
        sumout[17]) );
  FADDX1 U33 ( .A(in1[18]), .B(in2[18]), .CI(in3[18]), .CO(cout[18]), .S(
        sumout[18]) );
  FADDX1 U34 ( .A(in1[19]), .B(in2[19]), .CI(in3[19]), .CO(cout[19]), .S(
        sumout[19]) );
  FADDX1 U35 ( .A(in1[20]), .B(in2[20]), .CI(in3[20]), .CO(cout[20]), .S(
        sumout[20]) );
  FADDX1 U36 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U37 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U38 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U39 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U40 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U41 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U42 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U43 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U44 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U45 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U46 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U47 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
  FADDX1 U48 ( .A(in1[33]), .B(in2[33]), .CI(in3[33]), .CO(cout[33]), .S(
        sumout[33]) );
  FADDX1 U49 ( .A(in1[34]), .B(in2[34]), .CI(in3[34]), .CO(cout[34]), .S(
        sumout[34]) );
  FADDX1 U50 ( .A(in1[35]), .B(in2[35]), .CI(in3[35]), .CO(cout[35]), .S(
        sumout[35]) );
  FADDX1 U51 ( .A(in1[36]), .B(in3[36]), .CI(n15), .CO(cout[36]), .S(
        sumout[36]) );
endmodule


module csa51squ_68 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36;

  NBUFFX2 U1 ( .INP(in3[46]), .Z(sumout[46]) );
  NBUFFX2 U2 ( .INP(in3[45]), .Z(sumout[45]) );
  NBUFFX2 U3 ( .INP(in3[44]), .Z(sumout[44]) );
  NBUFFX2 U4 ( .INP(in3[43]), .Z(sumout[43]) );
  NBUFFX2 U5 ( .INP(in3[42]), .Z(sumout[42]) );
  NBUFFX2 U6 ( .INP(in3[33]), .Z(sumout[33]) );
  NBUFFX2 U7 ( .INP(in3[32]), .Z(sumout[32]) );
  NBUFFX2 U8 ( .INP(in3[37]), .Z(sumout[37]) );
  NBUFFX2 U9 ( .INP(in3[36]), .Z(sumout[36]) );
  NBUFFX2 U10 ( .INP(in3[35]), .Z(sumout[35]) );
  NBUFFX2 U11 ( .INP(in3[34]), .Z(sumout[34]) );
  NBUFFX2 U12 ( .INP(in3[41]), .Z(sumout[41]) );
  NBUFFX2 U13 ( .INP(in3[40]), .Z(sumout[40]) );
  NBUFFX2 U14 ( .INP(in3[39]), .Z(sumout[39]) );
  NBUFFX2 U15 ( .INP(in3[38]), .Z(sumout[38]) );
  AND2X1 U16 ( .IN1(in2[31]), .IN2(in3[31]), .Q(cout[31]) );
  INVX0 U17 ( .INP(in2[31]), .ZN(n36) );
  MUX21X1 U18 ( .IN1(in2[31]), .IN2(n36), .S(in3[31]), .Q(sumout[31]) );
  AND2X1 U19 ( .IN1(in2[3]), .IN2(in1[3]), .Q(cout[3]) );
  AND2X1 U20 ( .IN1(in2[4]), .IN2(in1[4]), .Q(cout[4]) );
  NOR2X0 U21 ( .IN1(in2[4]), .IN2(in1[4]), .QN(n16) );
  NOR2X0 U22 ( .IN1(n16), .IN2(cout[4]), .QN(sumout[4]) );
  AND2X1 U23 ( .IN1(in2[5]), .IN2(in1[5]), .Q(cout[5]) );
  NOR2X0 U24 ( .IN1(in2[5]), .IN2(in1[5]), .QN(n17) );
  NOR2X0 U25 ( .IN1(n17), .IN2(cout[5]), .QN(sumout[5]) );
  AND2X1 U26 ( .IN1(in2[6]), .IN2(in1[6]), .Q(cout[6]) );
  NOR2X0 U27 ( .IN1(in2[6]), .IN2(in1[6]), .QN(n18) );
  NOR2X0 U28 ( .IN1(n18), .IN2(cout[6]), .QN(sumout[6]) );
  AND2X1 U29 ( .IN1(in2[7]), .IN2(in1[7]), .Q(cout[7]) );
  NOR2X0 U30 ( .IN1(in2[7]), .IN2(in1[7]), .QN(n19) );
  NOR2X0 U31 ( .IN1(n19), .IN2(cout[7]), .QN(sumout[7]) );
  AND2X1 U32 ( .IN1(in2[8]), .IN2(in1[8]), .Q(cout[8]) );
  NOR2X0 U33 ( .IN1(in2[8]), .IN2(in1[8]), .QN(n20) );
  NOR2X0 U34 ( .IN1(n20), .IN2(cout[8]), .QN(sumout[8]) );
  AND2X1 U35 ( .IN1(in2[9]), .IN2(in1[9]), .Q(cout[9]) );
  NOR2X0 U36 ( .IN1(in2[9]), .IN2(in1[9]), .QN(n21) );
  NOR2X0 U37 ( .IN1(n21), .IN2(cout[9]), .QN(sumout[9]) );
  AND2X1 U38 ( .IN1(in2[10]), .IN2(in1[10]), .Q(cout[10]) );
  NOR2X0 U39 ( .IN1(in2[10]), .IN2(in1[10]), .QN(n22) );
  NOR2X0 U40 ( .IN1(n22), .IN2(cout[10]), .QN(sumout[10]) );
  AND2X1 U41 ( .IN1(in2[11]), .IN2(in1[11]), .Q(cout[11]) );
  NOR2X0 U42 ( .IN1(in2[11]), .IN2(in1[11]), .QN(n23) );
  NOR2X0 U43 ( .IN1(n23), .IN2(cout[11]), .QN(sumout[11]) );
  AND2X1 U44 ( .IN1(in2[12]), .IN2(in1[12]), .Q(cout[12]) );
  NOR2X0 U45 ( .IN1(in2[12]), .IN2(in1[12]), .QN(n24) );
  NOR2X0 U46 ( .IN1(n24), .IN2(cout[12]), .QN(sumout[12]) );
  AND2X1 U47 ( .IN1(in2[13]), .IN2(in1[13]), .Q(cout[13]) );
  NOR2X0 U48 ( .IN1(in2[13]), .IN2(in1[13]), .QN(n25) );
  NOR2X0 U49 ( .IN1(n25), .IN2(cout[13]), .QN(sumout[13]) );
  AND2X1 U50 ( .IN1(in2[14]), .IN2(in1[14]), .Q(cout[14]) );
  NOR2X0 U51 ( .IN1(in2[14]), .IN2(in1[14]), .QN(n26) );
  NOR2X0 U52 ( .IN1(n26), .IN2(cout[14]), .QN(sumout[14]) );
  AND2X1 U53 ( .IN1(in2[15]), .IN2(in1[15]), .Q(cout[15]) );
  NOR2X0 U54 ( .IN1(in2[15]), .IN2(in1[15]), .QN(n27) );
  NOR2X0 U55 ( .IN1(n27), .IN2(cout[15]), .QN(sumout[15]) );
  AND2X1 U56 ( .IN1(in2[16]), .IN2(in1[16]), .Q(cout[16]) );
  NOR2X0 U57 ( .IN1(in2[16]), .IN2(in1[16]), .QN(n28) );
  NOR2X0 U58 ( .IN1(n28), .IN2(cout[16]), .QN(sumout[16]) );
  AND2X1 U59 ( .IN1(in2[17]), .IN2(in1[17]), .Q(cout[17]) );
  NOR2X0 U60 ( .IN1(in2[17]), .IN2(in1[17]), .QN(n29) );
  NOR2X0 U61 ( .IN1(n29), .IN2(cout[17]), .QN(sumout[17]) );
  AND2X1 U62 ( .IN1(in2[18]), .IN2(in1[18]), .Q(cout[18]) );
  NOR2X0 U63 ( .IN1(in2[18]), .IN2(in1[18]), .QN(n30) );
  NOR2X0 U64 ( .IN1(n30), .IN2(cout[18]), .QN(sumout[18]) );
  AND2X1 U65 ( .IN1(in2[19]), .IN2(in1[19]), .Q(cout[19]) );
  NOR2X0 U66 ( .IN1(in2[19]), .IN2(in1[19]), .QN(n31) );
  NOR2X0 U67 ( .IN1(n31), .IN2(cout[19]), .QN(sumout[19]) );
  AND2X1 U68 ( .IN1(in2[20]), .IN2(in1[20]), .Q(cout[20]) );
  NOR2X0 U69 ( .IN1(in2[20]), .IN2(in1[20]), .QN(n32) );
  NOR2X0 U70 ( .IN1(n32), .IN2(cout[20]), .QN(sumout[20]) );
  AND2X1 U71 ( .IN1(in2[21]), .IN2(in1[21]), .Q(cout[21]) );
  NOR2X0 U72 ( .IN1(in2[21]), .IN2(in1[21]), .QN(n33) );
  NOR2X0 U73 ( .IN1(n33), .IN2(cout[21]), .QN(sumout[21]) );
  AND2X1 U74 ( .IN1(in2[22]), .IN2(in1[22]), .Q(cout[22]) );
  NOR2X0 U75 ( .IN1(in2[22]), .IN2(in1[22]), .QN(n34) );
  NOR2X0 U76 ( .IN1(n34), .IN2(cout[22]), .QN(sumout[22]) );
  AND2X1 U77 ( .IN1(in2[23]), .IN2(in1[23]), .Q(cout[23]) );
  NOR2X0 U78 ( .IN1(in2[23]), .IN2(in1[23]), .QN(n35) );
  NOR2X0 U79 ( .IN1(n35), .IN2(cout[23]), .QN(sumout[23]) );
  FADDX1 U80 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U81 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U82 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U83 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U84 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U85 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U86 ( .A(in1[30]), .B(in3[30]), .CI(n36), .CO(cout[30]), .S(
        sumout[30]) );
endmodule


module csa51squ_69 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n3, n4, n5, n6, n7;

  NBUFFX2 U1 ( .INP(in1[18]), .Z(sumout[18]) );
  NBUFFX2 U2 ( .INP(in1[19]), .Z(sumout[19]) );
  AND2X1 U3 ( .IN1(in2[20]), .IN2(in1[20]), .Q(cout[20]) );
  NOR2X0 U4 ( .IN1(in2[20]), .IN2(in1[20]), .QN(n3) );
  NOR2X0 U5 ( .IN1(n3), .IN2(cout[20]), .QN(sumout[20]) );
  AND2X1 U6 ( .IN1(in2[21]), .IN2(in1[21]), .Q(cout[21]) );
  NOR2X0 U7 ( .IN1(in2[21]), .IN2(in1[21]), .QN(n4) );
  NOR2X0 U8 ( .IN1(n4), .IN2(cout[21]), .QN(sumout[21]) );
  AND2X1 U9 ( .IN1(in2[46]), .IN2(in3[46]), .Q(cout[46]) );
  NOR2X0 U10 ( .IN1(in2[46]), .IN2(in3[46]), .QN(n5) );
  NOR2X0 U11 ( .IN1(n5), .IN2(cout[46]), .QN(sumout[46]) );
  INVX0 U12 ( .INP(in2[46]), .ZN(n6) );
  MUX21X1 U13 ( .IN1(n6), .IN2(in2[46]), .S(in3[47]), .Q(sumout[47]) );
  INVX0 U14 ( .INP(in1[44]), .ZN(n7) );
  FADDX1 U15 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U16 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U17 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U18 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U19 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U20 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U21 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U22 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U23 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U24 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U25 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
  FADDX1 U26 ( .A(in1[33]), .B(in2[33]), .CI(in3[33]), .CO(cout[33]), .S(
        sumout[33]) );
  FADDX1 U27 ( .A(in1[34]), .B(in2[34]), .CI(in3[34]), .CO(cout[34]), .S(
        sumout[34]) );
  FADDX1 U28 ( .A(in1[35]), .B(in2[35]), .CI(in3[35]), .CO(cout[35]), .S(
        sumout[35]) );
  FADDX1 U29 ( .A(in1[36]), .B(in2[36]), .CI(in3[36]), .CO(cout[36]), .S(
        sumout[36]) );
  FADDX1 U30 ( .A(in1[37]), .B(in2[37]), .CI(in3[37]), .CO(cout[37]), .S(
        sumout[37]) );
  FADDX1 U31 ( .A(in1[38]), .B(in2[38]), .CI(in3[38]), .CO(cout[38]), .S(
        sumout[38]) );
  FADDX1 U32 ( .A(in1[39]), .B(in2[39]), .CI(in3[39]), .CO(cout[39]), .S(
        sumout[39]) );
  FADDX1 U33 ( .A(in1[40]), .B(in2[40]), .CI(in3[40]), .CO(cout[40]), .S(
        sumout[40]) );
  FADDX1 U34 ( .A(in1[41]), .B(in2[41]), .CI(in3[41]), .CO(cout[41]), .S(
        sumout[41]) );
  FADDX1 U35 ( .A(in1[42]), .B(in2[42]), .CI(in3[42]), .CO(cout[42]), .S(
        sumout[42]) );
  FADDX1 U36 ( .A(in1[43]), .B(in2[43]), .CI(in3[43]), .CO(cout[43]), .S(
        sumout[43]) );
  FADDX1 U37 ( .A(in1[44]), .B(in2[44]), .CI(in3[44]), .CO(cout[44]), .S(
        sumout[44]) );
  FADDX1 U38 ( .A(in2[45]), .B(in3[45]), .CI(n7), .CO(cout[45]), .S(sumout[45]) );
endmodule


module csa51squ_70 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n5, n6, n7, n8, n9, n10;

  AND2X1 U1 ( .IN1(in3[37]), .IN2(in2[37]), .Q(cout[37]) );
  NAND2X0 U2 ( .IN1(n5), .IN2(cout[39]), .QN(sumout[39]) );
  NAND2X0 U3 ( .IN1(in2[39]), .IN2(in3[39]), .QN(n5) );
  NBUFFX2 U4 ( .INP(in1[12]), .Z(sumout[12]) );
  NBUFFX2 U5 ( .INP(in1[13]), .Z(sumout[13]) );
  NBUFFX2 U6 ( .INP(in3[42]), .Z(sumout[42]) );
  XOR2X1 U7 ( .IN1(in2[37]), .IN2(in3[37]), .Q(sumout[37]) );
  OR2X1 U8 ( .IN1(in3[39]), .IN2(in2[39]), .Q(cout[39]) );
  AND2X1 U9 ( .IN1(in3[38]), .IN2(in2[38]), .Q(cout[38]) );
  NOR2X0 U10 ( .IN1(in3[38]), .IN2(in2[38]), .QN(n6) );
  NOR2X0 U11 ( .IN1(n6), .IN2(cout[38]), .QN(sumout[38]) );
  AND2X1 U12 ( .IN1(in2[14]), .IN2(in1[14]), .Q(cout[14]) );
  NOR2X0 U13 ( .IN1(in2[14]), .IN2(in1[14]), .QN(n7) );
  NOR2X0 U14 ( .IN1(n7), .IN2(cout[14]), .QN(sumout[14]) );
  AND2X1 U15 ( .IN1(in2[15]), .IN2(in1[15]), .Q(cout[15]) );
  NOR2X0 U16 ( .IN1(in2[15]), .IN2(in1[15]), .QN(n8) );
  NOR2X0 U17 ( .IN1(n8), .IN2(cout[15]), .QN(sumout[15]) );
  AND2X1 U18 ( .IN1(in2[40]), .IN2(in3[40]), .Q(cout[40]) );
  NOR2X0 U19 ( .IN1(in2[40]), .IN2(in3[40]), .QN(n9) );
  NOR2X0 U20 ( .IN1(n9), .IN2(cout[40]), .QN(sumout[40]) );
  INVX0 U21 ( .INP(in3[41]), .ZN(n10) );
  NOR2X0 U22 ( .IN1(in2[40]), .IN2(n10), .QN(cout[41]) );
  MUX21X1 U23 ( .IN1(n10), .IN2(in3[41]), .S(in2[40]), .Q(sumout[41]) );
  FADDX1 U24 ( .A(in1[16]), .B(in2[16]), .CI(in3[16]), .CO(cout[16]), .S(
        sumout[16]) );
  FADDX1 U25 ( .A(in1[17]), .B(in2[17]), .CI(in3[17]), .CO(cout[17]), .S(
        sumout[17]) );
  FADDX1 U26 ( .A(in1[18]), .B(in2[18]), .CI(in3[18]), .CO(cout[18]), .S(
        sumout[18]) );
  FADDX1 U27 ( .A(in1[19]), .B(in2[19]), .CI(in3[19]), .CO(cout[19]), .S(
        sumout[19]) );
  FADDX1 U28 ( .A(in1[20]), .B(in2[20]), .CI(in3[20]), .CO(cout[20]), .S(
        sumout[20]) );
  FADDX1 U29 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U30 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U31 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U32 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U33 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U34 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U35 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U36 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U37 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U38 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U39 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U40 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
  FADDX1 U41 ( .A(in1[33]), .B(in2[33]), .CI(in3[33]), .CO(cout[33]), .S(
        sumout[33]) );
  FADDX1 U42 ( .A(in1[34]), .B(in2[34]), .CI(in3[34]), .CO(cout[34]), .S(
        sumout[34]) );
  FADDX1 U43 ( .A(in1[35]), .B(in2[35]), .CI(in3[35]), .CO(cout[35]), .S(
        sumout[35]) );
  FADDX1 U44 ( .A(in1[36]), .B(in2[36]), .CI(in3[36]), .CO(cout[36]), .S(
        sumout[36]) );
endmodule


module csa51squ_71 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n4, n5, n6, n7, n8;

  NBUFFX2 U1 ( .INP(in1[6]), .Z(sumout[6]) );
  NBUFFX2 U2 ( .INP(in1[7]), .Z(sumout[7]) );
  NBUFFX2 U3 ( .INP(in3[37]), .Z(sumout[37]) );
  AND2X1 U4 ( .IN1(in2[8]), .IN2(in1[8]), .Q(cout[8]) );
  NOR2X0 U5 ( .IN1(in2[8]), .IN2(in1[8]), .QN(n4) );
  NOR2X0 U6 ( .IN1(n4), .IN2(cout[8]), .QN(sumout[8]) );
  AND2X1 U7 ( .IN1(in2[9]), .IN2(in1[9]), .Q(cout[9]) );
  NOR2X0 U8 ( .IN1(in2[9]), .IN2(in1[9]), .QN(n5) );
  NOR2X0 U9 ( .IN1(n5), .IN2(cout[9]), .QN(sumout[9]) );
  AND2X1 U10 ( .IN1(in2[34]), .IN2(in3[34]), .Q(cout[34]) );
  NOR2X0 U11 ( .IN1(in2[34]), .IN2(in3[34]), .QN(n6) );
  NOR2X0 U12 ( .IN1(n6), .IN2(cout[34]), .QN(sumout[34]) );
  INVX0 U13 ( .INP(in3[35]), .ZN(n7) );
  NOR2X0 U14 ( .IN1(in2[34]), .IN2(n7), .QN(cout[35]) );
  MUX21X1 U15 ( .IN1(n7), .IN2(in3[35]), .S(in2[34]), .Q(sumout[35]) );
  INVX0 U16 ( .INP(in1[32]), .ZN(n8) );
  FADDX1 U17 ( .A(in1[10]), .B(in2[10]), .CI(in3[10]), .CO(cout[10]), .S(
        sumout[10]) );
  FADDX1 U18 ( .A(in1[11]), .B(in2[11]), .CI(in3[11]), .CO(cout[11]), .S(
        sumout[11]) );
  FADDX1 U19 ( .A(in1[12]), .B(in2[12]), .CI(in3[12]), .CO(cout[12]), .S(
        sumout[12]) );
  FADDX1 U20 ( .A(in1[13]), .B(in2[13]), .CI(in3[13]), .CO(cout[13]), .S(
        sumout[13]) );
  FADDX1 U21 ( .A(in1[14]), .B(in2[14]), .CI(in3[14]), .CO(cout[14]), .S(
        sumout[14]) );
  FADDX1 U22 ( .A(in1[15]), .B(in2[15]), .CI(in3[15]), .CO(cout[15]), .S(
        sumout[15]) );
  FADDX1 U23 ( .A(in1[16]), .B(in2[16]), .CI(in3[16]), .CO(cout[16]), .S(
        sumout[16]) );
  FADDX1 U24 ( .A(in1[17]), .B(in2[17]), .CI(in3[17]), .CO(cout[17]), .S(
        sumout[17]) );
  FADDX1 U25 ( .A(in1[18]), .B(in2[18]), .CI(in3[18]), .CO(cout[18]), .S(
        sumout[18]) );
  FADDX1 U26 ( .A(in1[19]), .B(in2[19]), .CI(in3[19]), .CO(cout[19]), .S(
        sumout[19]) );
  FADDX1 U27 ( .A(in1[20]), .B(in2[20]), .CI(in3[20]), .CO(cout[20]), .S(
        sumout[20]) );
  FADDX1 U28 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U29 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U30 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U31 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U32 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U33 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U34 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U35 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U36 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U37 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U38 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U39 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
  FADDX1 U40 ( .A(in2[33]), .B(in3[33]), .CI(n8), .CO(cout[33]), .S(sumout[33]) );
endmodule


module csa51squ_72 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n2, n3, n4, n5;

  NBUFFX2 U1 ( .INP(in3[31]), .Z(sumout[31]) );
  AND2X1 U2 ( .IN1(in2[2]), .IN2(in1[2]), .Q(cout[2]) );
  AND2X1 U3 ( .IN1(in2[3]), .IN2(in1[3]), .Q(cout[3]) );
  NOR2X0 U4 ( .IN1(in2[3]), .IN2(in1[3]), .QN(n2) );
  NOR2X0 U5 ( .IN1(n2), .IN2(cout[3]), .QN(sumout[3]) );
  AND2X1 U6 ( .IN1(in2[28]), .IN2(in3[28]), .Q(cout[28]) );
  NOR2X0 U7 ( .IN1(in2[28]), .IN2(in3[28]), .QN(n3) );
  NOR2X0 U8 ( .IN1(n3), .IN2(cout[28]), .QN(sumout[28]) );
  INVX0 U9 ( .INP(in3[29]), .ZN(n4) );
  NOR2X0 U10 ( .IN1(in2[28]), .IN2(n4), .QN(cout[29]) );
  MUX21X1 U11 ( .IN1(n4), .IN2(in3[29]), .S(in2[28]), .Q(sumout[29]) );
  INVX0 U12 ( .INP(in1[26]), .ZN(n5) );
  FADDX1 U13 ( .A(in1[10]), .B(in2[10]), .CI(in3[10]), .CO(cout[10]), .S(
        sumout[10]) );
  FADDX1 U14 ( .A(in1[11]), .B(in2[11]), .CI(in3[11]), .CO(cout[11]), .S(
        sumout[11]) );
  FADDX1 U15 ( .A(in1[12]), .B(in2[12]), .CI(in3[12]), .CO(cout[12]), .S(
        sumout[12]) );
  FADDX1 U16 ( .A(in1[13]), .B(in2[13]), .CI(in3[13]), .CO(cout[13]), .S(
        sumout[13]) );
  FADDX1 U17 ( .A(in1[14]), .B(in2[14]), .CI(in3[14]), .CO(cout[14]), .S(
        sumout[14]) );
  FADDX1 U18 ( .A(in1[15]), .B(in2[15]), .CI(in3[15]), .CO(cout[15]), .S(
        sumout[15]) );
  FADDX1 U19 ( .A(in1[16]), .B(in2[16]), .CI(in3[16]), .CO(cout[16]), .S(
        sumout[16]) );
  FADDX1 U20 ( .A(in1[17]), .B(in2[17]), .CI(in3[17]), .CO(cout[17]), .S(
        sumout[17]) );
  FADDX1 U21 ( .A(in1[18]), .B(in2[18]), .CI(in3[18]), .CO(cout[18]), .S(
        sumout[18]) );
  FADDX1 U22 ( .A(in1[19]), .B(in2[19]), .CI(in3[19]), .CO(cout[19]), .S(
        sumout[19]) );
  FADDX1 U23 ( .A(in1[20]), .B(in2[20]), .CI(in3[20]), .CO(cout[20]), .S(
        sumout[20]) );
  FADDX1 U24 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U25 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U26 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U27 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U28 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U29 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U30 ( .A(in2[27]), .B(in3[27]), .CI(n5), .CO(cout[27]), .S(sumout[27]) );
  FADDX1 U31 ( .A(in1[4]), .B(in2[4]), .CI(in3[4]), .CO(cout[4]), .S(sumout[4]) );
  FADDX1 U32 ( .A(in1[5]), .B(in2[5]), .CI(in3[5]), .CO(cout[5]), .S(sumout[5]) );
  FADDX1 U33 ( .A(in1[6]), .B(in2[6]), .CI(in3[6]), .CO(cout[6]), .S(sumout[6]) );
  FADDX1 U34 ( .A(in1[7]), .B(in2[7]), .CI(in3[7]), .CO(cout[7]), .S(sumout[7]) );
  FADDX1 U35 ( .A(in1[8]), .B(in2[8]), .CI(in3[8]), .CO(cout[8]), .S(sumout[8]) );
  FADDX1 U36 ( .A(in1[9]), .B(in2[9]), .CI(in3[9]), .CO(cout[9]), .S(sumout[9]) );
endmodule


module booth27_66 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;


  NBUFFX2 U3 ( .INP(in2[22]), .Z(out1[22]) );
  NBUFFX2 U4 ( .INP(in2[21]), .Z(out1[21]) );
  NBUFFX2 U5 ( .INP(in2[20]), .Z(out1[20]) );
  NBUFFX2 U6 ( .INP(in2[0]), .Z(out1[0]) );
  NBUFFX2 U7 ( .INP(in2[19]), .Z(out1[19]) );
  NBUFFX2 U8 ( .INP(in2[18]), .Z(out1[18]) );
  NBUFFX2 U9 ( .INP(in2[4]), .Z(out1[4]) );
  NBUFFX2 U10 ( .INP(in2[3]), .Z(out1[3]) );
  NBUFFX2 U11 ( .INP(in2[2]), .Z(out1[2]) );
  NBUFFX2 U12 ( .INP(in2[1]), .Z(out1[1]) );
  NBUFFX2 U13 ( .INP(in2[6]), .Z(out1[6]) );
  NBUFFX2 U14 ( .INP(in2[5]), .Z(out1[5]) );
  NBUFFX2 U15 ( .INP(in2[9]), .Z(out1[9]) );
  NBUFFX2 U16 ( .INP(in2[8]), .Z(out1[8]) );
  NBUFFX2 U17 ( .INP(in2[7]), .Z(out1[7]) );
  NBUFFX2 U18 ( .INP(in2[13]), .Z(out1[13]) );
  NBUFFX2 U19 ( .INP(in2[12]), .Z(out1[12]) );
  NBUFFX2 U20 ( .INP(in2[11]), .Z(out1[11]) );
  NBUFFX2 U21 ( .INP(in2[10]), .Z(out1[10]) );
  NBUFFX2 U22 ( .INP(in2[17]), .Z(out1[17]) );
  NBUFFX2 U23 ( .INP(in2[16]), .Z(out1[16]) );
  NBUFFX2 U24 ( .INP(in2[15]), .Z(out1[15]) );
  NBUFFX2 U25 ( .INP(in2[14]), .Z(out1[14]) );
endmodule


module booth27_67 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76;

  NAND2X0 U3 ( .IN1(n1), .IN2(n2), .QN(n8) );
  NAND2X0 U4 ( .IN1(n71), .IN2(in2[0]), .QN(n15) );
  NAND2X0 U5 ( .IN1(n19), .IN2(in2[5]), .QN(n20) );
  NAND2X0 U6 ( .IN1(n25), .IN2(in2[7]), .QN(n26) );
  NAND2X0 U7 ( .IN1(n31), .IN2(in2[9]), .QN(n32) );
  NAND2X0 U8 ( .IN1(n37), .IN2(in2[11]), .QN(n38) );
  NAND2X0 U9 ( .IN1(n43), .IN2(in2[13]), .QN(n44) );
  NAND2X0 U10 ( .IN1(n46), .IN2(in2[14]), .QN(n47) );
  NAND2X0 U11 ( .IN1(n49), .IN2(in2[15]), .QN(n50) );
  NAND2X0 U12 ( .IN1(n52), .IN2(in2[16]), .QN(n53) );
  NAND2X0 U13 ( .IN1(n55), .IN2(in2[17]), .QN(n56) );
  NAND2X0 U14 ( .IN1(n7), .IN2(n15), .QN(out1[1]) );
  NAND2X0 U15 ( .IN1(n10), .IN2(n9), .QN(out1[2]) );
  NAND2X0 U16 ( .IN1(n58), .IN2(in2[18]), .QN(n59) );
  NAND2X0 U17 ( .IN1(n61), .IN2(in2[19]), .QN(n62) );
  NAND2X0 U18 ( .IN1(in1[1]), .IN2(in1[0]), .QN(out1[25]) );
  NOR2X0 U19 ( .IN1(in1[1]), .IN2(in1[0]), .QN(n71) );
  INVX0 U20 ( .INP(in2[0]), .ZN(n1) );
  INVX0 U21 ( .INP(in2[1]), .ZN(n2) );
  INVX0 U22 ( .INP(in2[3]), .ZN(n3) );
  INVX0 U23 ( .INP(in2[21]), .ZN(n4) );
  INVX0 U24 ( .INP(in2[22]), .ZN(n5) );
  INVX0 U25 ( .INP(in1[1]), .ZN(n6) );
  MUX21X1 U26 ( .IN1(in1[1]), .IN2(n6), .S(in1[0]), .Q(n74) );
  INVX0 U27 ( .INP(n74), .ZN(n76) );
  AO221X1 U28 ( .IN1(in2[0]), .IN2(in2[1]), .IN3(n1), .IN4(n2), .IN5(n76), .Q(
        n7) );
  MUX21X1 U29 ( .IN1(n2), .IN2(n8), .S(in2[2]), .Q(n12) );
  AO221X1 U30 ( .IN1(n12), .IN2(in2[2]), .IN3(n12), .IN4(n1), .IN5(n76), .Q(
        n10) );
  INVX0 U31 ( .INP(n71), .ZN(n13) );
  AO221X1 U32 ( .IN1(in2[0]), .IN2(in2[1]), .IN3(n1), .IN4(n2), .IN5(n13), .Q(
        n9) );
  NOR3X0 U33 ( .IN1(in2[0]), .IN2(in2[2]), .IN3(in2[1]), .QN(n11) );
  OR4X1 U34 ( .IN1(in2[3]), .IN2(in2[0]), .IN3(in2[2]), .IN4(in2[1]), .Q(n16)
         );
  OA21X1 U35 ( .IN1(n11), .IN2(n3), .IN3(n16), .Q(n18) );
  INVX0 U36 ( .INP(n18), .ZN(n14) );
  OAI222X1 U37 ( .IN1(n15), .IN2(in2[2]), .IN3(n14), .IN4(n76), .IN5(n13), 
        .IN6(n12), .QN(out1[3]) );
  OR2X1 U38 ( .IN1(in2[4]), .IN2(n16), .Q(n19) );
  NAND2X0 U39 ( .IN1(n16), .IN2(in2[4]), .QN(n17) );
  AND2X1 U40 ( .IN1(n19), .IN2(n17), .Q(n21) );
  AO22X1 U41 ( .IN1(n71), .IN2(n18), .IN3(n21), .IN4(n74), .Q(out1[4]) );
  OR2X1 U42 ( .IN1(in2[5]), .IN2(n19), .Q(n22) );
  AND2X1 U43 ( .IN1(n22), .IN2(n20), .Q(n24) );
  AO22X1 U44 ( .IN1(n71), .IN2(n21), .IN3(n24), .IN4(n74), .Q(out1[5]) );
  OR2X1 U45 ( .IN1(in2[6]), .IN2(n22), .Q(n25) );
  NAND2X0 U46 ( .IN1(n22), .IN2(in2[6]), .QN(n23) );
  AND2X1 U47 ( .IN1(n25), .IN2(n23), .Q(n27) );
  AO22X1 U48 ( .IN1(n71), .IN2(n24), .IN3(n27), .IN4(n74), .Q(out1[6]) );
  OR2X1 U49 ( .IN1(in2[7]), .IN2(n25), .Q(n28) );
  AND2X1 U50 ( .IN1(n28), .IN2(n26), .Q(n30) );
  AO22X1 U51 ( .IN1(n71), .IN2(n27), .IN3(n30), .IN4(n74), .Q(out1[7]) );
  OR2X1 U52 ( .IN1(in2[8]), .IN2(n28), .Q(n31) );
  NAND2X0 U53 ( .IN1(n28), .IN2(in2[8]), .QN(n29) );
  AND2X1 U54 ( .IN1(n31), .IN2(n29), .Q(n33) );
  AO22X1 U55 ( .IN1(n71), .IN2(n30), .IN3(n33), .IN4(n74), .Q(out1[8]) );
  OR2X1 U56 ( .IN1(in2[9]), .IN2(n31), .Q(n34) );
  AND2X1 U57 ( .IN1(n34), .IN2(n32), .Q(n36) );
  AO22X1 U58 ( .IN1(n71), .IN2(n33), .IN3(n36), .IN4(n74), .Q(out1[9]) );
  OR2X1 U59 ( .IN1(in2[10]), .IN2(n34), .Q(n37) );
  NAND2X0 U60 ( .IN1(n34), .IN2(in2[10]), .QN(n35) );
  AND2X1 U61 ( .IN1(n37), .IN2(n35), .Q(n39) );
  AO22X1 U62 ( .IN1(n71), .IN2(n36), .IN3(n39), .IN4(n74), .Q(out1[10]) );
  OR2X1 U63 ( .IN1(in2[11]), .IN2(n37), .Q(n40) );
  AND2X1 U64 ( .IN1(n40), .IN2(n38), .Q(n42) );
  AO22X1 U65 ( .IN1(n71), .IN2(n39), .IN3(n42), .IN4(n74), .Q(out1[11]) );
  OR2X1 U66 ( .IN1(in2[12]), .IN2(n40), .Q(n43) );
  NAND2X0 U67 ( .IN1(n40), .IN2(in2[12]), .QN(n41) );
  AND2X1 U68 ( .IN1(n43), .IN2(n41), .Q(n45) );
  AO22X1 U69 ( .IN1(n71), .IN2(n42), .IN3(n45), .IN4(n74), .Q(out1[12]) );
  OR2X1 U70 ( .IN1(in2[13]), .IN2(n43), .Q(n46) );
  AND2X1 U71 ( .IN1(n46), .IN2(n44), .Q(n48) );
  AO22X1 U72 ( .IN1(n71), .IN2(n45), .IN3(n48), .IN4(n74), .Q(out1[13]) );
  OR2X1 U73 ( .IN1(in2[14]), .IN2(n46), .Q(n49) );
  AND2X1 U74 ( .IN1(n49), .IN2(n47), .Q(n51) );
  AO22X1 U75 ( .IN1(n71), .IN2(n48), .IN3(n51), .IN4(n74), .Q(out1[14]) );
  OR2X1 U76 ( .IN1(in2[15]), .IN2(n49), .Q(n52) );
  AND2X1 U77 ( .IN1(n52), .IN2(n50), .Q(n54) );
  AO22X1 U78 ( .IN1(n71), .IN2(n51), .IN3(n54), .IN4(n74), .Q(out1[15]) );
  OR2X1 U79 ( .IN1(in2[16]), .IN2(n52), .Q(n55) );
  AND2X1 U80 ( .IN1(n55), .IN2(n53), .Q(n57) );
  AO22X1 U81 ( .IN1(n71), .IN2(n54), .IN3(n57), .IN4(n74), .Q(out1[16]) );
  OR2X1 U82 ( .IN1(in2[17]), .IN2(n55), .Q(n58) );
  AND2X1 U83 ( .IN1(n58), .IN2(n56), .Q(n60) );
  AO22X1 U84 ( .IN1(n71), .IN2(n57), .IN3(n60), .IN4(n74), .Q(out1[17]) );
  OR2X1 U85 ( .IN1(in2[18]), .IN2(n58), .Q(n61) );
  AND2X1 U86 ( .IN1(n61), .IN2(n59), .Q(n63) );
  AO22X1 U87 ( .IN1(n71), .IN2(n60), .IN3(n63), .IN4(n74), .Q(out1[18]) );
  OR2X1 U88 ( .IN1(in2[19]), .IN2(n61), .Q(n64) );
  AND2X1 U89 ( .IN1(n64), .IN2(n62), .Q(n65) );
  AO22X1 U90 ( .IN1(n71), .IN2(n63), .IN3(n65), .IN4(n74), .Q(out1[19]) );
  NOR2X0 U91 ( .IN1(in2[20]), .IN2(n64), .QN(n72) );
  AOI21X1 U92 ( .IN1(in2[20]), .IN2(n64), .IN3(n72), .QN(n66) );
  AO22X1 U93 ( .IN1(n71), .IN2(n65), .IN3(n66), .IN4(n74), .Q(out1[20]) );
  MUX21X1 U94 ( .IN1(n4), .IN2(in2[21]), .S(n72), .Q(n69) );
  AO22X1 U95 ( .IN1(n71), .IN2(n66), .IN3(n69), .IN4(n74), .Q(out1[21]) );
  INVX0 U96 ( .INP(n72), .ZN(n67) );
  NOR2X0 U97 ( .IN1(in2[21]), .IN2(n67), .QN(n70) );
  MUX21X1 U98 ( .IN1(n5), .IN2(in2[22]), .S(n70), .Q(n68) );
  AO22X1 U99 ( .IN1(n71), .IN2(n69), .IN3(n68), .IN4(n74), .Q(out1[22]) );
  MUX21X1 U100 ( .IN1(n71), .IN2(n74), .S(n70), .Q(n73) );
  AND3X1 U101 ( .IN1(n72), .IN2(n71), .IN3(n4), .Q(n75) );
  MUX21X1 U102 ( .IN1(n73), .IN2(n75), .S(in2[22]), .Q(out1[23]) );
  AO21X1 U103 ( .IN1(n75), .IN2(n5), .IN3(n74), .Q(out1[24]) );
  NOR2X0 U104 ( .IN1(n76), .IN2(n1), .QN(out1[0]) );
endmodule


module booth27_68 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n25), .IN2(n6), .QN(n30) );
  NAND2X0 U4 ( .IN1(n33), .IN2(n7), .QN(n37) );
  NAND2X0 U5 ( .IN1(n41), .IN2(n8), .QN(n45) );
  NAND2X0 U6 ( .IN1(n49), .IN2(n9), .QN(n53) );
  NAND2X0 U7 ( .IN1(n57), .IN2(n10), .QN(n61) );
  NAND2X0 U8 ( .IN1(n65), .IN2(n11), .QN(n77) );
  NAND2X0 U9 ( .IN1(n81), .IN2(n13), .QN(n89) );
  NAND2X0 U10 ( .IN1(n93), .IN2(n15), .QN(n101) );
  NAND2X0 U11 ( .IN1(n105), .IN2(n17), .QN(n114) );
  NAND2X0 U12 ( .IN1(n27), .IN2(n132), .QN(n4) );
  NAND2X0 U13 ( .IN1(in1[2]), .IN2(n77), .QN(n71) );
  NAND2X0 U14 ( .IN1(n70), .IN2(n132), .QN(n74) );
  NAND2X0 U15 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U16 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U17 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U18 ( .IN1(n118), .IN2(n19), .QN(n125) );
  NAND2X0 U19 ( .IN1(n141), .IN2(n130), .QN(n24) );
  NAND2X0 U20 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NAND2X0 U21 ( .IN1(n32), .IN2(n31), .QN(out1[3]) );
  NAND2X0 U22 ( .IN1(n36), .IN2(n35), .QN(out1[4]) );
  NAND2X0 U23 ( .IN1(n40), .IN2(n39), .QN(out1[5]) );
  NAND2X0 U24 ( .IN1(n44), .IN2(n43), .QN(out1[6]) );
  NAND2X0 U25 ( .IN1(n48), .IN2(n47), .QN(out1[7]) );
  NAND2X0 U26 ( .IN1(n52), .IN2(n51), .QN(out1[8]) );
  NAND2X0 U27 ( .IN1(n56), .IN2(n55), .QN(out1[9]) );
  NAND2X0 U28 ( .IN1(n60), .IN2(n59), .QN(out1[10]) );
  NAND2X0 U29 ( .IN1(n64), .IN2(n63), .QN(out1[11]) );
  NAND2X0 U30 ( .IN1(n69), .IN2(n68), .QN(out1[12]) );
  NAND2X0 U31 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U32 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U33 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U34 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U35 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U36 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U37 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U38 ( .IN1(n23), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U39 ( .IN1(in1[2]), .IN2(n22), .QN(n23) );
  NOR2X0 U40 ( .IN1(n28), .IN2(n26), .QN(n3) );
  NOR2X0 U41 ( .IN1(n142), .IN2(n21), .QN(n1) );
  NOR2X0 U42 ( .IN1(n142), .IN2(n111), .QN(n138) );
  INVX0 U43 ( .INP(n130), .ZN(n137) );
  INVX0 U44 ( .INP(n132), .ZN(n141) );
  NOR3X0 U45 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  NAND3X0 U46 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  MUX21X1 U47 ( .IN1(n22), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  INVX0 U48 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U49 ( .INP(in2[2]), .ZN(n6) );
  INVX0 U50 ( .INP(in2[4]), .ZN(n7) );
  INVX0 U51 ( .INP(in2[6]), .ZN(n8) );
  INVX0 U52 ( .INP(in2[8]), .ZN(n9) );
  INVX0 U53 ( .INP(in2[10]), .ZN(n10) );
  INVX0 U54 ( .INP(in2[12]), .ZN(n11) );
  INVX0 U55 ( .INP(in2[13]), .ZN(n12) );
  INVX0 U56 ( .INP(in2[14]), .ZN(n13) );
  INVX0 U57 ( .INP(in2[15]), .ZN(n14) );
  INVX0 U58 ( .INP(in2[16]), .ZN(n15) );
  INVX0 U59 ( .INP(in2[17]), .ZN(n16) );
  INVX0 U60 ( .INP(in2[18]), .ZN(n17) );
  INVX0 U61 ( .INP(in2[19]), .ZN(n18) );
  INVX0 U62 ( .INP(in2[20]), .ZN(n19) );
  INVX0 U63 ( .INP(in2[21]), .ZN(n20) );
  INVX0 U64 ( .INP(in2[22]), .ZN(n21) );
  INVX0 U65 ( .INP(in1[1]), .ZN(n22) );
  INVX0 U66 ( .INP(in1[2]), .ZN(n111) );
  INVX0 U67 ( .INP(n138), .ZN(n140) );
  NOR2X0 U68 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n25) );
  AOI21X1 U69 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n25), .QN(n27) );
  NOR2X0 U70 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U71 ( .IN1(n24), .IN2(in2[0]), .IN3(n138), .IN4(n27), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U72 ( .INP(n133), .ZN(n67) );
  NOR2X0 U73 ( .IN1(n67), .IN2(n6), .QN(n28) );
  OA21X1 U74 ( .IN1(n25), .IN2(n6), .IN3(n30), .Q(n29) );
  AO22X1 U75 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n29), .Q(n26) );
  AOI22X1 U76 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n29), .QN(n32) );
  NOR2X0 U77 ( .IN1(in2[3]), .IN2(n30), .QN(n33) );
  AO21X1 U78 ( .IN1(in2[3]), .IN2(n30), .IN3(n33), .Q(n34) );
  OA22X1 U79 ( .IN1(n6), .IN2(n130), .IN3(n140), .IN4(n34), .Q(n31) );
  OA21X1 U80 ( .IN1(n33), .IN2(n7), .IN3(n37), .Q(n38) );
  AOI22X1 U81 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n38), .QN(n36) );
  OA22X1 U82 ( .IN1(n67), .IN2(n7), .IN3(n141), .IN4(n34), .Q(n35) );
  NOR2X0 U83 ( .IN1(in2[5]), .IN2(n37), .QN(n41) );
  AO21X1 U84 ( .IN1(in2[5]), .IN2(n37), .IN3(n41), .Q(n42) );
  OA22X1 U85 ( .IN1(n7), .IN2(n130), .IN3(n140), .IN4(n42), .Q(n40) );
  AOI22X1 U86 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n38), .QN(n39) );
  OA21X1 U87 ( .IN1(n41), .IN2(n8), .IN3(n45), .Q(n46) );
  AOI22X1 U88 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n46), .QN(n44) );
  OA22X1 U89 ( .IN1(n67), .IN2(n8), .IN3(n141), .IN4(n42), .Q(n43) );
  NOR2X0 U90 ( .IN1(in2[7]), .IN2(n45), .QN(n49) );
  AO21X1 U91 ( .IN1(in2[7]), .IN2(n45), .IN3(n49), .Q(n50) );
  OA22X1 U92 ( .IN1(n8), .IN2(n130), .IN3(n140), .IN4(n50), .Q(n48) );
  AOI22X1 U93 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n46), .QN(n47) );
  OA21X1 U94 ( .IN1(n49), .IN2(n9), .IN3(n53), .Q(n54) );
  AOI22X1 U95 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n54), .QN(n52) );
  OA22X1 U96 ( .IN1(n67), .IN2(n9), .IN3(n141), .IN4(n50), .Q(n51) );
  NOR2X0 U97 ( .IN1(in2[9]), .IN2(n53), .QN(n57) );
  AO21X1 U98 ( .IN1(in2[9]), .IN2(n53), .IN3(n57), .Q(n58) );
  OA22X1 U99 ( .IN1(n9), .IN2(n130), .IN3(n140), .IN4(n58), .Q(n56) );
  AOI22X1 U100 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n54), .QN(n55) );
  OA21X1 U101 ( .IN1(n57), .IN2(n10), .IN3(n61), .Q(n62) );
  AOI22X1 U102 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n62), .QN(n60) );
  OA22X1 U103 ( .IN1(n67), .IN2(n10), .IN3(n141), .IN4(n58), .Q(n59) );
  NOR2X0 U104 ( .IN1(in2[11]), .IN2(n61), .QN(n65) );
  AO21X1 U105 ( .IN1(in2[11]), .IN2(n61), .IN3(n65), .Q(n66) );
  OA22X1 U106 ( .IN1(n10), .IN2(n130), .IN3(n140), .IN4(n66), .Q(n64) );
  AOI22X1 U107 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n62), .QN(n63) );
  OA21X1 U108 ( .IN1(n65), .IN2(n11), .IN3(n77), .Q(n70) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n70), .QN(n69) );
  OA22X1 U110 ( .IN1(n67), .IN2(n11), .IN3(n141), .IN4(n66), .Q(n68) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n12), .S(n71), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n11), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n13), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n12), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n12), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n14), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n13), .IN4(n85), .IN5(n84), 
        .Q(out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n15), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n14), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n14), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n16), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n15), .IN4(n97), .IN5(n96), 
        .Q(out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n17), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n16), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n16), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n18), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n17), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n19), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n18), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n18), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n20), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n19), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n21), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n20), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n20), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n21), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_69 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n33), .IN2(n7), .QN(n37) );
  NAND2X0 U4 ( .IN1(n41), .IN2(n8), .QN(n45) );
  NAND2X0 U5 ( .IN1(n49), .IN2(n9), .QN(n53) );
  NAND2X0 U6 ( .IN1(n57), .IN2(n10), .QN(n61) );
  NAND2X0 U7 ( .IN1(n25), .IN2(n6), .QN(n30) );
  NAND2X0 U8 ( .IN1(n65), .IN2(n11), .QN(n77) );
  NAND2X0 U9 ( .IN1(n81), .IN2(n13), .QN(n89) );
  NAND2X0 U10 ( .IN1(n93), .IN2(n15), .QN(n101) );
  NAND2X0 U11 ( .IN1(n105), .IN2(n17), .QN(n114) );
  NAND2X0 U12 ( .IN1(n118), .IN2(n19), .QN(n125) );
  NAND2X0 U13 ( .IN1(in1[2]), .IN2(n77), .QN(n71) );
  NAND2X0 U14 ( .IN1(n70), .IN2(n132), .QN(n74) );
  NAND2X0 U15 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U16 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U17 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U18 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U19 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U20 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U21 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U22 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NAND2X0 U23 ( .IN1(n27), .IN2(n132), .QN(n4) );
  NAND2X0 U24 ( .IN1(n32), .IN2(n31), .QN(out1[3]) );
  NAND2X0 U25 ( .IN1(n36), .IN2(n35), .QN(out1[4]) );
  NAND2X0 U26 ( .IN1(n40), .IN2(n39), .QN(out1[5]) );
  NAND2X0 U27 ( .IN1(n44), .IN2(n43), .QN(out1[6]) );
  NAND2X0 U28 ( .IN1(n48), .IN2(n47), .QN(out1[7]) );
  NAND2X0 U29 ( .IN1(n52), .IN2(n51), .QN(out1[8]) );
  NAND2X0 U30 ( .IN1(n56), .IN2(n55), .QN(out1[9]) );
  NAND2X0 U31 ( .IN1(n60), .IN2(n59), .QN(out1[10]) );
  NAND2X0 U32 ( .IN1(n64), .IN2(n63), .QN(out1[11]) );
  NAND2X0 U33 ( .IN1(n69), .IN2(n68), .QN(out1[12]) );
  NAND2X0 U34 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U35 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U36 ( .IN1(n141), .IN2(n130), .QN(n24) );
  NAND2X0 U37 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U38 ( .IN1(n23), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U39 ( .IN1(in1[2]), .IN2(n22), .QN(n23) );
  NOR2X0 U40 ( .IN1(n28), .IN2(n26), .QN(n3) );
  NOR2X0 U41 ( .IN1(n142), .IN2(n111), .QN(n138) );
  NOR2X0 U42 ( .IN1(n142), .IN2(n21), .QN(n1) );
  INVX0 U43 ( .INP(n130), .ZN(n137) );
  INVX0 U44 ( .INP(n132), .ZN(n141) );
  NOR3X0 U45 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  NAND3X0 U46 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  MUX21X1 U47 ( .IN1(n22), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  INVX0 U48 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U49 ( .INP(in2[2]), .ZN(n6) );
  INVX0 U50 ( .INP(in2[4]), .ZN(n7) );
  INVX0 U51 ( .INP(in2[6]), .ZN(n8) );
  INVX0 U52 ( .INP(in2[8]), .ZN(n9) );
  INVX0 U53 ( .INP(in2[10]), .ZN(n10) );
  INVX0 U54 ( .INP(in2[12]), .ZN(n11) );
  INVX0 U55 ( .INP(in2[13]), .ZN(n12) );
  INVX0 U56 ( .INP(in2[14]), .ZN(n13) );
  INVX0 U57 ( .INP(in2[15]), .ZN(n14) );
  INVX0 U58 ( .INP(in2[16]), .ZN(n15) );
  INVX0 U59 ( .INP(in2[17]), .ZN(n16) );
  INVX0 U60 ( .INP(in2[18]), .ZN(n17) );
  INVX0 U61 ( .INP(in2[19]), .ZN(n18) );
  INVX0 U62 ( .INP(in2[20]), .ZN(n19) );
  INVX0 U63 ( .INP(in2[21]), .ZN(n20) );
  INVX0 U64 ( .INP(in2[22]), .ZN(n21) );
  INVX0 U65 ( .INP(in1[1]), .ZN(n22) );
  INVX0 U66 ( .INP(in1[2]), .ZN(n111) );
  INVX0 U67 ( .INP(n138), .ZN(n140) );
  NOR2X0 U68 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n25) );
  AOI21X1 U69 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n25), .QN(n27) );
  NOR2X0 U70 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U71 ( .IN1(n24), .IN2(in2[0]), .IN3(n138), .IN4(n27), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U72 ( .INP(n133), .ZN(n67) );
  NOR2X0 U73 ( .IN1(n67), .IN2(n6), .QN(n28) );
  OA21X1 U74 ( .IN1(n25), .IN2(n6), .IN3(n30), .Q(n29) );
  AO22X1 U75 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n29), .Q(n26) );
  AOI22X1 U76 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n29), .QN(n32) );
  NOR2X0 U77 ( .IN1(in2[3]), .IN2(n30), .QN(n33) );
  AO21X1 U78 ( .IN1(in2[3]), .IN2(n30), .IN3(n33), .Q(n34) );
  OA22X1 U79 ( .IN1(n6), .IN2(n130), .IN3(n140), .IN4(n34), .Q(n31) );
  OA21X1 U80 ( .IN1(n33), .IN2(n7), .IN3(n37), .Q(n38) );
  AOI22X1 U81 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n38), .QN(n36) );
  OA22X1 U82 ( .IN1(n67), .IN2(n7), .IN3(n141), .IN4(n34), .Q(n35) );
  NOR2X0 U83 ( .IN1(in2[5]), .IN2(n37), .QN(n41) );
  AO21X1 U84 ( .IN1(in2[5]), .IN2(n37), .IN3(n41), .Q(n42) );
  OA22X1 U85 ( .IN1(n7), .IN2(n130), .IN3(n140), .IN4(n42), .Q(n40) );
  AOI22X1 U86 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n38), .QN(n39) );
  OA21X1 U87 ( .IN1(n41), .IN2(n8), .IN3(n45), .Q(n46) );
  AOI22X1 U88 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n46), .QN(n44) );
  OA22X1 U89 ( .IN1(n67), .IN2(n8), .IN3(n141), .IN4(n42), .Q(n43) );
  NOR2X0 U90 ( .IN1(in2[7]), .IN2(n45), .QN(n49) );
  AO21X1 U91 ( .IN1(in2[7]), .IN2(n45), .IN3(n49), .Q(n50) );
  OA22X1 U92 ( .IN1(n8), .IN2(n130), .IN3(n140), .IN4(n50), .Q(n48) );
  AOI22X1 U93 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n46), .QN(n47) );
  OA21X1 U94 ( .IN1(n49), .IN2(n9), .IN3(n53), .Q(n54) );
  AOI22X1 U95 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n54), .QN(n52) );
  OA22X1 U96 ( .IN1(n67), .IN2(n9), .IN3(n141), .IN4(n50), .Q(n51) );
  NOR2X0 U97 ( .IN1(in2[9]), .IN2(n53), .QN(n57) );
  AO21X1 U98 ( .IN1(in2[9]), .IN2(n53), .IN3(n57), .Q(n58) );
  OA22X1 U99 ( .IN1(n9), .IN2(n130), .IN3(n140), .IN4(n58), .Q(n56) );
  AOI22X1 U100 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n54), .QN(n55) );
  OA21X1 U101 ( .IN1(n57), .IN2(n10), .IN3(n61), .Q(n62) );
  AOI22X1 U102 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n62), .QN(n60) );
  OA22X1 U103 ( .IN1(n67), .IN2(n10), .IN3(n141), .IN4(n58), .Q(n59) );
  NOR2X0 U104 ( .IN1(in2[11]), .IN2(n61), .QN(n65) );
  AO21X1 U105 ( .IN1(in2[11]), .IN2(n61), .IN3(n65), .Q(n66) );
  OA22X1 U106 ( .IN1(n10), .IN2(n130), .IN3(n140), .IN4(n66), .Q(n64) );
  AOI22X1 U107 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n62), .QN(n63) );
  OA21X1 U108 ( .IN1(n65), .IN2(n11), .IN3(n77), .Q(n70) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n70), .QN(n69) );
  OA22X1 U110 ( .IN1(n67), .IN2(n11), .IN3(n141), .IN4(n66), .Q(n68) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n12), .S(n71), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n11), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n13), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n12), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n12), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n14), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n13), .IN4(n85), .IN5(n84), 
        .Q(out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n15), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n14), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n14), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n16), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n15), .IN4(n97), .IN5(n96), 
        .Q(out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n17), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n16), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n16), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n18), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n17), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n19), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n18), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n18), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n20), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n19), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n21), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n20), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n20), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n21), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_70 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n41), .IN2(n8), .QN(n45) );
  NAND2X0 U4 ( .IN1(n49), .IN2(n9), .QN(n53) );
  NAND2X0 U5 ( .IN1(n57), .IN2(n10), .QN(n61) );
  NAND2X0 U6 ( .IN1(n33), .IN2(n7), .QN(n37) );
  NAND2X0 U7 ( .IN1(n25), .IN2(n6), .QN(n30) );
  NAND2X0 U8 ( .IN1(n65), .IN2(n11), .QN(n77) );
  NAND2X0 U9 ( .IN1(n81), .IN2(n13), .QN(n89) );
  NAND2X0 U10 ( .IN1(n93), .IN2(n15), .QN(n101) );
  NAND2X0 U11 ( .IN1(in1[2]), .IN2(n77), .QN(n71) );
  NAND2X0 U12 ( .IN1(n70), .IN2(n132), .QN(n74) );
  NAND2X0 U13 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U14 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U15 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U16 ( .IN1(n118), .IN2(n19), .QN(n125) );
  NAND2X0 U17 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U18 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U19 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U20 ( .IN1(n27), .IN2(n132), .QN(n4) );
  NAND2X0 U21 ( .IN1(n141), .IN2(n130), .QN(n24) );
  NAND2X0 U22 ( .IN1(n40), .IN2(n39), .QN(out1[5]) );
  NAND2X0 U23 ( .IN1(n44), .IN2(n43), .QN(out1[6]) );
  NAND2X0 U24 ( .IN1(n48), .IN2(n47), .QN(out1[7]) );
  NAND2X0 U25 ( .IN1(n52), .IN2(n51), .QN(out1[8]) );
  NAND2X0 U26 ( .IN1(n56), .IN2(n55), .QN(out1[9]) );
  NAND2X0 U27 ( .IN1(n60), .IN2(n59), .QN(out1[10]) );
  NAND2X0 U28 ( .IN1(n64), .IN2(n63), .QN(out1[11]) );
  NAND2X0 U29 ( .IN1(n69), .IN2(n68), .QN(out1[12]) );
  NAND2X0 U30 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U31 ( .IN1(n105), .IN2(n17), .QN(n114) );
  NAND2X0 U32 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U33 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U34 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U35 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NAND2X0 U36 ( .IN1(n32), .IN2(n31), .QN(out1[3]) );
  NAND2X0 U37 ( .IN1(n36), .IN2(n35), .QN(out1[4]) );
  NAND2X0 U38 ( .IN1(n23), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U39 ( .IN1(in1[2]), .IN2(n22), .QN(n23) );
  INVX0 U40 ( .INP(in1[2]), .ZN(n111) );
  NOR2X0 U41 ( .IN1(n28), .IN2(n26), .QN(n3) );
  NOR2X0 U42 ( .IN1(n142), .IN2(n21), .QN(n1) );
  INVX0 U43 ( .INP(n132), .ZN(n141) );
  INVX0 U44 ( .INP(n130), .ZN(n137) );
  NOR2X0 U45 ( .IN1(n142), .IN2(n111), .QN(n138) );
  MUX21X1 U46 ( .IN1(n22), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  NAND3X0 U47 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  NOR3X0 U48 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  INVX0 U49 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U50 ( .INP(in2[2]), .ZN(n6) );
  INVX0 U51 ( .INP(in2[4]), .ZN(n7) );
  INVX0 U52 ( .INP(in2[6]), .ZN(n8) );
  INVX0 U53 ( .INP(in2[8]), .ZN(n9) );
  INVX0 U54 ( .INP(in2[10]), .ZN(n10) );
  INVX0 U55 ( .INP(in2[12]), .ZN(n11) );
  INVX0 U56 ( .INP(in2[13]), .ZN(n12) );
  INVX0 U57 ( .INP(in2[14]), .ZN(n13) );
  INVX0 U58 ( .INP(in2[15]), .ZN(n14) );
  INVX0 U59 ( .INP(in2[16]), .ZN(n15) );
  INVX0 U60 ( .INP(in2[17]), .ZN(n16) );
  INVX0 U61 ( .INP(in2[18]), .ZN(n17) );
  INVX0 U62 ( .INP(in2[19]), .ZN(n18) );
  INVX0 U63 ( .INP(in2[20]), .ZN(n19) );
  INVX0 U64 ( .INP(in2[21]), .ZN(n20) );
  INVX0 U65 ( .INP(in2[22]), .ZN(n21) );
  INVX0 U66 ( .INP(in1[1]), .ZN(n22) );
  INVX0 U67 ( .INP(n138), .ZN(n140) );
  NOR2X0 U68 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n25) );
  AOI21X1 U69 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n25), .QN(n27) );
  NOR2X0 U70 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U71 ( .IN1(n24), .IN2(in2[0]), .IN3(n138), .IN4(n27), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U72 ( .INP(n133), .ZN(n67) );
  NOR2X0 U73 ( .IN1(n67), .IN2(n6), .QN(n28) );
  OA21X1 U74 ( .IN1(n25), .IN2(n6), .IN3(n30), .Q(n29) );
  AO22X1 U75 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n29), .Q(n26) );
  AOI22X1 U76 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n29), .QN(n32) );
  NOR2X0 U77 ( .IN1(in2[3]), .IN2(n30), .QN(n33) );
  AO21X1 U78 ( .IN1(in2[3]), .IN2(n30), .IN3(n33), .Q(n34) );
  OA22X1 U79 ( .IN1(n6), .IN2(n130), .IN3(n140), .IN4(n34), .Q(n31) );
  OA21X1 U80 ( .IN1(n33), .IN2(n7), .IN3(n37), .Q(n38) );
  AOI22X1 U81 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n38), .QN(n36) );
  OA22X1 U82 ( .IN1(n67), .IN2(n7), .IN3(n141), .IN4(n34), .Q(n35) );
  NOR2X0 U83 ( .IN1(in2[5]), .IN2(n37), .QN(n41) );
  AO21X1 U84 ( .IN1(in2[5]), .IN2(n37), .IN3(n41), .Q(n42) );
  OA22X1 U85 ( .IN1(n7), .IN2(n130), .IN3(n140), .IN4(n42), .Q(n40) );
  AOI22X1 U86 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n38), .QN(n39) );
  OA21X1 U87 ( .IN1(n41), .IN2(n8), .IN3(n45), .Q(n46) );
  AOI22X1 U88 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n46), .QN(n44) );
  OA22X1 U89 ( .IN1(n67), .IN2(n8), .IN3(n141), .IN4(n42), .Q(n43) );
  NOR2X0 U90 ( .IN1(in2[7]), .IN2(n45), .QN(n49) );
  AO21X1 U91 ( .IN1(in2[7]), .IN2(n45), .IN3(n49), .Q(n50) );
  OA22X1 U92 ( .IN1(n8), .IN2(n130), .IN3(n140), .IN4(n50), .Q(n48) );
  AOI22X1 U93 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n46), .QN(n47) );
  OA21X1 U94 ( .IN1(n49), .IN2(n9), .IN3(n53), .Q(n54) );
  AOI22X1 U95 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n54), .QN(n52) );
  OA22X1 U96 ( .IN1(n67), .IN2(n9), .IN3(n141), .IN4(n50), .Q(n51) );
  NOR2X0 U97 ( .IN1(in2[9]), .IN2(n53), .QN(n57) );
  AO21X1 U98 ( .IN1(in2[9]), .IN2(n53), .IN3(n57), .Q(n58) );
  OA22X1 U99 ( .IN1(n9), .IN2(n130), .IN3(n140), .IN4(n58), .Q(n56) );
  AOI22X1 U100 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n54), .QN(n55) );
  OA21X1 U101 ( .IN1(n57), .IN2(n10), .IN3(n61), .Q(n62) );
  AOI22X1 U102 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n62), .QN(n60) );
  OA22X1 U103 ( .IN1(n67), .IN2(n10), .IN3(n141), .IN4(n58), .Q(n59) );
  NOR2X0 U104 ( .IN1(in2[11]), .IN2(n61), .QN(n65) );
  AO21X1 U105 ( .IN1(in2[11]), .IN2(n61), .IN3(n65), .Q(n66) );
  OA22X1 U106 ( .IN1(n10), .IN2(n130), .IN3(n140), .IN4(n66), .Q(n64) );
  AOI22X1 U107 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n62), .QN(n63) );
  OA21X1 U108 ( .IN1(n65), .IN2(n11), .IN3(n77), .Q(n70) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n70), .QN(n69) );
  OA22X1 U110 ( .IN1(n67), .IN2(n11), .IN3(n141), .IN4(n66), .Q(n68) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n12), .S(n71), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n11), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n13), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n12), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n12), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n14), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n13), .IN4(n85), .IN5(n84), 
        .Q(out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n15), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n14), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n14), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n16), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n15), .IN4(n97), .IN5(n96), 
        .Q(out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n17), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n16), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n16), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n18), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n17), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n19), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n18), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n18), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n20), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n19), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n21), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n20), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n20), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n21), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_71 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90;

  NAND2X0 U3 ( .IN1(n31), .IN2(n6), .QN(n33) );
  NAND2X0 U4 ( .IN1(n35), .IN2(n7), .QN(n37) );
  NAND2X0 U5 ( .IN1(n39), .IN2(n8), .QN(n44) );
  NAND2X0 U6 ( .IN1(n23), .IN2(n4), .QN(n25) );
  NAND2X0 U7 ( .IN1(n27), .IN2(n5), .QN(n29) );
  NAND2X0 U8 ( .IN1(in1[2]), .IN2(n44), .QN(n41) );
  NAND2X0 U9 ( .IN1(n49), .IN2(n10), .QN(n52) );
  NAND2X0 U10 ( .IN1(in1[2]), .IN2(n52), .QN(n48) );
  NAND2X0 U11 ( .IN1(n57), .IN2(n12), .QN(n60) );
  NAND2X0 U12 ( .IN1(in1[2]), .IN2(n60), .QN(n56) );
  NAND2X0 U13 ( .IN1(n65), .IN2(n14), .QN(n68) );
  NAND2X0 U14 ( .IN1(in1[2]), .IN2(n68), .QN(n64) );
  NAND2X0 U15 ( .IN1(n75), .IN2(n16), .QN(n79) );
  NAND2X0 U16 ( .IN1(n72), .IN2(in1[2]), .QN(n83) );
  NAND2X0 U17 ( .IN1(in1[2]), .IN2(n79), .QN(n74) );
  NAND2X0 U18 ( .IN1(in2[21]), .IN2(n79), .QN(n80) );
  INVX0 U19 ( .INP(n83), .ZN(n86) );
  NOR2X0 U20 ( .IN1(n72), .IN2(n69), .QN(n89) );
  NOR2X0 U21 ( .IN1(in1[2]), .IN2(n72), .QN(n87) );
  NBUFFX2 U22 ( .INP(in1[2]), .Z(out1[26]) );
  NBUFFX2 U23 ( .INP(in1[2]), .Z(out1[25]) );
  INVX0 U24 ( .INP(in2[2]), .ZN(n3) );
  INVX0 U25 ( .INP(in2[4]), .ZN(n4) );
  INVX0 U26 ( .INP(in2[6]), .ZN(n5) );
  INVX0 U27 ( .INP(in2[8]), .ZN(n6) );
  INVX0 U28 ( .INP(in2[10]), .ZN(n7) );
  INVX0 U29 ( .INP(in2[12]), .ZN(n8) );
  INVX0 U30 ( .INP(in2[13]), .ZN(n9) );
  INVX0 U31 ( .INP(in2[14]), .ZN(n10) );
  INVX0 U32 ( .INP(in2[15]), .ZN(n11) );
  INVX0 U33 ( .INP(in2[16]), .ZN(n12) );
  INVX0 U34 ( .INP(in2[17]), .ZN(n13) );
  INVX0 U35 ( .INP(in2[18]), .ZN(n14) );
  INVX0 U36 ( .INP(in2[19]), .ZN(n15) );
  INVX0 U37 ( .INP(in2[20]), .ZN(n16) );
  INVX0 U38 ( .INP(in2[21]), .ZN(n17) );
  INVX0 U39 ( .INP(in2[22]), .ZN(n18) );
  INVX0 U40 ( .INP(in1[1]), .ZN(n72) );
  INVX0 U41 ( .INP(in1[2]), .ZN(n69) );
  NOR2X0 U42 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n19) );
  AOI21X1 U43 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n19), .QN(n20) );
  AO222X1 U44 ( .IN1(in2[0]), .IN2(n86), .IN3(in2[1]), .IN4(n87), .IN5(n89), 
        .IN6(n20), .Q(out1[1]) );
  OR3X1 U45 ( .IN1(in2[2]), .IN2(in2[0]), .IN3(in2[1]), .Q(n21) );
  OA21X1 U46 ( .IN1(n19), .IN2(n3), .IN3(n21), .Q(n22) );
  AO222X1 U47 ( .IN1(in2[2]), .IN2(n87), .IN3(n86), .IN4(n20), .IN5(n22), 
        .IN6(n89), .Q(out1[2]) );
  NOR2X0 U48 ( .IN1(in2[3]), .IN2(n21), .QN(n23) );
  AOI21X1 U49 ( .IN1(in2[3]), .IN2(n21), .IN3(n23), .QN(n24) );
  AO222X1 U50 ( .IN1(in2[3]), .IN2(n87), .IN3(n86), .IN4(n22), .IN5(n24), 
        .IN6(n89), .Q(out1[3]) );
  OA21X1 U51 ( .IN1(n23), .IN2(n4), .IN3(n25), .Q(n26) );
  AO222X1 U52 ( .IN1(in2[4]), .IN2(n87), .IN3(n86), .IN4(n24), .IN5(n26), 
        .IN6(n89), .Q(out1[4]) );
  NOR2X0 U53 ( .IN1(in2[5]), .IN2(n25), .QN(n27) );
  AOI21X1 U54 ( .IN1(in2[5]), .IN2(n25), .IN3(n27), .QN(n28) );
  AO222X1 U55 ( .IN1(in2[5]), .IN2(n87), .IN3(n86), .IN4(n26), .IN5(n28), 
        .IN6(n89), .Q(out1[5]) );
  OA21X1 U56 ( .IN1(n27), .IN2(n5), .IN3(n29), .Q(n30) );
  AO222X1 U57 ( .IN1(in2[6]), .IN2(n87), .IN3(n86), .IN4(n28), .IN5(n30), 
        .IN6(n89), .Q(out1[6]) );
  NOR2X0 U58 ( .IN1(in2[7]), .IN2(n29), .QN(n31) );
  AOI21X1 U59 ( .IN1(in2[7]), .IN2(n29), .IN3(n31), .QN(n32) );
  AO222X1 U60 ( .IN1(in2[7]), .IN2(n87), .IN3(n86), .IN4(n30), .IN5(n32), 
        .IN6(n89), .Q(out1[7]) );
  OA21X1 U61 ( .IN1(n31), .IN2(n6), .IN3(n33), .Q(n34) );
  AO222X1 U62 ( .IN1(in2[8]), .IN2(n87), .IN3(n86), .IN4(n32), .IN5(n34), 
        .IN6(n89), .Q(out1[8]) );
  NOR2X0 U63 ( .IN1(in2[9]), .IN2(n33), .QN(n35) );
  AOI21X1 U64 ( .IN1(in2[9]), .IN2(n33), .IN3(n35), .QN(n36) );
  AO222X1 U65 ( .IN1(in2[9]), .IN2(n87), .IN3(n86), .IN4(n34), .IN5(n36), 
        .IN6(n89), .Q(out1[9]) );
  OA21X1 U66 ( .IN1(n35), .IN2(n7), .IN3(n37), .Q(n38) );
  AO222X1 U67 ( .IN1(in2[10]), .IN2(n87), .IN3(n86), .IN4(n36), .IN5(n38), 
        .IN6(n89), .Q(out1[10]) );
  NOR2X0 U68 ( .IN1(in2[11]), .IN2(n37), .QN(n39) );
  AOI21X1 U69 ( .IN1(in2[11]), .IN2(n37), .IN3(n39), .QN(n40) );
  AO222X1 U70 ( .IN1(in2[11]), .IN2(n87), .IN3(n86), .IN4(n38), .IN5(n40), 
        .IN6(n89), .Q(out1[11]) );
  OA21X1 U71 ( .IN1(n39), .IN2(n8), .IN3(n44), .Q(n42) );
  AO222X1 U72 ( .IN1(in2[12]), .IN2(n87), .IN3(n86), .IN4(n40), .IN5(n42), 
        .IN6(n89), .Q(out1[12]) );
  MUX21X1 U73 ( .IN1(n9), .IN2(in2[13]), .S(n41), .Q(n43) );
  AO22X1 U74 ( .IN1(in1[1]), .IN2(n43), .IN3(n86), .IN4(n42), .Q(out1[13]) );
  NOR2X0 U75 ( .IN1(in2[13]), .IN2(n44), .QN(n49) );
  AO21X1 U76 ( .IN1(in2[13]), .IN2(n44), .IN3(n83), .Q(n47) );
  NOR2X0 U77 ( .IN1(n49), .IN2(n69), .QN(n45) );
  MUX21X1 U78 ( .IN1(n10), .IN2(in2[14]), .S(n45), .Q(n46) );
  OAI22X1 U79 ( .IN1(n49), .IN2(n47), .IN3(n72), .IN4(n46), .QN(out1[14]) );
  MUX21X1 U80 ( .IN1(n11), .IN2(in2[15]), .S(n48), .Q(n51) );
  OA21X1 U81 ( .IN1(n49), .IN2(n10), .IN3(n86), .Q(n50) );
  AO22X1 U82 ( .IN1(in1[1]), .IN2(n51), .IN3(n50), .IN4(n52), .Q(out1[15]) );
  NOR2X0 U83 ( .IN1(in2[15]), .IN2(n52), .QN(n57) );
  AO21X1 U84 ( .IN1(in2[15]), .IN2(n52), .IN3(n83), .Q(n55) );
  NOR2X0 U85 ( .IN1(n57), .IN2(n69), .QN(n53) );
  MUX21X1 U86 ( .IN1(n12), .IN2(in2[16]), .S(n53), .Q(n54) );
  OAI22X1 U87 ( .IN1(n57), .IN2(n55), .IN3(n72), .IN4(n54), .QN(out1[16]) );
  MUX21X1 U88 ( .IN1(n13), .IN2(in2[17]), .S(n56), .Q(n59) );
  OA21X1 U89 ( .IN1(n57), .IN2(n12), .IN3(n86), .Q(n58) );
  AO22X1 U90 ( .IN1(in1[1]), .IN2(n59), .IN3(n58), .IN4(n60), .Q(out1[17]) );
  NOR2X0 U91 ( .IN1(in2[17]), .IN2(n60), .QN(n65) );
  AO21X1 U92 ( .IN1(in2[17]), .IN2(n60), .IN3(n83), .Q(n63) );
  NOR2X0 U93 ( .IN1(n65), .IN2(n69), .QN(n61) );
  MUX21X1 U94 ( .IN1(n14), .IN2(in2[18]), .S(n61), .Q(n62) );
  OAI22X1 U95 ( .IN1(n65), .IN2(n63), .IN3(n72), .IN4(n62), .QN(out1[18]) );
  MUX21X1 U96 ( .IN1(n15), .IN2(in2[19]), .S(n64), .Q(n67) );
  OA21X1 U97 ( .IN1(n65), .IN2(n14), .IN3(n86), .Q(n66) );
  AO22X1 U98 ( .IN1(in1[1]), .IN2(n67), .IN3(n66), .IN4(n68), .Q(out1[19]) );
  NOR2X0 U99 ( .IN1(in2[19]), .IN2(n68), .QN(n75) );
  AO21X1 U100 ( .IN1(in2[19]), .IN2(n68), .IN3(n83), .Q(n73) );
  NOR2X0 U101 ( .IN1(n75), .IN2(n69), .QN(n70) );
  MUX21X1 U102 ( .IN1(n16), .IN2(in2[20]), .S(n70), .Q(n71) );
  OAI22X1 U103 ( .IN1(n75), .IN2(n73), .IN3(n72), .IN4(n71), .QN(out1[20]) );
  MUX21X1 U104 ( .IN1(n17), .IN2(in2[21]), .S(n74), .Q(n77) );
  MUX21X1 U105 ( .IN1(n16), .IN2(in2[20]), .S(n75), .Q(n76) );
  AO22X1 U106 ( .IN1(in1[1]), .IN2(n77), .IN3(n86), .IN4(n76), .Q(out1[21]) );
  INVX0 U107 ( .INP(n89), .ZN(n78) );
  OR2X1 U108 ( .IN1(n79), .IN2(in2[21]), .Q(n85) );
  NOR2X0 U109 ( .IN1(n78), .IN2(n85), .QN(n84) );
  NOR2X0 U110 ( .IN1(in2[22]), .IN2(n78), .QN(n81) );
  OA221X1 U111 ( .IN1(n81), .IN2(n86), .IN3(n81), .IN4(n80), .IN5(n85), .Q(n82) );
  AO221X1 U112 ( .IN1(in2[22]), .IN2(n87), .IN3(in2[22]), .IN4(n84), .IN5(n82), 
        .Q(out1[22]) );
  NOR2X0 U113 ( .IN1(n83), .IN2(n85), .QN(n90) );
  AO21X1 U114 ( .IN1(n86), .IN2(n85), .IN3(n84), .Q(n88) );
  AO221X1 U115 ( .IN1(in2[22]), .IN2(n90), .IN3(n18), .IN4(n88), .IN5(n87), 
        .Q(out1[23]) );
  AO21X1 U116 ( .IN1(n90), .IN2(n18), .IN3(n89), .Q(out1[24]) );
  AND2X1 U117 ( .IN1(in1[1]), .IN2(in2[0]), .Q(out1[0]) );
endmodule


module booth27_72 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2;

  AND2X1 U3 ( .IN1(in1[1]), .IN2(in1[0]), .Q(out1[24]) );
  INVX0 U4 ( .INP(in1[1]), .ZN(n1) );
  MUX21X1 U5 ( .IN1(in1[1]), .IN2(n1), .S(in1[0]), .Q(n2) );
  AO22X1 U6 ( .IN1(in2[0]), .IN2(out1[24]), .IN3(in2[1]), .IN4(n2), .Q(out1[1]) );
  AO22X1 U7 ( .IN1(out1[24]), .IN2(in2[1]), .IN3(in2[2]), .IN4(n2), .Q(out1[2]) );
  AO22X1 U8 ( .IN1(out1[24]), .IN2(in2[2]), .IN3(in2[3]), .IN4(n2), .Q(out1[3]) );
  AO22X1 U9 ( .IN1(out1[24]), .IN2(in2[3]), .IN3(in2[4]), .IN4(n2), .Q(out1[4]) );
  AO22X1 U10 ( .IN1(out1[24]), .IN2(in2[4]), .IN3(in2[5]), .IN4(n2), .Q(
        out1[5]) );
  AO22X1 U11 ( .IN1(out1[24]), .IN2(in2[5]), .IN3(in2[6]), .IN4(n2), .Q(
        out1[6]) );
  AO22X1 U12 ( .IN1(out1[24]), .IN2(in2[6]), .IN3(in2[7]), .IN4(n2), .Q(
        out1[7]) );
  AO22X1 U13 ( .IN1(out1[24]), .IN2(in2[7]), .IN3(in2[8]), .IN4(n2), .Q(
        out1[8]) );
  AO22X1 U14 ( .IN1(out1[24]), .IN2(in2[8]), .IN3(in2[9]), .IN4(n2), .Q(
        out1[9]) );
  AO22X1 U15 ( .IN1(out1[24]), .IN2(in2[9]), .IN3(in2[10]), .IN4(n2), .Q(
        out1[10]) );
  AO22X1 U16 ( .IN1(out1[24]), .IN2(in2[10]), .IN3(in2[11]), .IN4(n2), .Q(
        out1[11]) );
  AO22X1 U17 ( .IN1(out1[24]), .IN2(in2[11]), .IN3(in2[12]), .IN4(n2), .Q(
        out1[12]) );
  AO22X1 U18 ( .IN1(out1[24]), .IN2(in2[12]), .IN3(in2[13]), .IN4(n2), .Q(
        out1[13]) );
  AO22X1 U19 ( .IN1(out1[24]), .IN2(in2[13]), .IN3(in2[14]), .IN4(n2), .Q(
        out1[14]) );
  AO22X1 U20 ( .IN1(out1[24]), .IN2(in2[14]), .IN3(in2[15]), .IN4(n2), .Q(
        out1[15]) );
  AO22X1 U21 ( .IN1(out1[24]), .IN2(in2[15]), .IN3(in2[16]), .IN4(n2), .Q(
        out1[16]) );
  AO22X1 U22 ( .IN1(out1[24]), .IN2(in2[16]), .IN3(in2[17]), .IN4(n2), .Q(
        out1[17]) );
  AO22X1 U23 ( .IN1(out1[24]), .IN2(in2[17]), .IN3(in2[18]), .IN4(n2), .Q(
        out1[18]) );
  AO22X1 U24 ( .IN1(out1[24]), .IN2(in2[18]), .IN3(in2[19]), .IN4(n2), .Q(
        out1[19]) );
  AO22X1 U25 ( .IN1(out1[24]), .IN2(in2[19]), .IN3(in2[20]), .IN4(n2), .Q(
        out1[20]) );
  AO22X1 U26 ( .IN1(out1[24]), .IN2(in2[20]), .IN3(in2[21]), .IN4(n2), .Q(
        out1[21]) );
  AO22X1 U27 ( .IN1(out1[24]), .IN2(in2[21]), .IN3(in2[22]), .IN4(n2), .Q(
        out1[22]) );
  AO21X1 U28 ( .IN1(out1[24]), .IN2(in2[22]), .IN3(n2), .Q(out1[23]) );
  AND2X1 U29 ( .IN1(in2[0]), .IN2(n2), .Q(out1[0]) );
endmodule


module booth27_73 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n57), .IN2(n10), .QN(n61) );
  NAND2X0 U4 ( .IN1(n25), .IN2(n6), .QN(n30) );
  NAND2X0 U5 ( .IN1(n33), .IN2(n7), .QN(n37) );
  NAND2X0 U6 ( .IN1(n49), .IN2(n9), .QN(n53) );
  NAND2X0 U7 ( .IN1(n41), .IN2(n8), .QN(n45) );
  NAND2X0 U8 ( .IN1(n65), .IN2(n11), .QN(n77) );
  NAND2X0 U9 ( .IN1(n81), .IN2(n13), .QN(n89) );
  NAND2X0 U10 ( .IN1(n93), .IN2(n15), .QN(n101) );
  NAND2X0 U11 ( .IN1(n105), .IN2(n17), .QN(n114) );
  NAND2X0 U12 ( .IN1(in1[2]), .IN2(n77), .QN(n71) );
  NAND2X0 U13 ( .IN1(n70), .IN2(n132), .QN(n74) );
  NAND2X0 U14 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U15 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U16 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U17 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U18 ( .IN1(n118), .IN2(n19), .QN(n125) );
  NAND2X0 U19 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U20 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U21 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U22 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U23 ( .IN1(n141), .IN2(n130), .QN(n24) );
  NAND2X0 U24 ( .IN1(n27), .IN2(n132), .QN(n4) );
  NAND2X0 U25 ( .IN1(n56), .IN2(n55), .QN(out1[9]) );
  NAND2X0 U26 ( .IN1(n60), .IN2(n59), .QN(out1[10]) );
  NAND2X0 U27 ( .IN1(n64), .IN2(n63), .QN(out1[11]) );
  NAND2X0 U28 ( .IN1(n69), .IN2(n68), .QN(out1[12]) );
  NAND2X0 U29 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U30 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U31 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NAND2X0 U32 ( .IN1(n32), .IN2(n31), .QN(out1[3]) );
  NAND2X0 U33 ( .IN1(n36), .IN2(n35), .QN(out1[4]) );
  NAND2X0 U34 ( .IN1(n40), .IN2(n39), .QN(out1[5]) );
  NAND2X0 U35 ( .IN1(n44), .IN2(n43), .QN(out1[6]) );
  NAND2X0 U36 ( .IN1(n48), .IN2(n47), .QN(out1[7]) );
  NAND2X0 U37 ( .IN1(n52), .IN2(n51), .QN(out1[8]) );
  NAND2X0 U38 ( .IN1(n23), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U39 ( .IN1(in1[2]), .IN2(n22), .QN(n23) );
  NOR2X0 U40 ( .IN1(n28), .IN2(n26), .QN(n3) );
  INVX0 U41 ( .INP(n130), .ZN(n137) );
  NAND3X0 U42 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  NOR2X0 U43 ( .IN1(n142), .IN2(n21), .QN(n1) );
  INVX0 U44 ( .INP(n132), .ZN(n141) );
  NOR3X0 U45 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  NOR2X0 U46 ( .IN1(n142), .IN2(n111), .QN(n138) );
  MUX21X1 U47 ( .IN1(n22), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  INVX0 U48 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U49 ( .INP(in2[2]), .ZN(n6) );
  INVX0 U50 ( .INP(in2[4]), .ZN(n7) );
  INVX0 U51 ( .INP(in2[6]), .ZN(n8) );
  INVX0 U52 ( .INP(in2[8]), .ZN(n9) );
  INVX0 U53 ( .INP(in2[10]), .ZN(n10) );
  INVX0 U54 ( .INP(in2[12]), .ZN(n11) );
  INVX0 U55 ( .INP(in2[13]), .ZN(n12) );
  INVX0 U56 ( .INP(in2[14]), .ZN(n13) );
  INVX0 U57 ( .INP(in2[15]), .ZN(n14) );
  INVX0 U58 ( .INP(in2[16]), .ZN(n15) );
  INVX0 U59 ( .INP(in2[17]), .ZN(n16) );
  INVX0 U60 ( .INP(in2[18]), .ZN(n17) );
  INVX0 U61 ( .INP(in2[19]), .ZN(n18) );
  INVX0 U62 ( .INP(in2[20]), .ZN(n19) );
  INVX0 U63 ( .INP(in2[21]), .ZN(n20) );
  INVX0 U64 ( .INP(in2[22]), .ZN(n21) );
  INVX0 U65 ( .INP(in1[1]), .ZN(n22) );
  INVX0 U66 ( .INP(in1[2]), .ZN(n111) );
  INVX0 U67 ( .INP(n138), .ZN(n140) );
  NOR2X0 U68 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n25) );
  AOI21X1 U69 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n25), .QN(n27) );
  NOR2X0 U70 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U71 ( .IN1(n24), .IN2(in2[0]), .IN3(n138), .IN4(n27), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U72 ( .INP(n133), .ZN(n67) );
  NOR2X0 U73 ( .IN1(n67), .IN2(n6), .QN(n28) );
  OA21X1 U74 ( .IN1(n25), .IN2(n6), .IN3(n30), .Q(n29) );
  AO22X1 U75 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n29), .Q(n26) );
  AOI22X1 U76 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n29), .QN(n32) );
  NOR2X0 U77 ( .IN1(in2[3]), .IN2(n30), .QN(n33) );
  AO21X1 U78 ( .IN1(in2[3]), .IN2(n30), .IN3(n33), .Q(n34) );
  OA22X1 U79 ( .IN1(n6), .IN2(n130), .IN3(n140), .IN4(n34), .Q(n31) );
  OA21X1 U80 ( .IN1(n33), .IN2(n7), .IN3(n37), .Q(n38) );
  AOI22X1 U81 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n38), .QN(n36) );
  OA22X1 U82 ( .IN1(n67), .IN2(n7), .IN3(n141), .IN4(n34), .Q(n35) );
  NOR2X0 U83 ( .IN1(in2[5]), .IN2(n37), .QN(n41) );
  AO21X1 U84 ( .IN1(in2[5]), .IN2(n37), .IN3(n41), .Q(n42) );
  OA22X1 U85 ( .IN1(n7), .IN2(n130), .IN3(n140), .IN4(n42), .Q(n40) );
  AOI22X1 U86 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n38), .QN(n39) );
  OA21X1 U87 ( .IN1(n41), .IN2(n8), .IN3(n45), .Q(n46) );
  AOI22X1 U88 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n46), .QN(n44) );
  OA22X1 U89 ( .IN1(n67), .IN2(n8), .IN3(n141), .IN4(n42), .Q(n43) );
  NOR2X0 U90 ( .IN1(in2[7]), .IN2(n45), .QN(n49) );
  AO21X1 U91 ( .IN1(in2[7]), .IN2(n45), .IN3(n49), .Q(n50) );
  OA22X1 U92 ( .IN1(n8), .IN2(n130), .IN3(n140), .IN4(n50), .Q(n48) );
  AOI22X1 U93 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n46), .QN(n47) );
  OA21X1 U94 ( .IN1(n49), .IN2(n9), .IN3(n53), .Q(n54) );
  AOI22X1 U95 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n54), .QN(n52) );
  OA22X1 U96 ( .IN1(n67), .IN2(n9), .IN3(n141), .IN4(n50), .Q(n51) );
  NOR2X0 U97 ( .IN1(in2[9]), .IN2(n53), .QN(n57) );
  AO21X1 U98 ( .IN1(in2[9]), .IN2(n53), .IN3(n57), .Q(n58) );
  OA22X1 U99 ( .IN1(n9), .IN2(n130), .IN3(n140), .IN4(n58), .Q(n56) );
  AOI22X1 U100 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n54), .QN(n55) );
  OA21X1 U101 ( .IN1(n57), .IN2(n10), .IN3(n61), .Q(n62) );
  AOI22X1 U102 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n62), .QN(n60) );
  OA22X1 U103 ( .IN1(n67), .IN2(n10), .IN3(n141), .IN4(n58), .Q(n59) );
  NOR2X0 U104 ( .IN1(in2[11]), .IN2(n61), .QN(n65) );
  AO21X1 U105 ( .IN1(in2[11]), .IN2(n61), .IN3(n65), .Q(n66) );
  OA22X1 U106 ( .IN1(n10), .IN2(n130), .IN3(n140), .IN4(n66), .Q(n64) );
  AOI22X1 U107 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n62), .QN(n63) );
  OA21X1 U108 ( .IN1(n65), .IN2(n11), .IN3(n77), .Q(n70) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n70), .QN(n69) );
  OA22X1 U110 ( .IN1(n67), .IN2(n11), .IN3(n141), .IN4(n66), .Q(n68) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n12), .S(n71), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n11), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n13), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n12), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n12), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n14), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n13), .IN4(n85), .IN5(n84), 
        .Q(out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n15), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n14), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n14), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n16), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n15), .IN4(n97), .IN5(n96), 
        .Q(out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n17), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n16), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n16), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n18), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n17), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n19), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n18), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n18), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n20), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n19), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n21), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n20), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n20), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n21), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_74 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n25), .IN2(n6), .QN(n30) );
  NAND2X0 U4 ( .IN1(n33), .IN2(n7), .QN(n37) );
  NAND2X0 U5 ( .IN1(n41), .IN2(n8), .QN(n45) );
  NAND2X0 U6 ( .IN1(n57), .IN2(n10), .QN(n61) );
  NAND2X0 U7 ( .IN1(n49), .IN2(n9), .QN(n53) );
  NAND2X0 U8 ( .IN1(n65), .IN2(n11), .QN(n77) );
  NAND2X0 U9 ( .IN1(n81), .IN2(n13), .QN(n89) );
  NAND2X0 U10 ( .IN1(n93), .IN2(n15), .QN(n101) );
  NAND2X0 U11 ( .IN1(n105), .IN2(n17), .QN(n114) );
  NAND2X0 U12 ( .IN1(n118), .IN2(n19), .QN(n125) );
  NAND2X0 U13 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U14 ( .IN1(in1[2]), .IN2(n77), .QN(n71) );
  NAND2X0 U15 ( .IN1(n70), .IN2(n132), .QN(n74) );
  NAND2X0 U16 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U17 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U18 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U19 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U20 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U21 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U22 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U23 ( .IN1(n141), .IN2(n130), .QN(n24) );
  NAND2X0 U24 ( .IN1(n27), .IN2(n132), .QN(n4) );
  NAND2X0 U25 ( .IN1(n64), .IN2(n63), .QN(out1[11]) );
  NAND2X0 U26 ( .IN1(n69), .IN2(n68), .QN(out1[12]) );
  NAND2X0 U27 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U28 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U29 ( .IN1(n23), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U30 ( .IN1(in1[2]), .IN2(n22), .QN(n23) );
  NAND2X0 U31 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NAND2X0 U32 ( .IN1(n32), .IN2(n31), .QN(out1[3]) );
  NAND2X0 U33 ( .IN1(n36), .IN2(n35), .QN(out1[4]) );
  NAND2X0 U34 ( .IN1(n40), .IN2(n39), .QN(out1[5]) );
  NAND2X0 U35 ( .IN1(n44), .IN2(n43), .QN(out1[6]) );
  NAND2X0 U36 ( .IN1(n48), .IN2(n47), .QN(out1[7]) );
  NAND2X0 U37 ( .IN1(n52), .IN2(n51), .QN(out1[8]) );
  NAND2X0 U38 ( .IN1(n56), .IN2(n55), .QN(out1[9]) );
  NAND2X0 U39 ( .IN1(n60), .IN2(n59), .QN(out1[10]) );
  NOR2X0 U40 ( .IN1(n28), .IN2(n26), .QN(n3) );
  NOR2X0 U41 ( .IN1(n142), .IN2(n21), .QN(n1) );
  INVX0 U42 ( .INP(n132), .ZN(n141) );
  INVX0 U43 ( .INP(n130), .ZN(n137) );
  NAND3X0 U44 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  NOR3X0 U45 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  NOR2X0 U46 ( .IN1(n142), .IN2(n111), .QN(n138) );
  MUX21X1 U47 ( .IN1(n22), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  INVX0 U48 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U49 ( .INP(in2[2]), .ZN(n6) );
  INVX0 U50 ( .INP(in2[4]), .ZN(n7) );
  INVX0 U51 ( .INP(in2[6]), .ZN(n8) );
  INVX0 U52 ( .INP(in2[8]), .ZN(n9) );
  INVX0 U53 ( .INP(in2[10]), .ZN(n10) );
  INVX0 U54 ( .INP(in2[12]), .ZN(n11) );
  INVX0 U55 ( .INP(in2[13]), .ZN(n12) );
  INVX0 U56 ( .INP(in2[14]), .ZN(n13) );
  INVX0 U57 ( .INP(in2[15]), .ZN(n14) );
  INVX0 U58 ( .INP(in2[16]), .ZN(n15) );
  INVX0 U59 ( .INP(in2[17]), .ZN(n16) );
  INVX0 U60 ( .INP(in2[18]), .ZN(n17) );
  INVX0 U61 ( .INP(in2[19]), .ZN(n18) );
  INVX0 U62 ( .INP(in2[20]), .ZN(n19) );
  INVX0 U63 ( .INP(in2[21]), .ZN(n20) );
  INVX0 U64 ( .INP(in2[22]), .ZN(n21) );
  INVX0 U65 ( .INP(in1[1]), .ZN(n22) );
  INVX0 U66 ( .INP(in1[2]), .ZN(n111) );
  INVX0 U67 ( .INP(n138), .ZN(n140) );
  NOR2X0 U68 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n25) );
  AOI21X1 U69 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n25), .QN(n27) );
  NOR2X0 U70 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U71 ( .IN1(n24), .IN2(in2[0]), .IN3(n138), .IN4(n27), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U72 ( .INP(n133), .ZN(n67) );
  NOR2X0 U73 ( .IN1(n67), .IN2(n6), .QN(n28) );
  OA21X1 U74 ( .IN1(n25), .IN2(n6), .IN3(n30), .Q(n29) );
  AO22X1 U75 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n29), .Q(n26) );
  AOI22X1 U76 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n29), .QN(n32) );
  NOR2X0 U77 ( .IN1(in2[3]), .IN2(n30), .QN(n33) );
  AO21X1 U78 ( .IN1(in2[3]), .IN2(n30), .IN3(n33), .Q(n34) );
  OA22X1 U79 ( .IN1(n6), .IN2(n130), .IN3(n140), .IN4(n34), .Q(n31) );
  OA21X1 U80 ( .IN1(n33), .IN2(n7), .IN3(n37), .Q(n38) );
  AOI22X1 U81 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n38), .QN(n36) );
  OA22X1 U82 ( .IN1(n67), .IN2(n7), .IN3(n141), .IN4(n34), .Q(n35) );
  NOR2X0 U83 ( .IN1(in2[5]), .IN2(n37), .QN(n41) );
  AO21X1 U84 ( .IN1(in2[5]), .IN2(n37), .IN3(n41), .Q(n42) );
  OA22X1 U85 ( .IN1(n7), .IN2(n130), .IN3(n140), .IN4(n42), .Q(n40) );
  AOI22X1 U86 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n38), .QN(n39) );
  OA21X1 U87 ( .IN1(n41), .IN2(n8), .IN3(n45), .Q(n46) );
  AOI22X1 U88 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n46), .QN(n44) );
  OA22X1 U89 ( .IN1(n67), .IN2(n8), .IN3(n141), .IN4(n42), .Q(n43) );
  NOR2X0 U90 ( .IN1(in2[7]), .IN2(n45), .QN(n49) );
  AO21X1 U91 ( .IN1(in2[7]), .IN2(n45), .IN3(n49), .Q(n50) );
  OA22X1 U92 ( .IN1(n8), .IN2(n130), .IN3(n140), .IN4(n50), .Q(n48) );
  AOI22X1 U93 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n46), .QN(n47) );
  OA21X1 U94 ( .IN1(n49), .IN2(n9), .IN3(n53), .Q(n54) );
  AOI22X1 U95 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n54), .QN(n52) );
  OA22X1 U96 ( .IN1(n67), .IN2(n9), .IN3(n141), .IN4(n50), .Q(n51) );
  NOR2X0 U97 ( .IN1(in2[9]), .IN2(n53), .QN(n57) );
  AO21X1 U98 ( .IN1(in2[9]), .IN2(n53), .IN3(n57), .Q(n58) );
  OA22X1 U99 ( .IN1(n9), .IN2(n130), .IN3(n140), .IN4(n58), .Q(n56) );
  AOI22X1 U100 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n54), .QN(n55) );
  OA21X1 U101 ( .IN1(n57), .IN2(n10), .IN3(n61), .Q(n62) );
  AOI22X1 U102 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n62), .QN(n60) );
  OA22X1 U103 ( .IN1(n67), .IN2(n10), .IN3(n141), .IN4(n58), .Q(n59) );
  NOR2X0 U104 ( .IN1(in2[11]), .IN2(n61), .QN(n65) );
  AO21X1 U105 ( .IN1(in2[11]), .IN2(n61), .IN3(n65), .Q(n66) );
  OA22X1 U106 ( .IN1(n10), .IN2(n130), .IN3(n140), .IN4(n66), .Q(n64) );
  AOI22X1 U107 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n62), .QN(n63) );
  OA21X1 U108 ( .IN1(n65), .IN2(n11), .IN3(n77), .Q(n70) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n70), .QN(n69) );
  OA22X1 U110 ( .IN1(n67), .IN2(n11), .IN3(n141), .IN4(n66), .Q(n68) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n12), .S(n71), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n11), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n13), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n12), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n12), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n14), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n13), .IN4(n85), .IN5(n84), 
        .Q(out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n15), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n14), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n14), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n16), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n15), .IN4(n97), .IN5(n96), 
        .Q(out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n17), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n16), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n16), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n18), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n17), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n19), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n18), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n18), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n20), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n19), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n21), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n20), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n20), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n21), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_75 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90;

  NAND2X0 U3 ( .IN1(n75), .IN2(n16), .QN(n79) );
  NAND2X0 U4 ( .IN1(n23), .IN2(n4), .QN(n25) );
  NAND2X0 U5 ( .IN1(n27), .IN2(n5), .QN(n29) );
  NAND2X0 U6 ( .IN1(n31), .IN2(n6), .QN(n33) );
  NAND2X0 U7 ( .IN1(n35), .IN2(n7), .QN(n37) );
  NAND2X0 U8 ( .IN1(n39), .IN2(n8), .QN(n44) );
  NAND2X0 U9 ( .IN1(in1[2]), .IN2(n44), .QN(n41) );
  NAND2X0 U10 ( .IN1(n49), .IN2(n10), .QN(n52) );
  NAND2X0 U11 ( .IN1(in1[2]), .IN2(n52), .QN(n48) );
  NAND2X0 U12 ( .IN1(n57), .IN2(n12), .QN(n60) );
  NAND2X0 U13 ( .IN1(in1[2]), .IN2(n60), .QN(n56) );
  NAND2X0 U14 ( .IN1(n65), .IN2(n14), .QN(n68) );
  NAND2X0 U15 ( .IN1(in1[2]), .IN2(n68), .QN(n64) );
  NAND2X0 U16 ( .IN1(in1[2]), .IN2(n79), .QN(n74) );
  NAND2X0 U17 ( .IN1(in2[21]), .IN2(n79), .QN(n80) );
  NAND2X0 U18 ( .IN1(n72), .IN2(in1[2]), .QN(n83) );
  INVX0 U19 ( .INP(n83), .ZN(n86) );
  INVX0 U20 ( .INP(in1[0]), .ZN(n72) );
  NOR2X0 U21 ( .IN1(in1[2]), .IN2(n72), .QN(n87) );
  NOR2X0 U22 ( .IN1(n72), .IN2(n69), .QN(n89) );
  NBUFFX2 U23 ( .INP(in1[2]), .Z(out1[25]) );
  NBUFFX2 U24 ( .INP(in1[2]), .Z(out1[26]) );
  INVX0 U25 ( .INP(in2[2]), .ZN(n3) );
  INVX0 U26 ( .INP(in2[4]), .ZN(n4) );
  INVX0 U27 ( .INP(in2[6]), .ZN(n5) );
  INVX0 U28 ( .INP(in2[8]), .ZN(n6) );
  INVX0 U29 ( .INP(in2[10]), .ZN(n7) );
  INVX0 U30 ( .INP(in2[12]), .ZN(n8) );
  INVX0 U31 ( .INP(in2[13]), .ZN(n9) );
  INVX0 U32 ( .INP(in2[14]), .ZN(n10) );
  INVX0 U33 ( .INP(in2[15]), .ZN(n11) );
  INVX0 U34 ( .INP(in2[16]), .ZN(n12) );
  INVX0 U35 ( .INP(in2[17]), .ZN(n13) );
  INVX0 U36 ( .INP(in2[18]), .ZN(n14) );
  INVX0 U37 ( .INP(in2[19]), .ZN(n15) );
  INVX0 U38 ( .INP(in2[20]), .ZN(n16) );
  INVX0 U39 ( .INP(in2[21]), .ZN(n17) );
  INVX0 U40 ( .INP(in2[22]), .ZN(n18) );
  INVX0 U41 ( .INP(in1[2]), .ZN(n69) );
  NOR2X0 U42 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n19) );
  AOI21X1 U43 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n19), .QN(n20) );
  AO222X1 U44 ( .IN1(in2[0]), .IN2(n86), .IN3(in2[1]), .IN4(n87), .IN5(n89), 
        .IN6(n20), .Q(out1[1]) );
  OR3X1 U45 ( .IN1(in2[2]), .IN2(in2[0]), .IN3(in2[1]), .Q(n21) );
  OA21X1 U46 ( .IN1(n19), .IN2(n3), .IN3(n21), .Q(n22) );
  AO222X1 U47 ( .IN1(in2[2]), .IN2(n87), .IN3(n86), .IN4(n20), .IN5(n22), 
        .IN6(n89), .Q(out1[2]) );
  NOR2X0 U48 ( .IN1(in2[3]), .IN2(n21), .QN(n23) );
  AOI21X1 U49 ( .IN1(in2[3]), .IN2(n21), .IN3(n23), .QN(n24) );
  AO222X1 U50 ( .IN1(in2[3]), .IN2(n87), .IN3(n86), .IN4(n22), .IN5(n24), 
        .IN6(n89), .Q(out1[3]) );
  OA21X1 U51 ( .IN1(n23), .IN2(n4), .IN3(n25), .Q(n26) );
  AO222X1 U52 ( .IN1(in2[4]), .IN2(n87), .IN3(n86), .IN4(n24), .IN5(n26), 
        .IN6(n89), .Q(out1[4]) );
  NOR2X0 U53 ( .IN1(in2[5]), .IN2(n25), .QN(n27) );
  AOI21X1 U54 ( .IN1(in2[5]), .IN2(n25), .IN3(n27), .QN(n28) );
  AO222X1 U55 ( .IN1(in2[5]), .IN2(n87), .IN3(n86), .IN4(n26), .IN5(n28), 
        .IN6(n89), .Q(out1[5]) );
  OA21X1 U56 ( .IN1(n27), .IN2(n5), .IN3(n29), .Q(n30) );
  AO222X1 U57 ( .IN1(in2[6]), .IN2(n87), .IN3(n86), .IN4(n28), .IN5(n30), 
        .IN6(n89), .Q(out1[6]) );
  NOR2X0 U58 ( .IN1(in2[7]), .IN2(n29), .QN(n31) );
  AOI21X1 U59 ( .IN1(in2[7]), .IN2(n29), .IN3(n31), .QN(n32) );
  AO222X1 U60 ( .IN1(in2[7]), .IN2(n87), .IN3(n86), .IN4(n30), .IN5(n32), 
        .IN6(n89), .Q(out1[7]) );
  OA21X1 U61 ( .IN1(n31), .IN2(n6), .IN3(n33), .Q(n34) );
  AO222X1 U62 ( .IN1(in2[8]), .IN2(n87), .IN3(n86), .IN4(n32), .IN5(n34), 
        .IN6(n89), .Q(out1[8]) );
  NOR2X0 U63 ( .IN1(in2[9]), .IN2(n33), .QN(n35) );
  AOI21X1 U64 ( .IN1(in2[9]), .IN2(n33), .IN3(n35), .QN(n36) );
  AO222X1 U65 ( .IN1(in2[9]), .IN2(n87), .IN3(n86), .IN4(n34), .IN5(n36), 
        .IN6(n89), .Q(out1[9]) );
  OA21X1 U66 ( .IN1(n35), .IN2(n7), .IN3(n37), .Q(n38) );
  AO222X1 U67 ( .IN1(in2[10]), .IN2(n87), .IN3(n86), .IN4(n36), .IN5(n38), 
        .IN6(n89), .Q(out1[10]) );
  NOR2X0 U68 ( .IN1(in2[11]), .IN2(n37), .QN(n39) );
  AOI21X1 U69 ( .IN1(in2[11]), .IN2(n37), .IN3(n39), .QN(n40) );
  AO222X1 U70 ( .IN1(in2[11]), .IN2(n87), .IN3(n86), .IN4(n38), .IN5(n40), 
        .IN6(n89), .Q(out1[11]) );
  OA21X1 U71 ( .IN1(n39), .IN2(n8), .IN3(n44), .Q(n42) );
  AO222X1 U72 ( .IN1(in2[12]), .IN2(n87), .IN3(n86), .IN4(n40), .IN5(n42), 
        .IN6(n89), .Q(out1[12]) );
  MUX21X1 U73 ( .IN1(n9), .IN2(in2[13]), .S(n41), .Q(n43) );
  AO22X1 U74 ( .IN1(in1[0]), .IN2(n43), .IN3(n86), .IN4(n42), .Q(out1[13]) );
  NOR2X0 U75 ( .IN1(in2[13]), .IN2(n44), .QN(n49) );
  AO21X1 U76 ( .IN1(in2[13]), .IN2(n44), .IN3(n83), .Q(n47) );
  NOR2X0 U77 ( .IN1(n49), .IN2(n69), .QN(n45) );
  MUX21X1 U78 ( .IN1(n10), .IN2(in2[14]), .S(n45), .Q(n46) );
  OAI22X1 U79 ( .IN1(n49), .IN2(n47), .IN3(n72), .IN4(n46), .QN(out1[14]) );
  MUX21X1 U80 ( .IN1(n11), .IN2(in2[15]), .S(n48), .Q(n51) );
  OA21X1 U81 ( .IN1(n49), .IN2(n10), .IN3(n86), .Q(n50) );
  AO22X1 U82 ( .IN1(in1[0]), .IN2(n51), .IN3(n50), .IN4(n52), .Q(out1[15]) );
  NOR2X0 U83 ( .IN1(in2[15]), .IN2(n52), .QN(n57) );
  AO21X1 U84 ( .IN1(in2[15]), .IN2(n52), .IN3(n83), .Q(n55) );
  NOR2X0 U85 ( .IN1(n57), .IN2(n69), .QN(n53) );
  MUX21X1 U86 ( .IN1(n12), .IN2(in2[16]), .S(n53), .Q(n54) );
  OAI22X1 U87 ( .IN1(n57), .IN2(n55), .IN3(n72), .IN4(n54), .QN(out1[16]) );
  MUX21X1 U88 ( .IN1(n13), .IN2(in2[17]), .S(n56), .Q(n59) );
  OA21X1 U89 ( .IN1(n57), .IN2(n12), .IN3(n86), .Q(n58) );
  AO22X1 U90 ( .IN1(in1[0]), .IN2(n59), .IN3(n58), .IN4(n60), .Q(out1[17]) );
  NOR2X0 U91 ( .IN1(in2[17]), .IN2(n60), .QN(n65) );
  AO21X1 U92 ( .IN1(in2[17]), .IN2(n60), .IN3(n83), .Q(n63) );
  NOR2X0 U93 ( .IN1(n65), .IN2(n69), .QN(n61) );
  MUX21X1 U94 ( .IN1(n14), .IN2(in2[18]), .S(n61), .Q(n62) );
  OAI22X1 U95 ( .IN1(n65), .IN2(n63), .IN3(n72), .IN4(n62), .QN(out1[18]) );
  MUX21X1 U96 ( .IN1(n15), .IN2(in2[19]), .S(n64), .Q(n67) );
  OA21X1 U97 ( .IN1(n65), .IN2(n14), .IN3(n86), .Q(n66) );
  AO22X1 U98 ( .IN1(in1[0]), .IN2(n67), .IN3(n66), .IN4(n68), .Q(out1[19]) );
  NOR2X0 U99 ( .IN1(in2[19]), .IN2(n68), .QN(n75) );
  AO21X1 U100 ( .IN1(in2[19]), .IN2(n68), .IN3(n83), .Q(n73) );
  NOR2X0 U101 ( .IN1(n75), .IN2(n69), .QN(n70) );
  MUX21X1 U102 ( .IN1(n16), .IN2(in2[20]), .S(n70), .Q(n71) );
  OAI22X1 U103 ( .IN1(n75), .IN2(n73), .IN3(n72), .IN4(n71), .QN(out1[20]) );
  MUX21X1 U104 ( .IN1(n17), .IN2(in2[21]), .S(n74), .Q(n77) );
  MUX21X1 U105 ( .IN1(n16), .IN2(in2[20]), .S(n75), .Q(n76) );
  AO22X1 U106 ( .IN1(in1[0]), .IN2(n77), .IN3(n86), .IN4(n76), .Q(out1[21]) );
  INVX0 U107 ( .INP(n89), .ZN(n78) );
  OR2X1 U108 ( .IN1(n79), .IN2(in2[21]), .Q(n85) );
  NOR2X0 U109 ( .IN1(n78), .IN2(n85), .QN(n84) );
  NOR2X0 U110 ( .IN1(in2[22]), .IN2(n78), .QN(n81) );
  OA221X1 U111 ( .IN1(n81), .IN2(n86), .IN3(n81), .IN4(n80), .IN5(n85), .Q(n82) );
  AO221X1 U112 ( .IN1(in2[22]), .IN2(n87), .IN3(in2[22]), .IN4(n84), .IN5(n82), 
        .Q(out1[22]) );
  NOR2X0 U113 ( .IN1(n83), .IN2(n85), .QN(n90) );
  AO21X1 U114 ( .IN1(n86), .IN2(n85), .IN3(n84), .Q(n88) );
  AO221X1 U115 ( .IN1(in2[22]), .IN2(n90), .IN3(n18), .IN4(n88), .IN5(n87), 
        .Q(out1[23]) );
  AO21X1 U116 ( .IN1(n90), .IN2(n18), .IN3(n89), .Q(out1[24]) );
  AND2X1 U117 ( .IN1(in1[0]), .IN2(in2[0]), .Q(out1[0]) );
endmodule


module booth27_76 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n25), .IN2(n6), .QN(n30) );
  NAND2X0 U4 ( .IN1(n33), .IN2(n7), .QN(n37) );
  NAND2X0 U5 ( .IN1(n41), .IN2(n8), .QN(n45) );
  NAND2X0 U6 ( .IN1(n49), .IN2(n9), .QN(n53) );
  NAND2X0 U7 ( .IN1(n57), .IN2(n10), .QN(n61) );
  NAND2X0 U8 ( .IN1(n65), .IN2(n11), .QN(n77) );
  NAND2X0 U9 ( .IN1(n81), .IN2(n13), .QN(n89) );
  NAND2X0 U10 ( .IN1(n105), .IN2(n17), .QN(n114) );
  NAND2X0 U11 ( .IN1(n93), .IN2(n15), .QN(n101) );
  NAND2X0 U12 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U13 ( .IN1(n118), .IN2(n19), .QN(n125) );
  NAND2X0 U14 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U15 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U16 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U17 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U18 ( .IN1(n27), .IN2(n132), .QN(n4) );
  NAND2X0 U19 ( .IN1(n141), .IN2(n130), .QN(n24) );
  NAND2X0 U20 ( .IN1(n32), .IN2(n31), .QN(out1[3]) );
  NAND2X0 U21 ( .IN1(n36), .IN2(n35), .QN(out1[4]) );
  NAND2X0 U22 ( .IN1(in1[2]), .IN2(n77), .QN(n71) );
  NAND2X0 U23 ( .IN1(n70), .IN2(n132), .QN(n74) );
  NAND2X0 U24 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U25 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U26 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U27 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U28 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NAND2X0 U29 ( .IN1(n40), .IN2(n39), .QN(out1[5]) );
  NAND2X0 U30 ( .IN1(n44), .IN2(n43), .QN(out1[6]) );
  NAND2X0 U31 ( .IN1(n48), .IN2(n47), .QN(out1[7]) );
  NAND2X0 U32 ( .IN1(n52), .IN2(n51), .QN(out1[8]) );
  NAND2X0 U33 ( .IN1(n56), .IN2(n55), .QN(out1[9]) );
  NAND2X0 U34 ( .IN1(n60), .IN2(n59), .QN(out1[10]) );
  NAND2X0 U35 ( .IN1(n64), .IN2(n63), .QN(out1[11]) );
  NAND2X0 U36 ( .IN1(n69), .IN2(n68), .QN(out1[12]) );
  NAND2X0 U37 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U38 ( .IN1(n23), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U39 ( .IN1(in1[2]), .IN2(n22), .QN(n23) );
  NOR2X0 U40 ( .IN1(n28), .IN2(n26), .QN(n3) );
  NOR2X0 U41 ( .IN1(n142), .IN2(n21), .QN(n1) );
  INVX0 U42 ( .INP(n132), .ZN(n141) );
  INVX0 U43 ( .INP(n130), .ZN(n137) );
  NAND3X0 U44 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  NOR3X0 U45 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  NOR2X0 U46 ( .IN1(n142), .IN2(n111), .QN(n138) );
  MUX21X1 U47 ( .IN1(n22), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  INVX0 U48 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U49 ( .INP(in2[2]), .ZN(n6) );
  INVX0 U50 ( .INP(in2[4]), .ZN(n7) );
  INVX0 U51 ( .INP(in2[6]), .ZN(n8) );
  INVX0 U52 ( .INP(in2[8]), .ZN(n9) );
  INVX0 U53 ( .INP(in2[10]), .ZN(n10) );
  INVX0 U54 ( .INP(in2[12]), .ZN(n11) );
  INVX0 U55 ( .INP(in2[13]), .ZN(n12) );
  INVX0 U56 ( .INP(in2[14]), .ZN(n13) );
  INVX0 U57 ( .INP(in2[15]), .ZN(n14) );
  INVX0 U58 ( .INP(in2[16]), .ZN(n15) );
  INVX0 U59 ( .INP(in2[17]), .ZN(n16) );
  INVX0 U60 ( .INP(in2[18]), .ZN(n17) );
  INVX0 U61 ( .INP(in2[19]), .ZN(n18) );
  INVX0 U62 ( .INP(in2[20]), .ZN(n19) );
  INVX0 U63 ( .INP(in2[21]), .ZN(n20) );
  INVX0 U64 ( .INP(in2[22]), .ZN(n21) );
  INVX0 U65 ( .INP(in1[1]), .ZN(n22) );
  INVX0 U66 ( .INP(in1[2]), .ZN(n111) );
  INVX0 U67 ( .INP(n138), .ZN(n140) );
  NOR2X0 U68 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n25) );
  AOI21X1 U69 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n25), .QN(n27) );
  NOR2X0 U70 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U71 ( .IN1(n24), .IN2(in2[0]), .IN3(n138), .IN4(n27), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U72 ( .INP(n133), .ZN(n67) );
  NOR2X0 U73 ( .IN1(n67), .IN2(n6), .QN(n28) );
  OA21X1 U74 ( .IN1(n25), .IN2(n6), .IN3(n30), .Q(n29) );
  AO22X1 U75 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n29), .Q(n26) );
  AOI22X1 U76 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n29), .QN(n32) );
  NOR2X0 U77 ( .IN1(in2[3]), .IN2(n30), .QN(n33) );
  AO21X1 U78 ( .IN1(in2[3]), .IN2(n30), .IN3(n33), .Q(n34) );
  OA22X1 U79 ( .IN1(n6), .IN2(n130), .IN3(n140), .IN4(n34), .Q(n31) );
  OA21X1 U80 ( .IN1(n33), .IN2(n7), .IN3(n37), .Q(n38) );
  AOI22X1 U81 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n38), .QN(n36) );
  OA22X1 U82 ( .IN1(n67), .IN2(n7), .IN3(n141), .IN4(n34), .Q(n35) );
  NOR2X0 U83 ( .IN1(in2[5]), .IN2(n37), .QN(n41) );
  AO21X1 U84 ( .IN1(in2[5]), .IN2(n37), .IN3(n41), .Q(n42) );
  OA22X1 U85 ( .IN1(n7), .IN2(n130), .IN3(n140), .IN4(n42), .Q(n40) );
  AOI22X1 U86 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n38), .QN(n39) );
  OA21X1 U87 ( .IN1(n41), .IN2(n8), .IN3(n45), .Q(n46) );
  AOI22X1 U88 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n46), .QN(n44) );
  OA22X1 U89 ( .IN1(n67), .IN2(n8), .IN3(n141), .IN4(n42), .Q(n43) );
  NOR2X0 U90 ( .IN1(in2[7]), .IN2(n45), .QN(n49) );
  AO21X1 U91 ( .IN1(in2[7]), .IN2(n45), .IN3(n49), .Q(n50) );
  OA22X1 U92 ( .IN1(n8), .IN2(n130), .IN3(n140), .IN4(n50), .Q(n48) );
  AOI22X1 U93 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n46), .QN(n47) );
  OA21X1 U94 ( .IN1(n49), .IN2(n9), .IN3(n53), .Q(n54) );
  AOI22X1 U95 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n54), .QN(n52) );
  OA22X1 U96 ( .IN1(n67), .IN2(n9), .IN3(n141), .IN4(n50), .Q(n51) );
  NOR2X0 U97 ( .IN1(in2[9]), .IN2(n53), .QN(n57) );
  AO21X1 U98 ( .IN1(in2[9]), .IN2(n53), .IN3(n57), .Q(n58) );
  OA22X1 U99 ( .IN1(n9), .IN2(n130), .IN3(n140), .IN4(n58), .Q(n56) );
  AOI22X1 U100 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n54), .QN(n55) );
  OA21X1 U101 ( .IN1(n57), .IN2(n10), .IN3(n61), .Q(n62) );
  AOI22X1 U102 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n62), .QN(n60) );
  OA22X1 U103 ( .IN1(n67), .IN2(n10), .IN3(n141), .IN4(n58), .Q(n59) );
  NOR2X0 U104 ( .IN1(in2[11]), .IN2(n61), .QN(n65) );
  AO21X1 U105 ( .IN1(in2[11]), .IN2(n61), .IN3(n65), .Q(n66) );
  OA22X1 U106 ( .IN1(n10), .IN2(n130), .IN3(n140), .IN4(n66), .Q(n64) );
  AOI22X1 U107 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n62), .QN(n63) );
  OA21X1 U108 ( .IN1(n65), .IN2(n11), .IN3(n77), .Q(n70) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n70), .QN(n69) );
  OA22X1 U110 ( .IN1(n67), .IN2(n11), .IN3(n141), .IN4(n66), .Q(n68) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n12), .S(n71), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n11), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n13), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n12), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n12), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n14), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n13), .IN4(n85), .IN5(n84), 
        .Q(out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n15), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n14), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n14), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n16), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n15), .IN4(n97), .IN5(n96), 
        .Q(out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n17), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n16), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n16), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n18), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n17), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n19), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n18), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n18), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n20), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n19), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n21), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n20), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n20), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n21), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_77 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n33), .IN2(n7), .QN(n37) );
  NAND2X0 U4 ( .IN1(n41), .IN2(n8), .QN(n45) );
  NAND2X0 U5 ( .IN1(n49), .IN2(n9), .QN(n53) );
  NAND2X0 U6 ( .IN1(n57), .IN2(n10), .QN(n61) );
  NAND2X0 U7 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U8 ( .IN1(n25), .IN2(n6), .QN(n30) );
  NAND2X0 U9 ( .IN1(n65), .IN2(n11), .QN(n77) );
  NAND2X0 U10 ( .IN1(n81), .IN2(n13), .QN(n89) );
  NAND2X0 U11 ( .IN1(n93), .IN2(n15), .QN(n101) );
  NAND2X0 U12 ( .IN1(n118), .IN2(n19), .QN(n125) );
  NAND2X0 U13 ( .IN1(n105), .IN2(n17), .QN(n114) );
  NAND2X0 U14 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U15 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U16 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U17 ( .IN1(n40), .IN2(n39), .QN(out1[5]) );
  NAND2X0 U18 ( .IN1(n44), .IN2(n43), .QN(out1[6]) );
  NAND2X0 U19 ( .IN1(in1[2]), .IN2(n77), .QN(n71) );
  NAND2X0 U20 ( .IN1(n70), .IN2(n132), .QN(n74) );
  NAND2X0 U21 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U22 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U23 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U24 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U25 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U26 ( .IN1(n23), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U27 ( .IN1(in1[2]), .IN2(n22), .QN(n23) );
  NAND2X0 U28 ( .IN1(n36), .IN2(n35), .QN(out1[4]) );
  NAND2X0 U29 ( .IN1(n32), .IN2(n31), .QN(out1[3]) );
  NAND2X0 U30 ( .IN1(n27), .IN2(n132), .QN(n4) );
  NAND2X0 U31 ( .IN1(n48), .IN2(n47), .QN(out1[7]) );
  NAND2X0 U32 ( .IN1(n52), .IN2(n51), .QN(out1[8]) );
  NAND2X0 U33 ( .IN1(n56), .IN2(n55), .QN(out1[9]) );
  NAND2X0 U34 ( .IN1(n60), .IN2(n59), .QN(out1[10]) );
  NAND2X0 U35 ( .IN1(n64), .IN2(n63), .QN(out1[11]) );
  NAND2X0 U36 ( .IN1(n69), .IN2(n68), .QN(out1[12]) );
  NAND2X0 U37 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U38 ( .IN1(n141), .IN2(n130), .QN(n24) );
  NAND2X0 U39 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NOR2X0 U40 ( .IN1(n28), .IN2(n26), .QN(n3) );
  INVX0 U41 ( .INP(n130), .ZN(n137) );
  INVX0 U42 ( .INP(n132), .ZN(n141) );
  NOR3X0 U43 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  NAND3X0 U44 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  NOR2X0 U45 ( .IN1(n142), .IN2(n21), .QN(n1) );
  NOR2X0 U46 ( .IN1(n142), .IN2(n111), .QN(n138) );
  MUX21X1 U47 ( .IN1(n22), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  INVX0 U48 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U49 ( .INP(in2[2]), .ZN(n6) );
  INVX0 U50 ( .INP(in2[4]), .ZN(n7) );
  INVX0 U51 ( .INP(in2[6]), .ZN(n8) );
  INVX0 U52 ( .INP(in2[8]), .ZN(n9) );
  INVX0 U53 ( .INP(in2[10]), .ZN(n10) );
  INVX0 U54 ( .INP(in2[12]), .ZN(n11) );
  INVX0 U55 ( .INP(in2[13]), .ZN(n12) );
  INVX0 U56 ( .INP(in2[14]), .ZN(n13) );
  INVX0 U57 ( .INP(in2[15]), .ZN(n14) );
  INVX0 U58 ( .INP(in2[16]), .ZN(n15) );
  INVX0 U59 ( .INP(in2[17]), .ZN(n16) );
  INVX0 U60 ( .INP(in2[18]), .ZN(n17) );
  INVX0 U61 ( .INP(in2[19]), .ZN(n18) );
  INVX0 U62 ( .INP(in2[20]), .ZN(n19) );
  INVX0 U63 ( .INP(in2[21]), .ZN(n20) );
  INVX0 U64 ( .INP(in2[22]), .ZN(n21) );
  INVX0 U65 ( .INP(in1[1]), .ZN(n22) );
  INVX0 U66 ( .INP(in1[2]), .ZN(n111) );
  INVX0 U67 ( .INP(n138), .ZN(n140) );
  NOR2X0 U68 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n25) );
  AOI21X1 U69 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n25), .QN(n27) );
  NOR2X0 U70 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U71 ( .IN1(n24), .IN2(in2[0]), .IN3(n138), .IN4(n27), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U72 ( .INP(n133), .ZN(n67) );
  NOR2X0 U73 ( .IN1(n67), .IN2(n6), .QN(n28) );
  OA21X1 U74 ( .IN1(n25), .IN2(n6), .IN3(n30), .Q(n29) );
  AO22X1 U75 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n29), .Q(n26) );
  AOI22X1 U76 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n29), .QN(n32) );
  NOR2X0 U77 ( .IN1(in2[3]), .IN2(n30), .QN(n33) );
  AO21X1 U78 ( .IN1(in2[3]), .IN2(n30), .IN3(n33), .Q(n34) );
  OA22X1 U79 ( .IN1(n6), .IN2(n130), .IN3(n140), .IN4(n34), .Q(n31) );
  OA21X1 U80 ( .IN1(n33), .IN2(n7), .IN3(n37), .Q(n38) );
  AOI22X1 U81 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n38), .QN(n36) );
  OA22X1 U82 ( .IN1(n67), .IN2(n7), .IN3(n141), .IN4(n34), .Q(n35) );
  NOR2X0 U83 ( .IN1(in2[5]), .IN2(n37), .QN(n41) );
  AO21X1 U84 ( .IN1(in2[5]), .IN2(n37), .IN3(n41), .Q(n42) );
  OA22X1 U85 ( .IN1(n7), .IN2(n130), .IN3(n140), .IN4(n42), .Q(n40) );
  AOI22X1 U86 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n38), .QN(n39) );
  OA21X1 U87 ( .IN1(n41), .IN2(n8), .IN3(n45), .Q(n46) );
  AOI22X1 U88 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n46), .QN(n44) );
  OA22X1 U89 ( .IN1(n67), .IN2(n8), .IN3(n141), .IN4(n42), .Q(n43) );
  NOR2X0 U90 ( .IN1(in2[7]), .IN2(n45), .QN(n49) );
  AO21X1 U91 ( .IN1(in2[7]), .IN2(n45), .IN3(n49), .Q(n50) );
  OA22X1 U92 ( .IN1(n8), .IN2(n130), .IN3(n140), .IN4(n50), .Q(n48) );
  AOI22X1 U93 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n46), .QN(n47) );
  OA21X1 U94 ( .IN1(n49), .IN2(n9), .IN3(n53), .Q(n54) );
  AOI22X1 U95 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n54), .QN(n52) );
  OA22X1 U96 ( .IN1(n67), .IN2(n9), .IN3(n141), .IN4(n50), .Q(n51) );
  NOR2X0 U97 ( .IN1(in2[9]), .IN2(n53), .QN(n57) );
  AO21X1 U98 ( .IN1(in2[9]), .IN2(n53), .IN3(n57), .Q(n58) );
  OA22X1 U99 ( .IN1(n9), .IN2(n130), .IN3(n140), .IN4(n58), .Q(n56) );
  AOI22X1 U100 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n54), .QN(n55) );
  OA21X1 U101 ( .IN1(n57), .IN2(n10), .IN3(n61), .Q(n62) );
  AOI22X1 U102 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n62), .QN(n60) );
  OA22X1 U103 ( .IN1(n67), .IN2(n10), .IN3(n141), .IN4(n58), .Q(n59) );
  NOR2X0 U104 ( .IN1(in2[11]), .IN2(n61), .QN(n65) );
  AO21X1 U105 ( .IN1(in2[11]), .IN2(n61), .IN3(n65), .Q(n66) );
  OA22X1 U106 ( .IN1(n10), .IN2(n130), .IN3(n140), .IN4(n66), .Q(n64) );
  AOI22X1 U107 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n62), .QN(n63) );
  OA21X1 U108 ( .IN1(n65), .IN2(n11), .IN3(n77), .Q(n70) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n70), .QN(n69) );
  OA22X1 U110 ( .IN1(n67), .IN2(n11), .IN3(n141), .IN4(n66), .Q(n68) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n12), .S(n71), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n11), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n13), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n12), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n12), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n14), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n13), .IN4(n85), .IN5(n84), 
        .Q(out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n15), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n14), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n14), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n16), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n15), .IN4(n97), .IN5(n96), 
        .Q(out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n17), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n16), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n16), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n18), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n17), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n19), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n18), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n18), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n20), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n19), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n21), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n20), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n20), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n21), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_78 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93;

  NAND2X0 U3 ( .IN1(n30), .IN2(n7), .QN(n32) );
  NAND2X0 U4 ( .IN1(n34), .IN2(n8), .QN(n36) );
  NAND2X0 U5 ( .IN1(n38), .IN2(n9), .QN(n40) );
  NAND2X0 U6 ( .IN1(n42), .IN2(n10), .QN(n47) );
  NAND2X0 U7 ( .IN1(n78), .IN2(n18), .QN(n82) );
  NAND2X0 U8 ( .IN1(n26), .IN2(n6), .QN(n28) );
  NAND2X0 U9 ( .IN1(in1[2]), .IN2(n47), .QN(n44) );
  NAND2X0 U10 ( .IN1(n52), .IN2(n12), .QN(n55) );
  NAND2X0 U11 ( .IN1(in1[2]), .IN2(n55), .QN(n51) );
  NAND2X0 U12 ( .IN1(n60), .IN2(n14), .QN(n63) );
  NAND2X0 U13 ( .IN1(in1[2]), .IN2(n63), .QN(n59) );
  NAND2X0 U14 ( .IN1(n68), .IN2(n16), .QN(n71) );
  NAND2X0 U15 ( .IN1(in1[2]), .IN2(n71), .QN(n67) );
  NAND2X0 U16 ( .IN1(in1[2]), .IN2(n82), .QN(n77) );
  NAND2X0 U17 ( .IN1(in2[21]), .IN2(n82), .QN(n83) );
  NAND2X0 U18 ( .IN1(n75), .IN2(in1[2]), .QN(n86) );
  NAND2X0 U19 ( .IN1(n3), .IN2(n4), .QN(n22) );
  NAND2X0 U20 ( .IN1(n23), .IN2(n22), .QN(out1[2]) );
  INVX0 U21 ( .INP(n86), .ZN(n89) );
  NAND2X0 U22 ( .IN1(in2[1]), .IN2(in2[0]), .QN(n4) );
  NOR2X0 U23 ( .IN1(n21), .IN2(n86), .QN(n3) );
  NOR2X0 U24 ( .IN1(in1[2]), .IN2(n75), .QN(n90) );
  NOR2X0 U25 ( .IN1(n75), .IN2(n72), .QN(n92) );
  NBUFFX2 U26 ( .INP(in1[2]), .Z(out1[26]) );
  NBUFFX2 U27 ( .INP(in1[2]), .Z(out1[25]) );
  INVX0 U28 ( .INP(in2[2]), .ZN(n5) );
  INVX0 U29 ( .INP(in2[4]), .ZN(n6) );
  INVX0 U30 ( .INP(in2[6]), .ZN(n7) );
  INVX0 U31 ( .INP(in2[8]), .ZN(n8) );
  INVX0 U32 ( .INP(in2[10]), .ZN(n9) );
  INVX0 U33 ( .INP(in2[12]), .ZN(n10) );
  INVX0 U34 ( .INP(in2[13]), .ZN(n11) );
  INVX0 U35 ( .INP(in2[14]), .ZN(n12) );
  INVX0 U36 ( .INP(in2[15]), .ZN(n13) );
  INVX0 U37 ( .INP(in2[16]), .ZN(n14) );
  INVX0 U38 ( .INP(in2[17]), .ZN(n15) );
  INVX0 U39 ( .INP(in2[18]), .ZN(n16) );
  INVX0 U40 ( .INP(in2[19]), .ZN(n17) );
  INVX0 U41 ( .INP(in2[20]), .ZN(n18) );
  INVX0 U42 ( .INP(in2[21]), .ZN(n19) );
  INVX0 U43 ( .INP(in2[22]), .ZN(n20) );
  INVX0 U44 ( .INP(in1[1]), .ZN(n75) );
  INVX0 U45 ( .INP(in1[2]), .ZN(n72) );
  NOR2X0 U46 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n21) );
  OR3X1 U47 ( .IN1(in2[2]), .IN2(in2[0]), .IN3(in2[1]), .Q(n24) );
  OA21X1 U48 ( .IN1(n21), .IN2(n5), .IN3(n24), .Q(n25) );
  AOI22X1 U49 ( .IN1(in2[2]), .IN2(n90), .IN3(n92), .IN4(n25), .QN(n23) );
  NOR2X0 U50 ( .IN1(in2[3]), .IN2(n24), .QN(n26) );
  AOI21X1 U51 ( .IN1(in2[3]), .IN2(n24), .IN3(n26), .QN(n27) );
  AO222X1 U52 ( .IN1(in2[3]), .IN2(n90), .IN3(n92), .IN4(n27), .IN5(n89), 
        .IN6(n25), .Q(out1[3]) );
  OA21X1 U53 ( .IN1(n26), .IN2(n6), .IN3(n28), .Q(n29) );
  AO222X1 U54 ( .IN1(in2[4]), .IN2(n90), .IN3(n92), .IN4(n29), .IN5(n89), 
        .IN6(n27), .Q(out1[4]) );
  NOR2X0 U55 ( .IN1(in2[5]), .IN2(n28), .QN(n30) );
  AOI21X1 U56 ( .IN1(in2[5]), .IN2(n28), .IN3(n30), .QN(n31) );
  AO222X1 U57 ( .IN1(in2[5]), .IN2(n90), .IN3(n92), .IN4(n31), .IN5(n89), 
        .IN6(n29), .Q(out1[5]) );
  OA21X1 U58 ( .IN1(n30), .IN2(n7), .IN3(n32), .Q(n33) );
  AO222X1 U59 ( .IN1(in2[6]), .IN2(n90), .IN3(n92), .IN4(n33), .IN5(n89), 
        .IN6(n31), .Q(out1[6]) );
  NOR2X0 U60 ( .IN1(in2[7]), .IN2(n32), .QN(n34) );
  AOI21X1 U61 ( .IN1(in2[7]), .IN2(n32), .IN3(n34), .QN(n35) );
  AO222X1 U62 ( .IN1(in2[7]), .IN2(n90), .IN3(n92), .IN4(n35), .IN5(n89), 
        .IN6(n33), .Q(out1[7]) );
  OA21X1 U63 ( .IN1(n34), .IN2(n8), .IN3(n36), .Q(n37) );
  AO222X1 U64 ( .IN1(in2[8]), .IN2(n90), .IN3(n92), .IN4(n37), .IN5(n89), 
        .IN6(n35), .Q(out1[8]) );
  NOR2X0 U65 ( .IN1(in2[9]), .IN2(n36), .QN(n38) );
  AOI21X1 U66 ( .IN1(in2[9]), .IN2(n36), .IN3(n38), .QN(n39) );
  AO222X1 U67 ( .IN1(in2[9]), .IN2(n90), .IN3(n92), .IN4(n39), .IN5(n89), 
        .IN6(n37), .Q(out1[9]) );
  OA21X1 U68 ( .IN1(n38), .IN2(n9), .IN3(n40), .Q(n41) );
  AO222X1 U69 ( .IN1(in2[10]), .IN2(n90), .IN3(n92), .IN4(n41), .IN5(n89), 
        .IN6(n39), .Q(out1[10]) );
  NOR2X0 U70 ( .IN1(in2[11]), .IN2(n40), .QN(n42) );
  AOI21X1 U71 ( .IN1(in2[11]), .IN2(n40), .IN3(n42), .QN(n43) );
  AO222X1 U72 ( .IN1(in2[11]), .IN2(n90), .IN3(n92), .IN4(n43), .IN5(n89), 
        .IN6(n41), .Q(out1[11]) );
  OA21X1 U73 ( .IN1(n42), .IN2(n10), .IN3(n47), .Q(n45) );
  AO222X1 U74 ( .IN1(in2[12]), .IN2(n90), .IN3(n92), .IN4(n45), .IN5(n89), 
        .IN6(n43), .Q(out1[12]) );
  MUX21X1 U75 ( .IN1(n11), .IN2(in2[13]), .S(n44), .Q(n46) );
  AO22X1 U76 ( .IN1(in1[1]), .IN2(n46), .IN3(n89), .IN4(n45), .Q(out1[13]) );
  NOR2X0 U77 ( .IN1(in2[13]), .IN2(n47), .QN(n52) );
  AO21X1 U78 ( .IN1(in2[13]), .IN2(n47), .IN3(n86), .Q(n50) );
  NOR2X0 U79 ( .IN1(n52), .IN2(n72), .QN(n48) );
  MUX21X1 U80 ( .IN1(n12), .IN2(in2[14]), .S(n48), .Q(n49) );
  OAI22X1 U81 ( .IN1(n52), .IN2(n50), .IN3(n75), .IN4(n49), .QN(out1[14]) );
  MUX21X1 U82 ( .IN1(n13), .IN2(in2[15]), .S(n51), .Q(n54) );
  OA21X1 U83 ( .IN1(n52), .IN2(n12), .IN3(n89), .Q(n53) );
  AO22X1 U84 ( .IN1(in1[1]), .IN2(n54), .IN3(n53), .IN4(n55), .Q(out1[15]) );
  NOR2X0 U85 ( .IN1(in2[15]), .IN2(n55), .QN(n60) );
  AO21X1 U86 ( .IN1(in2[15]), .IN2(n55), .IN3(n86), .Q(n58) );
  NOR2X0 U87 ( .IN1(n60), .IN2(n72), .QN(n56) );
  MUX21X1 U88 ( .IN1(n14), .IN2(in2[16]), .S(n56), .Q(n57) );
  OAI22X1 U89 ( .IN1(n60), .IN2(n58), .IN3(n75), .IN4(n57), .QN(out1[16]) );
  MUX21X1 U90 ( .IN1(n15), .IN2(in2[17]), .S(n59), .Q(n62) );
  OA21X1 U91 ( .IN1(n60), .IN2(n14), .IN3(n89), .Q(n61) );
  AO22X1 U92 ( .IN1(in1[1]), .IN2(n62), .IN3(n61), .IN4(n63), .Q(out1[17]) );
  NOR2X0 U93 ( .IN1(in2[17]), .IN2(n63), .QN(n68) );
  AO21X1 U94 ( .IN1(in2[17]), .IN2(n63), .IN3(n86), .Q(n66) );
  NOR2X0 U95 ( .IN1(n68), .IN2(n72), .QN(n64) );
  MUX21X1 U96 ( .IN1(n16), .IN2(in2[18]), .S(n64), .Q(n65) );
  OAI22X1 U97 ( .IN1(n68), .IN2(n66), .IN3(n75), .IN4(n65), .QN(out1[18]) );
  MUX21X1 U98 ( .IN1(n17), .IN2(in2[19]), .S(n67), .Q(n70) );
  OA21X1 U99 ( .IN1(n68), .IN2(n16), .IN3(n89), .Q(n69) );
  AO22X1 U100 ( .IN1(in1[1]), .IN2(n70), .IN3(n69), .IN4(n71), .Q(out1[19]) );
  NOR2X0 U101 ( .IN1(in2[19]), .IN2(n71), .QN(n78) );
  AO21X1 U102 ( .IN1(in2[19]), .IN2(n71), .IN3(n86), .Q(n76) );
  NOR2X0 U103 ( .IN1(n78), .IN2(n72), .QN(n73) );
  MUX21X1 U104 ( .IN1(n18), .IN2(in2[20]), .S(n73), .Q(n74) );
  OAI22X1 U105 ( .IN1(n78), .IN2(n76), .IN3(n75), .IN4(n74), .QN(out1[20]) );
  MUX21X1 U106 ( .IN1(n19), .IN2(in2[21]), .S(n77), .Q(n80) );
  MUX21X1 U107 ( .IN1(n18), .IN2(in2[20]), .S(n78), .Q(n79) );
  AO22X1 U108 ( .IN1(in1[1]), .IN2(n80), .IN3(n89), .IN4(n79), .Q(out1[21]) );
  INVX0 U109 ( .INP(n92), .ZN(n81) );
  OR2X1 U110 ( .IN1(n82), .IN2(in2[21]), .Q(n88) );
  NOR2X0 U111 ( .IN1(n81), .IN2(n88), .QN(n87) );
  NOR2X0 U112 ( .IN1(in2[22]), .IN2(n81), .QN(n84) );
  OA221X1 U113 ( .IN1(n84), .IN2(n89), .IN3(n84), .IN4(n83), .IN5(n88), .Q(n85) );
  AO221X1 U114 ( .IN1(in2[22]), .IN2(n87), .IN3(in2[22]), .IN4(n90), .IN5(n85), 
        .Q(out1[22]) );
  NOR2X0 U115 ( .IN1(n86), .IN2(n88), .QN(n93) );
  AO21X1 U116 ( .IN1(n89), .IN2(n88), .IN3(n87), .Q(n91) );
  AO221X1 U117 ( .IN1(in2[22]), .IN2(n93), .IN3(n20), .IN4(n91), .IN5(n90), 
        .Q(out1[23]) );
  AO21X1 U118 ( .IN1(n93), .IN2(n20), .IN3(n92), .Q(out1[24]) );
endmodule


module mul26_6 ( clk, rst_n, in1, in2, en, mulout );
  input [25:0] in1;
  input [25:0] in2;
  output [50:0] mulout;
  input clk, rst_n, en;
  wire   N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24,
         N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38,
         N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N62, N63,
         N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77,
         N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91,
         N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n129, n130,
         SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22,
         SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24,
         SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26,
         SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28,
         SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30,
         SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32,
         SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34,
         SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36,
         SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38,
         SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40,
         SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42,
         SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44,
         SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46,
         SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48,
         SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50,
         SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52,
         SYNOPSYS_UNCONNECTED_53, SYNOPSYS_UNCONNECTED_54,
         SYNOPSYS_UNCONNECTED_55, SYNOPSYS_UNCONNECTED_56,
         SYNOPSYS_UNCONNECTED_57, SYNOPSYS_UNCONNECTED_58,
         SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_60,
         SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_62,
         SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_64,
         SYNOPSYS_UNCONNECTED_65, SYNOPSYS_UNCONNECTED_66,
         SYNOPSYS_UNCONNECTED_67, SYNOPSYS_UNCONNECTED_68,
         SYNOPSYS_UNCONNECTED_69, SYNOPSYS_UNCONNECTED_70,
         SYNOPSYS_UNCONNECTED_71, SYNOPSYS_UNCONNECTED_72,
         SYNOPSYS_UNCONNECTED_73, SYNOPSYS_UNCONNECTED_74,
         SYNOPSYS_UNCONNECTED_75, SYNOPSYS_UNCONNECTED_76,
         SYNOPSYS_UNCONNECTED_77, SYNOPSYS_UNCONNECTED_78,
         SYNOPSYS_UNCONNECTED_79, SYNOPSYS_UNCONNECTED_80,
         SYNOPSYS_UNCONNECTED_81, SYNOPSYS_UNCONNECTED_82,
         SYNOPSYS_UNCONNECTED_83, SYNOPSYS_UNCONNECTED_84,
         SYNOPSYS_UNCONNECTED_85, SYNOPSYS_UNCONNECTED_86,
         SYNOPSYS_UNCONNECTED_87, SYNOPSYS_UNCONNECTED_88,
         SYNOPSYS_UNCONNECTED_89, SYNOPSYS_UNCONNECTED_90,
         SYNOPSYS_UNCONNECTED_91, SYNOPSYS_UNCONNECTED_92,
         SYNOPSYS_UNCONNECTED_93, SYNOPSYS_UNCONNECTED_94,
         SYNOPSYS_UNCONNECTED_95, SYNOPSYS_UNCONNECTED_96,
         SYNOPSYS_UNCONNECTED_97, SYNOPSYS_UNCONNECTED_98,
         SYNOPSYS_UNCONNECTED_99, SYNOPSYS_UNCONNECTED_100,
         SYNOPSYS_UNCONNECTED_101, SYNOPSYS_UNCONNECTED_102,
         SYNOPSYS_UNCONNECTED_103, SYNOPSYS_UNCONNECTED_104,
         SYNOPSYS_UNCONNECTED_105, SYNOPSYS_UNCONNECTED_106,
         SYNOPSYS_UNCONNECTED_107, SYNOPSYS_UNCONNECTED_108,
         SYNOPSYS_UNCONNECTED_109, SYNOPSYS_UNCONNECTED_110,
         SYNOPSYS_UNCONNECTED_111, SYNOPSYS_UNCONNECTED_112,
         SYNOPSYS_UNCONNECTED_113, SYNOPSYS_UNCONNECTED_114,
         SYNOPSYS_UNCONNECTED_115, SYNOPSYS_UNCONNECTED_116,
         SYNOPSYS_UNCONNECTED_117, SYNOPSYS_UNCONNECTED_118,
         SYNOPSYS_UNCONNECTED_119, SYNOPSYS_UNCONNECTED_120,
         SYNOPSYS_UNCONNECTED_121, SYNOPSYS_UNCONNECTED_122,
         SYNOPSYS_UNCONNECTED_123, SYNOPSYS_UNCONNECTED_124,
         SYNOPSYS_UNCONNECTED_125, SYNOPSYS_UNCONNECTED_126,
         SYNOPSYS_UNCONNECTED_127, SYNOPSYS_UNCONNECTED_128,
         SYNOPSYS_UNCONNECTED_129, SYNOPSYS_UNCONNECTED_130,
         SYNOPSYS_UNCONNECTED_131, SYNOPSYS_UNCONNECTED_132,
         SYNOPSYS_UNCONNECTED_133, SYNOPSYS_UNCONNECTED_134,
         SYNOPSYS_UNCONNECTED_135, SYNOPSYS_UNCONNECTED_136,
         SYNOPSYS_UNCONNECTED_137, SYNOPSYS_UNCONNECTED_138,
         SYNOPSYS_UNCONNECTED_139, SYNOPSYS_UNCONNECTED_140,
         SYNOPSYS_UNCONNECTED_141, SYNOPSYS_UNCONNECTED_142,
         SYNOPSYS_UNCONNECTED_143, SYNOPSYS_UNCONNECTED_144,
         SYNOPSYS_UNCONNECTED_145, SYNOPSYS_UNCONNECTED_146,
         SYNOPSYS_UNCONNECTED_147, SYNOPSYS_UNCONNECTED_148,
         SYNOPSYS_UNCONNECTED_149, SYNOPSYS_UNCONNECTED_150,
         SYNOPSYS_UNCONNECTED_151, SYNOPSYS_UNCONNECTED_152,
         SYNOPSYS_UNCONNECTED_153, SYNOPSYS_UNCONNECTED_154,
         SYNOPSYS_UNCONNECTED_155, SYNOPSYS_UNCONNECTED_156,
         SYNOPSYS_UNCONNECTED_157, SYNOPSYS_UNCONNECTED_158,
         SYNOPSYS_UNCONNECTED_159, SYNOPSYS_UNCONNECTED_160,
         SYNOPSYS_UNCONNECTED_161, SYNOPSYS_UNCONNECTED_162,
         SYNOPSYS_UNCONNECTED_163, SYNOPSYS_UNCONNECTED_164,
         SYNOPSYS_UNCONNECTED_165, SYNOPSYS_UNCONNECTED_166,
         SYNOPSYS_UNCONNECTED_167, SYNOPSYS_UNCONNECTED_168,
         SYNOPSYS_UNCONNECTED_169, SYNOPSYS_UNCONNECTED_170,
         SYNOPSYS_UNCONNECTED_171, SYNOPSYS_UNCONNECTED_172,
         SYNOPSYS_UNCONNECTED_173, SYNOPSYS_UNCONNECTED_174,
         SYNOPSYS_UNCONNECTED_175, SYNOPSYS_UNCONNECTED_176,
         SYNOPSYS_UNCONNECTED_177, SYNOPSYS_UNCONNECTED_178,
         SYNOPSYS_UNCONNECTED_179, SYNOPSYS_UNCONNECTED_180,
         SYNOPSYS_UNCONNECTED_181, SYNOPSYS_UNCONNECTED_182,
         SYNOPSYS_UNCONNECTED_183, SYNOPSYS_UNCONNECTED_184,
         SYNOPSYS_UNCONNECTED_185, SYNOPSYS_UNCONNECTED_186,
         SYNOPSYS_UNCONNECTED_187, SYNOPSYS_UNCONNECTED_188,
         SYNOPSYS_UNCONNECTED_189, SYNOPSYS_UNCONNECTED_190,
         SYNOPSYS_UNCONNECTED_191, SYNOPSYS_UNCONNECTED_192,
         SYNOPSYS_UNCONNECTED_193, SYNOPSYS_UNCONNECTED_194,
         SYNOPSYS_UNCONNECTED_195, SYNOPSYS_UNCONNECTED_196,
         SYNOPSYS_UNCONNECTED_197, SYNOPSYS_UNCONNECTED_198,
         SYNOPSYS_UNCONNECTED_199, SYNOPSYS_UNCONNECTED_200,
         SYNOPSYS_UNCONNECTED_201, SYNOPSYS_UNCONNECTED_202,
         SYNOPSYS_UNCONNECTED_203, SYNOPSYS_UNCONNECTED_204,
         SYNOPSYS_UNCONNECTED_205, SYNOPSYS_UNCONNECTED_206,
         SYNOPSYS_UNCONNECTED_207, SYNOPSYS_UNCONNECTED_208,
         SYNOPSYS_UNCONNECTED_209, SYNOPSYS_UNCONNECTED_210,
         SYNOPSYS_UNCONNECTED_211, SYNOPSYS_UNCONNECTED_212,
         SYNOPSYS_UNCONNECTED_213, SYNOPSYS_UNCONNECTED_214,
         SYNOPSYS_UNCONNECTED_215, SYNOPSYS_UNCONNECTED_216,
         SYNOPSYS_UNCONNECTED_217, SYNOPSYS_UNCONNECTED_218,
         SYNOPSYS_UNCONNECTED_219, SYNOPSYS_UNCONNECTED_220,
         SYNOPSYS_UNCONNECTED_221, SYNOPSYS_UNCONNECTED_222,
         SYNOPSYS_UNCONNECTED_223, SYNOPSYS_UNCONNECTED_224,
         SYNOPSYS_UNCONNECTED_225, SYNOPSYS_UNCONNECTED_226,
         SYNOPSYS_UNCONNECTED_227, SYNOPSYS_UNCONNECTED_228,
         SYNOPSYS_UNCONNECTED_229, SYNOPSYS_UNCONNECTED_230,
         SYNOPSYS_UNCONNECTED_231, SYNOPSYS_UNCONNECTED_232,
         SYNOPSYS_UNCONNECTED_233, SYNOPSYS_UNCONNECTED_234,
         SYNOPSYS_UNCONNECTED_235, SYNOPSYS_UNCONNECTED_236,
         SYNOPSYS_UNCONNECTED_237, SYNOPSYS_UNCONNECTED_238,
         SYNOPSYS_UNCONNECTED_239, SYNOPSYS_UNCONNECTED_240,
         SYNOPSYS_UNCONNECTED_241, SYNOPSYS_UNCONNECTED_242,
         SYNOPSYS_UNCONNECTED_243, SYNOPSYS_UNCONNECTED_244,
         SYNOPSYS_UNCONNECTED_245, SYNOPSYS_UNCONNECTED_246,
         SYNOPSYS_UNCONNECTED_247, SYNOPSYS_UNCONNECTED_248,
         SYNOPSYS_UNCONNECTED_249, SYNOPSYS_UNCONNECTED_250,
         SYNOPSYS_UNCONNECTED_251, SYNOPSYS_UNCONNECTED_252,
         SYNOPSYS_UNCONNECTED_253, SYNOPSYS_UNCONNECTED_254,
         SYNOPSYS_UNCONNECTED_255, SYNOPSYS_UNCONNECTED_256,
         SYNOPSYS_UNCONNECTED_257, SYNOPSYS_UNCONNECTED_258,
         SYNOPSYS_UNCONNECTED_259, SYNOPSYS_UNCONNECTED_260,
         SYNOPSYS_UNCONNECTED_261, SYNOPSYS_UNCONNECTED_262,
         SYNOPSYS_UNCONNECTED_263, SYNOPSYS_UNCONNECTED_264,
         SYNOPSYS_UNCONNECTED_265, SYNOPSYS_UNCONNECTED_266,
         SYNOPSYS_UNCONNECTED_267, SYNOPSYS_UNCONNECTED_268,
         SYNOPSYS_UNCONNECTED_269, SYNOPSYS_UNCONNECTED_270,
         SYNOPSYS_UNCONNECTED_271, SYNOPSYS_UNCONNECTED_272,
         SYNOPSYS_UNCONNECTED_273, SYNOPSYS_UNCONNECTED_274,
         SYNOPSYS_UNCONNECTED_275, SYNOPSYS_UNCONNECTED_276,
         SYNOPSYS_UNCONNECTED_277, SYNOPSYS_UNCONNECTED_278,
         SYNOPSYS_UNCONNECTED_279, SYNOPSYS_UNCONNECTED_280,
         SYNOPSYS_UNCONNECTED_281, SYNOPSYS_UNCONNECTED_282,
         SYNOPSYS_UNCONNECTED_283, SYNOPSYS_UNCONNECTED_284,
         SYNOPSYS_UNCONNECTED_285, SYNOPSYS_UNCONNECTED_286,
         SYNOPSYS_UNCONNECTED_287, SYNOPSYS_UNCONNECTED_288,
         SYNOPSYS_UNCONNECTED_289, SYNOPSYS_UNCONNECTED_290,
         SYNOPSYS_UNCONNECTED_291, SYNOPSYS_UNCONNECTED_292,
         SYNOPSYS_UNCONNECTED_293, SYNOPSYS_UNCONNECTED_294,
         SYNOPSYS_UNCONNECTED_295, SYNOPSYS_UNCONNECTED_296,
         SYNOPSYS_UNCONNECTED_297, SYNOPSYS_UNCONNECTED_298,
         SYNOPSYS_UNCONNECTED_299, SYNOPSYS_UNCONNECTED_300,
         SYNOPSYS_UNCONNECTED_301, SYNOPSYS_UNCONNECTED_302,
         SYNOPSYS_UNCONNECTED_303, SYNOPSYS_UNCONNECTED_304,
         SYNOPSYS_UNCONNECTED_305, SYNOPSYS_UNCONNECTED_306,
         SYNOPSYS_UNCONNECTED_307, SYNOPSYS_UNCONNECTED_308,
         SYNOPSYS_UNCONNECTED_309, SYNOPSYS_UNCONNECTED_310,
         SYNOPSYS_UNCONNECTED_311, SYNOPSYS_UNCONNECTED_312,
         SYNOPSYS_UNCONNECTED_313, SYNOPSYS_UNCONNECTED_314,
         SYNOPSYS_UNCONNECTED_315, SYNOPSYS_UNCONNECTED_316,
         SYNOPSYS_UNCONNECTED_317, SYNOPSYS_UNCONNECTED_318,
         SYNOPSYS_UNCONNECTED_319, SYNOPSYS_UNCONNECTED_320,
         SYNOPSYS_UNCONNECTED_321, SYNOPSYS_UNCONNECTED_322,
         SYNOPSYS_UNCONNECTED_323, SYNOPSYS_UNCONNECTED_324,
         SYNOPSYS_UNCONNECTED_325, SYNOPSYS_UNCONNECTED_326,
         SYNOPSYS_UNCONNECTED_327, SYNOPSYS_UNCONNECTED_328,
         SYNOPSYS_UNCONNECTED_329, SYNOPSYS_UNCONNECTED_330,
         SYNOPSYS_UNCONNECTED_331, SYNOPSYS_UNCONNECTED_332,
         SYNOPSYS_UNCONNECTED_333, SYNOPSYS_UNCONNECTED_334,
         SYNOPSYS_UNCONNECTED_335, SYNOPSYS_UNCONNECTED_336,
         SYNOPSYS_UNCONNECTED_337, SYNOPSYS_UNCONNECTED_338,
         SYNOPSYS_UNCONNECTED_339, SYNOPSYS_UNCONNECTED_340,
         SYNOPSYS_UNCONNECTED_341, SYNOPSYS_UNCONNECTED_342,
         SYNOPSYS_UNCONNECTED_343, SYNOPSYS_UNCONNECTED_344,
         SYNOPSYS_UNCONNECTED_345, SYNOPSYS_UNCONNECTED_346,
         SYNOPSYS_UNCONNECTED_347, SYNOPSYS_UNCONNECTED_348,
         SYNOPSYS_UNCONNECTED_349, SYNOPSYS_UNCONNECTED_350,
         SYNOPSYS_UNCONNECTED_351, SYNOPSYS_UNCONNECTED_352,
         SYNOPSYS_UNCONNECTED_353, SYNOPSYS_UNCONNECTED_354,
         SYNOPSYS_UNCONNECTED_355, SYNOPSYS_UNCONNECTED_356,
         SYNOPSYS_UNCONNECTED_357, SYNOPSYS_UNCONNECTED_358,
         SYNOPSYS_UNCONNECTED_359, SYNOPSYS_UNCONNECTED_360,
         SYNOPSYS_UNCONNECTED_361, SYNOPSYS_UNCONNECTED_362,
         SYNOPSYS_UNCONNECTED_363, SYNOPSYS_UNCONNECTED_364,
         SYNOPSYS_UNCONNECTED_365, SYNOPSYS_UNCONNECTED_366,
         SYNOPSYS_UNCONNECTED_367, SYNOPSYS_UNCONNECTED_368,
         SYNOPSYS_UNCONNECTED_369, SYNOPSYS_UNCONNECTED_370,
         SYNOPSYS_UNCONNECTED_371, SYNOPSYS_UNCONNECTED_372,
         SYNOPSYS_UNCONNECTED_373, SYNOPSYS_UNCONNECTED_374,
         SYNOPSYS_UNCONNECTED_375, SYNOPSYS_UNCONNECTED_376,
         SYNOPSYS_UNCONNECTED_377, SYNOPSYS_UNCONNECTED_378,
         SYNOPSYS_UNCONNECTED_379, SYNOPSYS_UNCONNECTED_380,
         SYNOPSYS_UNCONNECTED_381, SYNOPSYS_UNCONNECTED_382,
         SYNOPSYS_UNCONNECTED_383, SYNOPSYS_UNCONNECTED_384,
         SYNOPSYS_UNCONNECTED_385, SYNOPSYS_UNCONNECTED_386,
         SYNOPSYS_UNCONNECTED_387, SYNOPSYS_UNCONNECTED_388,
         SYNOPSYS_UNCONNECTED_389, SYNOPSYS_UNCONNECTED_390,
         SYNOPSYS_UNCONNECTED_391, SYNOPSYS_UNCONNECTED_392,
         SYNOPSYS_UNCONNECTED_393, SYNOPSYS_UNCONNECTED_394,
         SYNOPSYS_UNCONNECTED_395, SYNOPSYS_UNCONNECTED_396,
         SYNOPSYS_UNCONNECTED_397, SYNOPSYS_UNCONNECTED_398,
         SYNOPSYS_UNCONNECTED_399, SYNOPSYS_UNCONNECTED_400,
         SYNOPSYS_UNCONNECTED_401, SYNOPSYS_UNCONNECTED_402,
         SYNOPSYS_UNCONNECTED_403, SYNOPSYS_UNCONNECTED_404,
         SYNOPSYS_UNCONNECTED_405, SYNOPSYS_UNCONNECTED_406,
         SYNOPSYS_UNCONNECTED_407, SYNOPSYS_UNCONNECTED_408,
         SYNOPSYS_UNCONNECTED_409, SYNOPSYS_UNCONNECTED_410,
         SYNOPSYS_UNCONNECTED_411, SYNOPSYS_UNCONNECTED_412,
         SYNOPSYS_UNCONNECTED_413, SYNOPSYS_UNCONNECTED_414;
  wire   [26:2] boothout1;
  wire   [26:0] boothout2;
  wire   [26:0] boothout3;
  wire   [26:0] boothout4;
  wire   [26:0] boothout5;
  wire   [26:0] boothout6;
  wire   [24:0] boothout7;
  wire   [26:0] boothout8;
  wire   [26:0] boothout9;
  wire   [26:0] boothout10;
  wire   [26:0] boothout11;
  wire   [25:0] boothout12;
  wire   [22:0] boothout13;
  wire   [29:2] cout1;
  wire   [31:3] mulout1;
  wire   [35:8] cout2;
  wire   [37:6] mulout2;
  wire   [41:14] cout3;
  wire   [42:12] mulout3;
  wire   [46:20] cout4;
  wire   [47:18] mulout4;
  wire   [31:3] cout5;
  wire   [46:4] mulout5;
  wire   [37:9] cout6;
  wire   [42:6] mulout6;
  wire   [46:18] cout7;
  wire   [47:12] mulout7;
  wire   [38:4] cout8;
  wire   [46:5] mulout8;
  wire   [46:12] cout9;
  wire   [47:6] mulout9;
  wire   [46:5] cout10;
  wire   [47:6] mulout10;
  wire   [46:6] cout11;
  wire   [47:7] mulout11;
  wire   [47:0] a;
  wire   [47:8] b;

  booth27_78 booth1 ( .out1({boothout1, SYNOPSYS_UNCONNECTED_1, 
        SYNOPSYS_UNCONNECTED_2}), .in1({in1[1:0], 1'b0}), .in2({1'b0, 1'b0, 
        1'b1, n30, n29, n28, n27, n26, n25, in2[16], n24, in2[14], n23, 
        in2[12], n22, in2[10], n21, in2[8], n20, in2[6], n19, in2[4:1], n18})
         );
  booth27_77 booth2 ( .out1(boothout2), .in1(in1[3:1]), .in2({1'b0, 1'b0, 1'b1, 
        n30, n29, n28, n27, n26, n25, in2[16], n24, in2[14], n23, in2[12], n22, 
        in2[10], n21, in2[8], n20, in2[6], n19, in2[4:1], n18}) );
  booth27_76 booth3 ( .out1(boothout3), .in1(in1[5:3]), .in2({1'b0, 1'b0, 1'b1, 
        n30, n29, n28, n27, n26, n25, in2[16], n24, in2[14], n23, in2[12], n22, 
        in2[10], n21, in2[8], n20, in2[6], n19, in2[4:1], n18}) );
  booth27_75 booth4 ( .out1(boothout4), .in1({in1[7], 1'b0, in1[5]}), .in2({
        1'b0, 1'b0, 1'b1, n30, n29, n28, n27, n26, n25, in2[16], n24, in2[14], 
        n23, in2[12], n22, in2[10], n21, in2[8], n20, in2[6], n19, in2[4:1], 
        n18}) );
  booth27_74 booth5 ( .out1(boothout5), .in1(in1[9:7]), .in2({1'b0, 1'b0, 1'b1, 
        n30, n29, n28, n27, n26, n25, in2[16], n24, in2[14], n23, in2[12], n22, 
        in2[10], n21, in2[8], n20, in2[6], n19, in2[4:1], n18}) );
  booth27_73 booth6 ( .out1(boothout6), .in1(in1[11:9]), .in2({1'b0, 1'b0, 
        1'b1, n30, n29, n28, n27, n26, n25, in2[16], n24, in2[14], n23, 
        in2[12], n22, in2[10], n21, in2[8], n20, in2[6], n19, in2[4:1], n18})
         );
  booth27_72 booth7 ( .out1({SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4, 
        boothout7}), .in1({1'b0, in1[12:11]}), .in2({1'b0, 1'b0, 1'b1, n30, 
        n29, n28, n27, n26, n25, in2[16], n24, in2[14], n23, in2[12], n22, 
        in2[10], n21, in2[8], n20, in2[6], n19, in2[4:1], n18}) );
  booth27_71 booth8 ( .out1(boothout8), .in1({in1[15:14], 1'b0}), .in2({1'b0, 
        1'b0, 1'b1, n30, n29, n28, n27, n26, n25, in2[16], n24, in2[14], n23, 
        in2[12], n22, in2[10], n21, in2[8], n20, in2[6], n19, in2[4:1], n18})
         );
  booth27_70 booth9 ( .out1(boothout9), .in1(in1[17:15]), .in2({1'b0, 1'b0, 
        1'b1, n30, n29, n28, n27, n26, n25, in2[16], n24, in2[14], n23, 
        in2[12], n22, in2[10], n21, in2[8], n20, in2[6], n19, in2[4:1], n18})
         );
  booth27_69 booth10 ( .out1(boothout10), .in1(in1[19:17]), .in2({1'b0, 1'b0, 
        1'b1, n30, n29, n28, n27, n26, n25, in2[16], n24, in2[14], n23, 
        in2[12], n22, in2[10], n21, in2[8], n20, in2[6], n19, in2[4:1], n18})
         );
  booth27_68 booth11 ( .out1(boothout11), .in1(in1[21:19]), .in2({1'b0, 1'b0, 
        1'b1, n30, n29, n28, n27, n26, n25, in2[16], n24, in2[14], n23, 
        in2[12], n22, in2[10], n21, in2[8], n20, in2[6], n19, in2[4:1], n18})
         );
  booth27_67 booth12 ( .out1({SYNOPSYS_UNCONNECTED_5, boothout12}), .in1({1'b1, 
        in1[22:21]}), .in2({1'b0, 1'b0, 1'b1, n30, n29, n28, n27, n26, n25, 
        in2[16], n24, in2[14], n23, in2[12], n22, in2[10], n21, in2[8], n20, 
        in2[6], n19, in2[4:1], n18}) );
  booth27_66 booth13 ( .out1({SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, 
        SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, boothout13}), .in1({
        1'b0, 1'b0, 1'b1}), .in2({1'b0, 1'b0, 1'b1, n30, n29, n28, n27, n26, 
        n25, in2[16], n24, in2[14], n23, in2[12], n22, in2[10], n21, in2[8], 
        n20, in2[6], n19, in2[4:1], n18}) );
  csa51squ_72 csa51squ1 ( .cout({SYNOPSYS_UNCONNECTED_10, 
        SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12, 
        SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14, 
        SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16, 
        SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18, 
        SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20, 
        SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22, 
        SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24, 
        SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26, 
        SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28, 
        SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30, cout1, 
        SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32}), .sumout({
        SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34, 
        SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36, 
        SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38, 
        SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40, 
        SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42, 
        SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44, 
        SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46, 
        SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48, 
        SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50, 
        SYNOPSYS_UNCONNECTED_51, mulout1[31], SYNOPSYS_UNCONNECTED_52, 
        mulout1[29:3], SYNOPSYS_UNCONNECTED_53, SYNOPSYS_UNCONNECTED_54, 
        SYNOPSYS_UNCONNECTED_55}), .in1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, boothout1, 1'b0, 1'b0}), .in2({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, boothout2, 
        1'b0, 1'b0}), .in3({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n130, 
        1'b0, boothout3[25:0], 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_71 csa51squ2 ( .cout({SYNOPSYS_UNCONNECTED_56, 
        SYNOPSYS_UNCONNECTED_57, SYNOPSYS_UNCONNECTED_58, 
        SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_60, 
        SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_62, 
        SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_64, 
        SYNOPSYS_UNCONNECTED_65, SYNOPSYS_UNCONNECTED_66, 
        SYNOPSYS_UNCONNECTED_67, SYNOPSYS_UNCONNECTED_68, 
        SYNOPSYS_UNCONNECTED_69, SYNOPSYS_UNCONNECTED_70, cout2, 
        SYNOPSYS_UNCONNECTED_71, SYNOPSYS_UNCONNECTED_72, 
        SYNOPSYS_UNCONNECTED_73, SYNOPSYS_UNCONNECTED_74, 
        SYNOPSYS_UNCONNECTED_75, SYNOPSYS_UNCONNECTED_76, 
        SYNOPSYS_UNCONNECTED_77, SYNOPSYS_UNCONNECTED_78}), .sumout({
        SYNOPSYS_UNCONNECTED_79, SYNOPSYS_UNCONNECTED_80, 
        SYNOPSYS_UNCONNECTED_81, SYNOPSYS_UNCONNECTED_82, 
        SYNOPSYS_UNCONNECTED_83, SYNOPSYS_UNCONNECTED_84, 
        SYNOPSYS_UNCONNECTED_85, SYNOPSYS_UNCONNECTED_86, 
        SYNOPSYS_UNCONNECTED_87, SYNOPSYS_UNCONNECTED_88, 
        SYNOPSYS_UNCONNECTED_89, SYNOPSYS_UNCONNECTED_90, 
        SYNOPSYS_UNCONNECTED_91, mulout2[37], SYNOPSYS_UNCONNECTED_92, 
        mulout2[35:6], SYNOPSYS_UNCONNECTED_93, SYNOPSYS_UNCONNECTED_94, 
        SYNOPSYS_UNCONNECTED_95, SYNOPSYS_UNCONNECTED_96, 
        SYNOPSYS_UNCONNECTED_97, SYNOPSYS_UNCONNECTED_98}), .in1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, boothout4, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, boothout5, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .in3({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n129, 1'b0, boothout6[25:0], 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_70 csa51squ3 ( .cout({SYNOPSYS_UNCONNECTED_99, 
        SYNOPSYS_UNCONNECTED_100, SYNOPSYS_UNCONNECTED_101, 
        SYNOPSYS_UNCONNECTED_102, SYNOPSYS_UNCONNECTED_103, 
        SYNOPSYS_UNCONNECTED_104, SYNOPSYS_UNCONNECTED_105, 
        SYNOPSYS_UNCONNECTED_106, SYNOPSYS_UNCONNECTED_107, cout3, 
        SYNOPSYS_UNCONNECTED_108, SYNOPSYS_UNCONNECTED_109, 
        SYNOPSYS_UNCONNECTED_110, SYNOPSYS_UNCONNECTED_111, 
        SYNOPSYS_UNCONNECTED_112, SYNOPSYS_UNCONNECTED_113, 
        SYNOPSYS_UNCONNECTED_114, SYNOPSYS_UNCONNECTED_115, 
        SYNOPSYS_UNCONNECTED_116, SYNOPSYS_UNCONNECTED_117, 
        SYNOPSYS_UNCONNECTED_118, SYNOPSYS_UNCONNECTED_119, 
        SYNOPSYS_UNCONNECTED_120, SYNOPSYS_UNCONNECTED_121}), .sumout({
        SYNOPSYS_UNCONNECTED_122, SYNOPSYS_UNCONNECTED_123, 
        SYNOPSYS_UNCONNECTED_124, SYNOPSYS_UNCONNECTED_125, 
        SYNOPSYS_UNCONNECTED_126, SYNOPSYS_UNCONNECTED_127, 
        SYNOPSYS_UNCONNECTED_128, SYNOPSYS_UNCONNECTED_129, mulout3, 
        SYNOPSYS_UNCONNECTED_130, SYNOPSYS_UNCONNECTED_131, 
        SYNOPSYS_UNCONNECTED_132, SYNOPSYS_UNCONNECTED_133, 
        SYNOPSYS_UNCONNECTED_134, SYNOPSYS_UNCONNECTED_135, 
        SYNOPSYS_UNCONNECTED_136, SYNOPSYS_UNCONNECTED_137, 
        SYNOPSYS_UNCONNECTED_138, SYNOPSYS_UNCONNECTED_139, 
        SYNOPSYS_UNCONNECTED_140, SYNOPSYS_UNCONNECTED_141}), .in1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 
        boothout7, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .in2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, boothout8, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in3({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, boothout9, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_69 csa51squ4 ( .cout({SYNOPSYS_UNCONNECTED_142, 
        SYNOPSYS_UNCONNECTED_143, SYNOPSYS_UNCONNECTED_144, 
        SYNOPSYS_UNCONNECTED_145, cout4, SYNOPSYS_UNCONNECTED_146, 
        SYNOPSYS_UNCONNECTED_147, SYNOPSYS_UNCONNECTED_148, 
        SYNOPSYS_UNCONNECTED_149, SYNOPSYS_UNCONNECTED_150, 
        SYNOPSYS_UNCONNECTED_151, SYNOPSYS_UNCONNECTED_152, 
        SYNOPSYS_UNCONNECTED_153, SYNOPSYS_UNCONNECTED_154, 
        SYNOPSYS_UNCONNECTED_155, SYNOPSYS_UNCONNECTED_156, 
        SYNOPSYS_UNCONNECTED_157, SYNOPSYS_UNCONNECTED_158, 
        SYNOPSYS_UNCONNECTED_159, SYNOPSYS_UNCONNECTED_160, 
        SYNOPSYS_UNCONNECTED_161, SYNOPSYS_UNCONNECTED_162, 
        SYNOPSYS_UNCONNECTED_163, SYNOPSYS_UNCONNECTED_164, 
        SYNOPSYS_UNCONNECTED_165}), .sumout({SYNOPSYS_UNCONNECTED_166, 
        SYNOPSYS_UNCONNECTED_167, SYNOPSYS_UNCONNECTED_168, mulout4, 
        SYNOPSYS_UNCONNECTED_169, SYNOPSYS_UNCONNECTED_170, 
        SYNOPSYS_UNCONNECTED_171, SYNOPSYS_UNCONNECTED_172, 
        SYNOPSYS_UNCONNECTED_173, SYNOPSYS_UNCONNECTED_174, 
        SYNOPSYS_UNCONNECTED_175, SYNOPSYS_UNCONNECTED_176, 
        SYNOPSYS_UNCONNECTED_177, SYNOPSYS_UNCONNECTED_178, 
        SYNOPSYS_UNCONNECTED_179, SYNOPSYS_UNCONNECTED_180, 
        SYNOPSYS_UNCONNECTED_181, SYNOPSYS_UNCONNECTED_182, 
        SYNOPSYS_UNCONNECTED_183, SYNOPSYS_UNCONNECTED_184, 
        SYNOPSYS_UNCONNECTED_185, SYNOPSYS_UNCONNECTED_186}), .in1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, boothout10, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 1'b0, 1'b0, 1'b0, boothout11, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .in3({1'b0, 1'b0, 1'b0, boothout12, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_68 csa51squ5 ( .cout({SYNOPSYS_UNCONNECTED_187, 
        SYNOPSYS_UNCONNECTED_188, SYNOPSYS_UNCONNECTED_189, 
        SYNOPSYS_UNCONNECTED_190, SYNOPSYS_UNCONNECTED_191, 
        SYNOPSYS_UNCONNECTED_192, SYNOPSYS_UNCONNECTED_193, 
        SYNOPSYS_UNCONNECTED_194, SYNOPSYS_UNCONNECTED_195, 
        SYNOPSYS_UNCONNECTED_196, SYNOPSYS_UNCONNECTED_197, 
        SYNOPSYS_UNCONNECTED_198, SYNOPSYS_UNCONNECTED_199, 
        SYNOPSYS_UNCONNECTED_200, SYNOPSYS_UNCONNECTED_201, 
        SYNOPSYS_UNCONNECTED_202, SYNOPSYS_UNCONNECTED_203, 
        SYNOPSYS_UNCONNECTED_204, SYNOPSYS_UNCONNECTED_205, cout5, 
        SYNOPSYS_UNCONNECTED_206, SYNOPSYS_UNCONNECTED_207, 
        SYNOPSYS_UNCONNECTED_208}), .sumout({SYNOPSYS_UNCONNECTED_209, 
        SYNOPSYS_UNCONNECTED_210, SYNOPSYS_UNCONNECTED_211, 
        SYNOPSYS_UNCONNECTED_212, mulout5, SYNOPSYS_UNCONNECTED_213, 
        SYNOPSYS_UNCONNECTED_214, SYNOPSYS_UNCONNECTED_215, 
        SYNOPSYS_UNCONNECTED_216}), .in1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, cout1, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, mulout1[31], 1'b0, mulout1[29:3], 1'b0, 1'b0, 1'b0}), 
        .in3({1'b0, 1'b0, 1'b0, 1'b1, boothout13, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_67 csa51squ6 ( .cout({SYNOPSYS_UNCONNECTED_217, 
        SYNOPSYS_UNCONNECTED_218, SYNOPSYS_UNCONNECTED_219, 
        SYNOPSYS_UNCONNECTED_220, SYNOPSYS_UNCONNECTED_221, 
        SYNOPSYS_UNCONNECTED_222, SYNOPSYS_UNCONNECTED_223, 
        SYNOPSYS_UNCONNECTED_224, SYNOPSYS_UNCONNECTED_225, 
        SYNOPSYS_UNCONNECTED_226, SYNOPSYS_UNCONNECTED_227, 
        SYNOPSYS_UNCONNECTED_228, SYNOPSYS_UNCONNECTED_229, cout6, 
        SYNOPSYS_UNCONNECTED_230, SYNOPSYS_UNCONNECTED_231, 
        SYNOPSYS_UNCONNECTED_232, SYNOPSYS_UNCONNECTED_233, 
        SYNOPSYS_UNCONNECTED_234, SYNOPSYS_UNCONNECTED_235, 
        SYNOPSYS_UNCONNECTED_236, SYNOPSYS_UNCONNECTED_237, 
        SYNOPSYS_UNCONNECTED_238}), .sumout({SYNOPSYS_UNCONNECTED_239, 
        SYNOPSYS_UNCONNECTED_240, SYNOPSYS_UNCONNECTED_241, 
        SYNOPSYS_UNCONNECTED_242, SYNOPSYS_UNCONNECTED_243, 
        SYNOPSYS_UNCONNECTED_244, SYNOPSYS_UNCONNECTED_245, 
        SYNOPSYS_UNCONNECTED_246, mulout6, SYNOPSYS_UNCONNECTED_247, 
        SYNOPSYS_UNCONNECTED_248, SYNOPSYS_UNCONNECTED_249, 
        SYNOPSYS_UNCONNECTED_250, SYNOPSYS_UNCONNECTED_251, 
        SYNOPSYS_UNCONNECTED_252}), .in1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, cout2, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        mulout2[37], 1'b0, mulout2[35:6], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .in3({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, cout3, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  csa51squ_66 csa51squ7 ( .cout({SYNOPSYS_UNCONNECTED_253, 
        SYNOPSYS_UNCONNECTED_254, SYNOPSYS_UNCONNECTED_255, 
        SYNOPSYS_UNCONNECTED_256, cout7, SYNOPSYS_UNCONNECTED_257, 
        SYNOPSYS_UNCONNECTED_258, SYNOPSYS_UNCONNECTED_259, 
        SYNOPSYS_UNCONNECTED_260, SYNOPSYS_UNCONNECTED_261, 
        SYNOPSYS_UNCONNECTED_262, SYNOPSYS_UNCONNECTED_263, 
        SYNOPSYS_UNCONNECTED_264, SYNOPSYS_UNCONNECTED_265, 
        SYNOPSYS_UNCONNECTED_266, SYNOPSYS_UNCONNECTED_267, 
        SYNOPSYS_UNCONNECTED_268, SYNOPSYS_UNCONNECTED_269, 
        SYNOPSYS_UNCONNECTED_270, SYNOPSYS_UNCONNECTED_271, 
        SYNOPSYS_UNCONNECTED_272, SYNOPSYS_UNCONNECTED_273, 
        SYNOPSYS_UNCONNECTED_274}), .sumout({SYNOPSYS_UNCONNECTED_275, 
        SYNOPSYS_UNCONNECTED_276, SYNOPSYS_UNCONNECTED_277, mulout7, 
        SYNOPSYS_UNCONNECTED_278, SYNOPSYS_UNCONNECTED_279, 
        SYNOPSYS_UNCONNECTED_280, SYNOPSYS_UNCONNECTED_281, 
        SYNOPSYS_UNCONNECTED_282, SYNOPSYS_UNCONNECTED_283, 
        SYNOPSYS_UNCONNECTED_284, SYNOPSYS_UNCONNECTED_285, 
        SYNOPSYS_UNCONNECTED_286, SYNOPSYS_UNCONNECTED_287, 
        SYNOPSYS_UNCONNECTED_288, SYNOPSYS_UNCONNECTED_289}), .in1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mulout3, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 1'b0, 
        1'b0, cout4, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in3({1'b0, 1'b0, 1'b0, mulout4, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_65 csa51squ8 ( .cout({SYNOPSYS_UNCONNECTED_290, 
        SYNOPSYS_UNCONNECTED_291, SYNOPSYS_UNCONNECTED_292, 
        SYNOPSYS_UNCONNECTED_293, SYNOPSYS_UNCONNECTED_294, 
        SYNOPSYS_UNCONNECTED_295, SYNOPSYS_UNCONNECTED_296, 
        SYNOPSYS_UNCONNECTED_297, SYNOPSYS_UNCONNECTED_298, 
        SYNOPSYS_UNCONNECTED_299, SYNOPSYS_UNCONNECTED_300, 
        SYNOPSYS_UNCONNECTED_301, cout8, SYNOPSYS_UNCONNECTED_302, 
        SYNOPSYS_UNCONNECTED_303, SYNOPSYS_UNCONNECTED_304, 
        SYNOPSYS_UNCONNECTED_305}), .sumout({SYNOPSYS_UNCONNECTED_306, 
        SYNOPSYS_UNCONNECTED_307, SYNOPSYS_UNCONNECTED_308, 
        SYNOPSYS_UNCONNECTED_309, mulout8, SYNOPSYS_UNCONNECTED_310, 
        SYNOPSYS_UNCONNECTED_311, SYNOPSYS_UNCONNECTED_312, 
        SYNOPSYS_UNCONNECTED_313, SYNOPSYS_UNCONNECTED_314}), .in1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, cout5, 1'b0, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 
        1'b0, 1'b0, 1'b1, mulout5, 1'b0, 1'b0, 1'b0, 1'b0}), .in3({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, cout6, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_64 csa51squ9 ( .cout({SYNOPSYS_UNCONNECTED_315, 
        SYNOPSYS_UNCONNECTED_316, SYNOPSYS_UNCONNECTED_317, 
        SYNOPSYS_UNCONNECTED_318, cout9, SYNOPSYS_UNCONNECTED_319, 
        SYNOPSYS_UNCONNECTED_320, SYNOPSYS_UNCONNECTED_321, 
        SYNOPSYS_UNCONNECTED_322, SYNOPSYS_UNCONNECTED_323, 
        SYNOPSYS_UNCONNECTED_324, SYNOPSYS_UNCONNECTED_325, 
        SYNOPSYS_UNCONNECTED_326, SYNOPSYS_UNCONNECTED_327, 
        SYNOPSYS_UNCONNECTED_328, SYNOPSYS_UNCONNECTED_329, 
        SYNOPSYS_UNCONNECTED_330}), .sumout({SYNOPSYS_UNCONNECTED_331, 
        SYNOPSYS_UNCONNECTED_332, SYNOPSYS_UNCONNECTED_333, mulout9, 
        SYNOPSYS_UNCONNECTED_334, SYNOPSYS_UNCONNECTED_335, 
        SYNOPSYS_UNCONNECTED_336, SYNOPSYS_UNCONNECTED_337, 
        SYNOPSYS_UNCONNECTED_338, SYNOPSYS_UNCONNECTED_339}), .in1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mulout6, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .in2({1'b0, 1'b0, 1'b0, cout7, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .in3({1'b0, 1'b0, 1'b0, mulout7, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_63 csa51squ10 ( .cout({SYNOPSYS_UNCONNECTED_340, 
        SYNOPSYS_UNCONNECTED_341, SYNOPSYS_UNCONNECTED_342, 
        SYNOPSYS_UNCONNECTED_343, cout10, SYNOPSYS_UNCONNECTED_344, 
        SYNOPSYS_UNCONNECTED_345, SYNOPSYS_UNCONNECTED_346, 
        SYNOPSYS_UNCONNECTED_347, SYNOPSYS_UNCONNECTED_348}), .sumout({
        SYNOPSYS_UNCONNECTED_349, SYNOPSYS_UNCONNECTED_350, 
        SYNOPSYS_UNCONNECTED_351, mulout10, SYNOPSYS_UNCONNECTED_352, 
        SYNOPSYS_UNCONNECTED_353, SYNOPSYS_UNCONNECTED_354, 
        SYNOPSYS_UNCONNECTED_355, SYNOPSYS_UNCONNECTED_356, 
        SYNOPSYS_UNCONNECTED_357}), .in1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, cout8, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .in2({1'b0, 1'b0, 1'b0, 1'b1, mulout8, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .in3({1'b0, 1'b0, 1'b0, cout9, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_62 csa51squ11 ( .cout({SYNOPSYS_UNCONNECTED_358, 
        SYNOPSYS_UNCONNECTED_359, SYNOPSYS_UNCONNECTED_360, 
        SYNOPSYS_UNCONNECTED_361, cout11, SYNOPSYS_UNCONNECTED_362, 
        SYNOPSYS_UNCONNECTED_363, SYNOPSYS_UNCONNECTED_364, 
        SYNOPSYS_UNCONNECTED_365, SYNOPSYS_UNCONNECTED_366, 
        SYNOPSYS_UNCONNECTED_367}), .sumout({SYNOPSYS_UNCONNECTED_368, 
        SYNOPSYS_UNCONNECTED_369, SYNOPSYS_UNCONNECTED_370, mulout11, 
        SYNOPSYS_UNCONNECTED_371, SYNOPSYS_UNCONNECTED_372, 
        SYNOPSYS_UNCONNECTED_373, SYNOPSYS_UNCONNECTED_374, 
        SYNOPSYS_UNCONNECTED_375, SYNOPSYS_UNCONNECTED_376, 
        SYNOPSYS_UNCONNECTED_377}), .in1({1'b0, 1'b0, 1'b0, mulout9, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 1'b0, 1'b0, cout10, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in3({1'b0, 1'b0, 1'b0, mulout10, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_61 csa51squ12 ( .sumout({SYNOPSYS_UNCONNECTED_378, 
        SYNOPSYS_UNCONNECTED_379, SYNOPSYS_UNCONNECTED_380, N101, N100, N99, 
        N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, 
        N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, 
        N70, N69, N68, N67, N66, N65, N64, N63, N62, SYNOPSYS_UNCONNECTED_381, 
        SYNOPSYS_UNCONNECTED_382, SYNOPSYS_UNCONNECTED_383, 
        SYNOPSYS_UNCONNECTED_384, SYNOPSYS_UNCONNECTED_385, 
        SYNOPSYS_UNCONNECTED_386, SYNOPSYS_UNCONNECTED_387, 
        SYNOPSYS_UNCONNECTED_388}), .in1({1'b0, 1'b0, 1'b0, mulout11, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 1'b0, 1'b0, cout11, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in3({1'b1, 1'b0, 1'b1, 
        1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 
        1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .cout_46_(N50), .cout_44_(N48), .cout_42_(N46), .cout_40_(N44), .cout_38_(
        N42), .cout_36_(N40), .cout_34_(N38), .cout_32_(N36), .cout_30_(N34), 
        .cout_28_(N32), .cout_27_(N31), .cout_7__BAR(N11), .cout_8__BAR(N12), 
        .cout_9__BAR(N13), .cout_10__BAR(N14), .cout_11__BAR(N15), 
        .cout_12__BAR(N16), .cout_13__BAR(N17), .cout_14__BAR(N18), 
        .cout_15__BAR(N19), .cout_16__BAR(N20), .cout_17__BAR(N21), 
        .cout_18__BAR(N22), .cout_19__BAR(N23), .cout_20__BAR(N24), 
        .cout_21__BAR(N25), .cout_22__BAR(N26), .cout_23__BAR(N27), 
        .cout_24__BAR(N28), .cout_25__BAR(N29), .cout_26__BAR(N30), 
        .cout_29__BAR(N33), .cout_31__BAR(N35), .cout_33__BAR(N37), 
        .cout_35__BAR(N39), .cout_37__BAR(N41), .cout_39__BAR(N43), 
        .cout_41__BAR(N45), .cout_43__BAR(N47), .cout_45__BAR(N49) );
  cla51squ_6 cla51squ ( .out({SYNOPSYS_UNCONNECTED_389, 
        SYNOPSYS_UNCONNECTED_390, SYNOPSYS_UNCONNECTED_391, mulout[47:23], 
        SYNOPSYS_UNCONNECTED_392, SYNOPSYS_UNCONNECTED_393, 
        SYNOPSYS_UNCONNECTED_394, SYNOPSYS_UNCONNECTED_395, 
        SYNOPSYS_UNCONNECTED_396, SYNOPSYS_UNCONNECTED_397, 
        SYNOPSYS_UNCONNECTED_398, SYNOPSYS_UNCONNECTED_399, 
        SYNOPSYS_UNCONNECTED_400, SYNOPSYS_UNCONNECTED_401, 
        SYNOPSYS_UNCONNECTED_402, SYNOPSYS_UNCONNECTED_403, 
        SYNOPSYS_UNCONNECTED_404, SYNOPSYS_UNCONNECTED_405, 
        SYNOPSYS_UNCONNECTED_406, SYNOPSYS_UNCONNECTED_407, 
        SYNOPSYS_UNCONNECTED_408, SYNOPSYS_UNCONNECTED_409, 
        SYNOPSYS_UNCONNECTED_410, SYNOPSYS_UNCONNECTED_411, 
        SYNOPSYS_UNCONNECTED_412, SYNOPSYS_UNCONNECTED_413, 
        SYNOPSYS_UNCONNECTED_414}), .a({1'b0, 1'b0, 1'b0, a[47:8], 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({1'b0, 1'b0, 1'b0, b, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  DFFARX1 b_reg_47_ ( .D(N101), .CLK(clk), .RSTB(rst_n), .Q(b[47]) );
  DFFARX1 b_reg_46_ ( .D(N100), .CLK(clk), .RSTB(rst_n), .Q(b[46]) );
  DFFARX1 b_reg_45_ ( .D(N99), .CLK(clk), .RSTB(rst_n), .Q(b[45]) );
  DFFARX1 b_reg_44_ ( .D(N98), .CLK(clk), .RSTB(rst_n), .Q(b[44]) );
  DFFARX1 b_reg_43_ ( .D(N97), .CLK(clk), .RSTB(rst_n), .Q(b[43]) );
  DFFARX1 b_reg_42_ ( .D(N96), .CLK(clk), .RSTB(rst_n), .Q(b[42]) );
  DFFARX1 b_reg_41_ ( .D(N95), .CLK(clk), .RSTB(rst_n), .Q(b[41]) );
  DFFARX1 b_reg_40_ ( .D(N94), .CLK(clk), .RSTB(rst_n), .Q(b[40]) );
  DFFARX1 b_reg_39_ ( .D(N93), .CLK(clk), .RSTB(rst_n), .Q(b[39]) );
  DFFARX1 b_reg_38_ ( .D(N92), .CLK(clk), .RSTB(rst_n), .Q(b[38]) );
  DFFARX1 b_reg_37_ ( .D(N91), .CLK(clk), .RSTB(rst_n), .Q(b[37]) );
  DFFARX1 b_reg_36_ ( .D(N90), .CLK(clk), .RSTB(rst_n), .Q(b[36]) );
  DFFARX1 b_reg_35_ ( .D(N89), .CLK(clk), .RSTB(rst_n), .Q(b[35]) );
  DFFARX1 b_reg_34_ ( .D(N88), .CLK(clk), .RSTB(rst_n), .Q(b[34]) );
  DFFARX1 b_reg_33_ ( .D(N87), .CLK(clk), .RSTB(rst_n), .Q(b[33]) );
  DFFARX1 b_reg_32_ ( .D(N86), .CLK(clk), .RSTB(rst_n), .Q(b[32]) );
  DFFARX1 b_reg_31_ ( .D(N85), .CLK(clk), .RSTB(rst_n), .Q(b[31]) );
  DFFARX1 b_reg_30_ ( .D(N84), .CLK(clk), .RSTB(rst_n), .Q(b[30]) );
  DFFARX1 b_reg_29_ ( .D(N83), .CLK(clk), .RSTB(rst_n), .Q(b[29]) );
  DFFARX1 b_reg_28_ ( .D(N82), .CLK(clk), .RSTB(rst_n), .Q(b[28]) );
  DFFARX1 b_reg_27_ ( .D(N81), .CLK(clk), .RSTB(rst_n), .Q(b[27]) );
  DFFARX1 b_reg_26_ ( .D(N80), .CLK(clk), .RSTB(rst_n), .Q(b[26]) );
  DFFARX1 b_reg_25_ ( .D(N79), .CLK(clk), .RSTB(rst_n), .Q(b[25]) );
  DFFARX1 b_reg_24_ ( .D(N78), .CLK(clk), .RSTB(rst_n), .Q(b[24]) );
  DFFARX1 b_reg_23_ ( .D(N77), .CLK(clk), .RSTB(rst_n), .Q(b[23]) );
  DFFARX1 b_reg_22_ ( .D(N76), .CLK(clk), .RSTB(rst_n), .Q(b[22]) );
  DFFARX1 b_reg_21_ ( .D(N75), .CLK(clk), .RSTB(rst_n), .Q(b[21]) );
  DFFARX1 b_reg_20_ ( .D(N74), .CLK(clk), .RSTB(rst_n), .Q(b[20]) );
  DFFARX1 b_reg_19_ ( .D(N73), .CLK(clk), .RSTB(rst_n), .Q(b[19]) );
  DFFARX1 b_reg_18_ ( .D(N72), .CLK(clk), .RSTB(rst_n), .Q(b[18]) );
  DFFARX1 b_reg_17_ ( .D(N71), .CLK(clk), .RSTB(rst_n), .Q(b[17]) );
  DFFARX1 b_reg_16_ ( .D(N70), .CLK(clk), .RSTB(rst_n), .Q(b[16]) );
  DFFARX1 b_reg_15_ ( .D(N69), .CLK(clk), .RSTB(rst_n), .Q(b[15]) );
  DFFARX1 b_reg_14_ ( .D(N68), .CLK(clk), .RSTB(rst_n), .Q(b[14]) );
  DFFARX1 b_reg_13_ ( .D(N67), .CLK(clk), .RSTB(rst_n), .Q(b[13]) );
  DFFARX1 b_reg_12_ ( .D(N66), .CLK(clk), .RSTB(rst_n), .Q(b[12]) );
  DFFARX1 b_reg_11_ ( .D(N65), .CLK(clk), .RSTB(rst_n), .Q(b[11]) );
  DFFARX1 b_reg_10_ ( .D(N64), .CLK(clk), .RSTB(rst_n), .Q(b[10]) );
  DFFARX1 b_reg_9_ ( .D(N63), .CLK(clk), .RSTB(rst_n), .Q(b[9]) );
  DFFARX1 b_reg_8_ ( .D(N62), .CLK(clk), .RSTB(rst_n), .Q(b[8]) );
  DFFARX1 a_reg_47_ ( .D(N50), .CLK(clk), .RSTB(rst_n), .Q(a[47]) );
  DFFARX1 a_reg_46_ ( .D(n60), .CLK(clk), .RSTB(rst_n), .Q(a[46]) );
  DFFARX1 a_reg_45_ ( .D(N48), .CLK(clk), .RSTB(rst_n), .Q(a[45]) );
  DFFARX1 a_reg_44_ ( .D(n61), .CLK(clk), .RSTB(rst_n), .Q(a[44]) );
  DFFARX1 a_reg_43_ ( .D(N46), .CLK(clk), .RSTB(rst_n), .Q(a[43]) );
  DFFARX1 a_reg_42_ ( .D(n62), .CLK(clk), .RSTB(rst_n), .Q(a[42]) );
  DFFARX1 a_reg_41_ ( .D(N44), .CLK(clk), .RSTB(rst_n), .Q(a[41]) );
  DFFARX1 a_reg_40_ ( .D(n63), .CLK(clk), .RSTB(rst_n), .Q(a[40]) );
  DFFARX1 a_reg_39_ ( .D(N42), .CLK(clk), .RSTB(rst_n), .Q(a[39]) );
  DFFARX1 a_reg_38_ ( .D(n64), .CLK(clk), .RSTB(rst_n), .Q(a[38]) );
  DFFARX1 a_reg_37_ ( .D(N40), .CLK(clk), .RSTB(rst_n), .Q(a[37]) );
  DFFARX1 a_reg_36_ ( .D(n65), .CLK(clk), .RSTB(rst_n), .Q(a[36]) );
  DFFARX1 a_reg_35_ ( .D(N38), .CLK(clk), .RSTB(rst_n), .Q(a[35]) );
  DFFARX1 a_reg_34_ ( .D(n66), .CLK(clk), .RSTB(rst_n), .Q(a[34]) );
  DFFARX1 a_reg_33_ ( .D(N36), .CLK(clk), .RSTB(rst_n), .Q(a[33]) );
  DFFARX1 a_reg_32_ ( .D(n67), .CLK(clk), .RSTB(rst_n), .Q(a[32]) );
  DFFARX1 a_reg_31_ ( .D(N34), .CLK(clk), .RSTB(rst_n), .Q(a[31]) );
  DFFARX1 a_reg_30_ ( .D(n68), .CLK(clk), .RSTB(rst_n), .Q(a[30]) );
  DFFARX1 a_reg_29_ ( .D(N32), .CLK(clk), .RSTB(rst_n), .Q(a[29]) );
  DFFARX1 a_reg_28_ ( .D(N31), .CLK(clk), .RSTB(rst_n), .Q(a[28]) );
  DFFARX1 a_reg_27_ ( .D(n69), .CLK(clk), .RSTB(rst_n), .Q(a[27]) );
  DFFARX1 a_reg_26_ ( .D(n70), .CLK(clk), .RSTB(rst_n), .Q(a[26]) );
  DFFARX1 a_reg_25_ ( .D(n71), .CLK(clk), .RSTB(rst_n), .Q(a[25]) );
  DFFARX1 a_reg_24_ ( .D(n72), .CLK(clk), .RSTB(rst_n), .Q(a[24]) );
  DFFARX1 a_reg_23_ ( .D(n73), .CLK(clk), .RSTB(rst_n), .Q(a[23]) );
  DFFARX1 a_reg_22_ ( .D(n74), .CLK(clk), .RSTB(rst_n), .Q(a[22]) );
  DFFARX1 a_reg_21_ ( .D(n75), .CLK(clk), .RSTB(rst_n), .Q(a[21]) );
  DFFARX1 a_reg_20_ ( .D(n76), .CLK(clk), .RSTB(rst_n), .Q(a[20]) );
  DFFARX1 a_reg_19_ ( .D(n77), .CLK(clk), .RSTB(rst_n), .Q(a[19]) );
  DFFARX1 a_reg_18_ ( .D(n78), .CLK(clk), .RSTB(rst_n), .Q(a[18]) );
  DFFARX1 a_reg_17_ ( .D(n79), .CLK(clk), .RSTB(rst_n), .Q(a[17]) );
  DFFARX1 a_reg_16_ ( .D(n80), .CLK(clk), .RSTB(rst_n), .Q(a[16]) );
  DFFARX1 a_reg_15_ ( .D(n81), .CLK(clk), .RSTB(rst_n), .Q(a[15]) );
  DFFARX1 a_reg_14_ ( .D(n82), .CLK(clk), .RSTB(rst_n), .Q(a[14]) );
  DFFARX1 a_reg_13_ ( .D(n83), .CLK(clk), .RSTB(rst_n), .Q(a[13]) );
  DFFARX1 a_reg_12_ ( .D(n84), .CLK(clk), .RSTB(rst_n), .Q(a[12]) );
  DFFARX1 a_reg_11_ ( .D(n85), .CLK(clk), .RSTB(rst_n), .Q(a[11]) );
  DFFARX1 a_reg_10_ ( .D(n86), .CLK(clk), .RSTB(rst_n), .Q(a[10]) );
  DFFARX1 a_reg_9_ ( .D(n87), .CLK(clk), .RSTB(rst_n), .Q(a[9]) );
  DFFARX1 a_reg_8_ ( .D(n88), .CLK(clk), .RSTB(rst_n), .Q(a[8]) );
  INVX0 U5 ( .INP(boothout3[26]), .ZN(n130) );
  INVX0 U8 ( .INP(boothout6[26]), .ZN(n129) );
  NBUFFX8 U3 ( .INP(in2[18]), .Z(n26) );
  NBUFFX8 U4 ( .INP(in2[20]), .Z(n28) );
  NBUFFX8 U6 ( .INP(in2[11]), .Z(n22) );
  NBUFFX8 U7 ( .INP(in2[5]), .Z(n19) );
  NBUFFX8 U9 ( .INP(in2[9]), .Z(n21) );
  NBUFFX8 U10 ( .INP(in2[7]), .Z(n20) );
  NBUFFX8 U11 ( .INP(in2[19]), .Z(n27) );
  NBUFFX8 U12 ( .INP(in2[17]), .Z(n25) );
  NBUFFX8 U13 ( .INP(in2[15]), .Z(n24) );
  NBUFFX8 U14 ( .INP(in2[13]), .Z(n23) );
  NBUFFX8 U15 ( .INP(in2[21]), .Z(n29) );
  NBUFFX8 U16 ( .INP(in2[22]), .Z(n30) );
  NBUFFX8 U17 ( .INP(in2[0]), .Z(n18) );
  INVX0 U69 ( .INP(N49), .ZN(n60) );
  INVX0 U70 ( .INP(N47), .ZN(n61) );
  INVX0 U71 ( .INP(N45), .ZN(n62) );
  INVX0 U72 ( .INP(N43), .ZN(n63) );
  INVX0 U73 ( .INP(N41), .ZN(n64) );
  INVX0 U74 ( .INP(N39), .ZN(n65) );
  INVX0 U75 ( .INP(N37), .ZN(n66) );
  INVX0 U76 ( .INP(N35), .ZN(n67) );
  INVX0 U77 ( .INP(N33), .ZN(n68) );
  INVX0 U78 ( .INP(N30), .ZN(n69) );
  INVX0 U79 ( .INP(N29), .ZN(n70) );
  INVX0 U80 ( .INP(N28), .ZN(n71) );
  INVX0 U81 ( .INP(N27), .ZN(n72) );
  INVX0 U82 ( .INP(N26), .ZN(n73) );
  INVX0 U83 ( .INP(N25), .ZN(n74) );
  INVX0 U84 ( .INP(N24), .ZN(n75) );
  INVX0 U85 ( .INP(N23), .ZN(n76) );
  INVX0 U86 ( .INP(N22), .ZN(n77) );
  INVX0 U87 ( .INP(N21), .ZN(n78) );
  INVX0 U88 ( .INP(N20), .ZN(n79) );
  INVX0 U89 ( .INP(N19), .ZN(n80) );
  INVX0 U90 ( .INP(N18), .ZN(n81) );
  INVX0 U91 ( .INP(N17), .ZN(n82) );
  INVX0 U92 ( .INP(N16), .ZN(n83) );
  INVX0 U93 ( .INP(N15), .ZN(n84) );
  INVX0 U94 ( .INP(N14), .ZN(n85) );
  INVX0 U95 ( .INP(N13), .ZN(n86) );
  INVX0 U96 ( .INP(N12), .ZN(n87) );
  INVX0 U97 ( .INP(N11), .ZN(n88) );
endmodule


module add_657 ( s, a, b, co, ci_BAR );
  input a, b, ci_BAR;
  output s, co;


  XOR2X1 U1 ( .IN1(a), .IN2(ci_BAR), .Q(s) );
endmodule


module add_658 ( s, a, b, ci, co_BAR );
  input a, b, ci;
  output s, co_BAR;


  NAND2X0 U1 ( .IN1(ci), .IN2(a), .QN(co_BAR) );
  OA21X1 U2 ( .IN1(ci), .IN2(a), .IN3(co_BAR), .Q(s) );
endmodule


module add_659 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_660 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_661 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_662 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_663 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  INVX0 U1 ( .INP(a), .ZN(s) );
  NBUFFX2 U2 ( .INP(a), .Z(co) );
endmodule


module add_664 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  NBUFFX2 U1 ( .INP(a), .Z(s) );
endmodule


module adder8_47 ( out, a, b, cin );
  output [7:0] out;
  input [7:0] a;
  input [7:0] b;
  input cin;

  wire   [6:1] c;

  add_664 add_01 ( .s(out[0]), .a(a[0]), .b(1'b1), .ci(1'b1) );
  add_663 add_02 ( .s(out[1]), .a(a[1]), .b(1'b0), .ci(1'b1), .co(c[1]) );
  add_662 add_03 ( .s(out[2]), .a(a[2]), .b(1'b0), .ci(c[1]), .co(c[2]) );
  add_661 add_04 ( .s(out[3]), .a(a[3]), .b(1'b0), .ci(c[2]), .co(c[3]) );
  add_660 add_05 ( .s(out[4]), .a(a[4]), .b(1'b0), .ci(c[3]), .co(c[4]) );
  add_659 add_06 ( .s(out[5]), .a(a[5]), .b(1'b0), .ci(c[4]), .co(c[5]) );
  add_658 add_07 ( .s(out[6]), .a(a[6]), .b(1'b0), .ci(c[5]), .co_BAR(c[6]) );
  add_657 add_08 ( .s(out[7]), .a(a[7]), .b(1'b1), .ci_BAR(c[6]) );
endmodule


module add_665 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  XOR2X1 U1 ( .IN1(ci), .IN2(b), .Q(s) );
endmodule


module add_666 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_667 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_668 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_669 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_670 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_671 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_672 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(b), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(b), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module adder8_48 ( out, a, b, cin );
  output [7:0] out;
  input [7:0] a;
  input [7:0] b;
  input cin;

  wire   [6:0] c;

  add_672 add_01 ( .s(out[0]), .a(a[0]), .b(b[0]), .ci(1'b0), .co(c[0]) );
  add_671 add_02 ( .s(out[1]), .a(a[1]), .b(b[1]), .ci(c[0]), .co(c[1]) );
  add_670 add_03 ( .s(out[2]), .a(a[2]), .b(b[2]), .ci(c[1]), .co(c[2]) );
  add_669 add_04 ( .s(out[3]), .a(a[3]), .b(b[3]), .ci(c[2]), .co(c[3]) );
  add_668 add_05 ( .s(out[4]), .a(a[4]), .b(b[4]), .ci(c[3]), .co(c[4]) );
  add_667 add_06 ( .s(out[5]), .a(a[5]), .b(b[5]), .ci(c[4]), .co(c[5]) );
  add_666 add_07 ( .s(out[6]), .a(a[6]), .b(b[6]), .ci(c[5]), .co(c[6]) );
  add_665 add_08 ( .s(out[7]), .a(1'b0), .b(b[7]), .ci(c[6]) );
endmodule


module floating_point_multiple_6 ( clk, rst_n, input_factor_01, 
        input_factor_02, output_multiply );
  input [31:0] input_factor_01;
  input [31:0] input_factor_02;
  output [31:0] output_multiply;
  input clk, rst_n;
  wire   N5, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22,
         N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N48, N49, N50, N51,
         N52, N53, N54, N55, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22,
         SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24,
         SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26;
  wire   [47:23] base_multiply_result;
  wire   [47:23] mulout;
  wire   [7:0] exponent_factor_12;
  wire   [7:0] pre_mul_output_exponent;

  mul26_6 mul26_01 ( .clk(clk), .rst_n(rst_n), .in1({1'b0, 1'b0, 1'b1, 
        input_factor_01[22:14], 1'b0, input_factor_01[12:7], 1'b0, 
        input_factor_01[5:0]}), .in2({1'b0, 1'b0, 1'b1, input_factor_02[22:0]}), .en(1'b1), .mulout({SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, 
        SYNOPSYS_UNCONNECTED_3, mulout, SYNOPSYS_UNCONNECTED_4, 
        SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, 
        SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, 
        SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11, 
        SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13, 
        SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, 
        SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17, 
        SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19, 
        SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21, 
        SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_23, 
        SYNOPSYS_UNCONNECTED_24, SYNOPSYS_UNCONNECTED_25, 
        SYNOPSYS_UNCONNECTED_26}) );
  adder8_48 adder8_01 ( .out(exponent_factor_12), .a({1'b0, 
        input_factor_01[29:23]}), .b(input_factor_02[30:23]), .cin(1'b0) );
  adder8_47 adder8_02 ( .out(pre_mul_output_exponent), .a(exponent_factor_12), 
        .b({1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0}), .cin(1'b1) );
  DFFARX1 mul_output_sign_reg ( .D(N5), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[31]) );
  DFFARX1 base_multiply_result_reg_47_ ( .D(mulout[47]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[47]) );
  DFFARX1 base_multiply_result_reg_46_ ( .D(mulout[46]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[46]) );
  DFFARX1 base_multiply_result_reg_45_ ( .D(mulout[45]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[45]) );
  DFFARX1 base_multiply_result_reg_44_ ( .D(mulout[44]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[44]) );
  DFFARX1 base_multiply_result_reg_43_ ( .D(mulout[43]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[43]) );
  DFFARX1 base_multiply_result_reg_42_ ( .D(mulout[42]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[42]) );
  DFFARX1 base_multiply_result_reg_41_ ( .D(mulout[41]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[41]) );
  DFFARX1 base_multiply_result_reg_40_ ( .D(mulout[40]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[40]) );
  DFFARX1 base_multiply_result_reg_39_ ( .D(mulout[39]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[39]) );
  DFFARX1 base_multiply_result_reg_38_ ( .D(mulout[38]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[38]) );
  DFFARX1 base_multiply_result_reg_37_ ( .D(mulout[37]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[37]) );
  DFFARX1 base_multiply_result_reg_36_ ( .D(mulout[36]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[36]) );
  DFFARX1 base_multiply_result_reg_35_ ( .D(mulout[35]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[35]) );
  DFFARX1 base_multiply_result_reg_34_ ( .D(mulout[34]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[34]) );
  DFFARX1 base_multiply_result_reg_33_ ( .D(mulout[33]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[33]) );
  DFFARX1 base_multiply_result_reg_32_ ( .D(mulout[32]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[32]) );
  DFFARX1 base_multiply_result_reg_31_ ( .D(mulout[31]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[31]) );
  DFFARX1 base_multiply_result_reg_30_ ( .D(mulout[30]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[30]) );
  DFFARX1 base_multiply_result_reg_29_ ( .D(mulout[29]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[29]) );
  DFFARX1 base_multiply_result_reg_28_ ( .D(mulout[28]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[28]) );
  DFFARX1 base_multiply_result_reg_27_ ( .D(mulout[27]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[27]) );
  DFFARX1 base_multiply_result_reg_26_ ( .D(mulout[26]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[26]) );
  DFFARX1 base_multiply_result_reg_25_ ( .D(mulout[25]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[25]) );
  DFFARX1 base_multiply_result_reg_24_ ( .D(mulout[24]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[24]) );
  DFFARX1 base_multiply_result_reg_23_ ( .D(mulout[23]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[23]) );
  DFFARX1 mul_output_significand_reg_22_ ( .D(N32), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[22]) );
  DFFARX1 mul_output_significand_reg_21_ ( .D(N31), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[21]) );
  DFFARX1 mul_output_significand_reg_20_ ( .D(N30), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[20]) );
  DFFARX1 mul_output_significand_reg_19_ ( .D(N29), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[19]) );
  DFFARX1 mul_output_significand_reg_18_ ( .D(N28), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[18]) );
  DFFARX1 mul_output_significand_reg_17_ ( .D(N27), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[17]) );
  DFFARX1 mul_output_significand_reg_16_ ( .D(N26), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[16]) );
  DFFARX1 mul_output_significand_reg_15_ ( .D(N25), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[15]) );
  DFFARX1 mul_output_significand_reg_14_ ( .D(N24), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[14]) );
  DFFARX1 mul_output_significand_reg_13_ ( .D(N23), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[13]) );
  DFFARX1 mul_output_significand_reg_12_ ( .D(N22), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[12]) );
  DFFARX1 mul_output_significand_reg_11_ ( .D(N21), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[11]) );
  DFFARX1 mul_output_significand_reg_10_ ( .D(N20), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[10]) );
  DFFARX1 mul_output_significand_reg_9_ ( .D(N19), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[9]) );
  DFFARX1 mul_output_significand_reg_8_ ( .D(N18), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[8]) );
  DFFARX1 mul_output_significand_reg_7_ ( .D(N17), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[7]) );
  DFFARX1 mul_output_significand_reg_6_ ( .D(N16), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[6]) );
  DFFARX1 mul_output_significand_reg_5_ ( .D(N15), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[5]) );
  DFFARX1 mul_output_significand_reg_4_ ( .D(N14), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[4]) );
  DFFARX1 mul_output_significand_reg_3_ ( .D(N13), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[3]) );
  DFFARX1 mul_output_significand_reg_2_ ( .D(N12), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[2]) );
  DFFARX1 mul_output_significand_reg_1_ ( .D(N11), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[1]) );
  DFFARX1 mul_output_significand_reg_0_ ( .D(N10), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[0]) );
  DFFARX1 mul_output_exponent_reg_7_ ( .D(N55), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[30]) );
  DFFARX1 mul_output_exponent_reg_6_ ( .D(N54), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[29]) );
  DFFARX1 mul_output_exponent_reg_5_ ( .D(N53), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[28]) );
  DFFARX1 mul_output_exponent_reg_4_ ( .D(N52), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[27]) );
  DFFARX1 mul_output_exponent_reg_3_ ( .D(N51), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[26]) );
  DFFARX1 mul_output_exponent_reg_2_ ( .D(N50), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[25]) );
  DFFARX1 mul_output_exponent_reg_1_ ( .D(N49), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[24]) );
  DFFARX1 mul_output_exponent_reg_0_ ( .D(N48), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[23]) );
  AND2X1 U3 ( .IN1(base_multiply_result[47]), .IN2(n35), .Q(n32) );
  INVX0 U4 ( .INP(n1), .ZN(n2) );
  OR2X1 U5 ( .IN1(base_multiply_result[47]), .IN2(n24), .Q(n1) );
  INVX0 U6 ( .INP(input_factor_02[31]), .ZN(n3) );
  NOR4X0 U8 ( .IN1(input_factor_01[21]), .IN2(input_factor_01[23]), .IN3(
        input_factor_01[17]), .IN4(input_factor_01[18]), .QN(n7) );
  NOR4X0 U9 ( .IN1(input_factor_01[11]), .IN2(input_factor_01[12]), .IN3(
        input_factor_01[22]), .IN4(input_factor_01[20]), .QN(n6) );
  NOR4X0 U10 ( .IN1(input_factor_01[28]), .IN2(input_factor_01[15]), .IN3(
        input_factor_01[16]), .IN4(input_factor_01[14]), .QN(n5) );
  NOR4X0 U11 ( .IN1(input_factor_01[19]), .IN2(input_factor_01[2]), .IN3(
        input_factor_01[1]), .IN4(input_factor_01[29]), .QN(n4) );
  NAND4X0 U12 ( .IN1(n7), .IN2(n6), .IN3(n5), .IN4(n4), .QN(n23) );
  NOR4X0 U13 ( .IN1(input_factor_01[8]), .IN2(input_factor_01[9]), .IN3(
        input_factor_01[24]), .IN4(input_factor_01[25]), .QN(n11) );
  NOR4X0 U14 ( .IN1(input_factor_01[4]), .IN2(input_factor_01[5]), .IN3(
        input_factor_01[0]), .IN4(input_factor_01[10]), .QN(n10) );
  NOR4X0 U15 ( .IN1(input_factor_01[26]), .IN2(input_factor_01[27]), .IN3(
        input_factor_01[31]), .IN4(input_factor_01[3]), .QN(n9) );
  INVX0 U16 ( .INP(input_factor_01[7]), .ZN(n8) );
  NAND4X0 U17 ( .IN1(n11), .IN2(n10), .IN3(n9), .IN4(n8), .QN(n22) );
  NOR4X0 U18 ( .IN1(input_factor_02[0]), .IN2(input_factor_02[10]), .IN3(
        input_factor_02[11]), .IN4(input_factor_02[12]), .QN(n15) );
  NOR4X0 U19 ( .IN1(input_factor_02[13]), .IN2(input_factor_02[14]), .IN3(
        input_factor_02[15]), .IN4(input_factor_02[16]), .QN(n14) );
  NOR4X0 U20 ( .IN1(input_factor_02[17]), .IN2(input_factor_02[18]), .IN3(
        input_factor_02[19]), .IN4(input_factor_02[1]), .QN(n13) );
  NOR4X0 U21 ( .IN1(input_factor_02[20]), .IN2(input_factor_02[21]), .IN3(
        input_factor_02[22]), .IN4(input_factor_02[23]), .QN(n12) );
  NAND4X0 U22 ( .IN1(n15), .IN2(n14), .IN3(n13), .IN4(n12), .QN(n21) );
  NOR4X0 U23 ( .IN1(input_factor_02[24]), .IN2(input_factor_02[25]), .IN3(
        input_factor_02[26]), .IN4(input_factor_02[27]), .QN(n19) );
  NOR4X0 U24 ( .IN1(input_factor_02[28]), .IN2(input_factor_02[29]), .IN3(
        input_factor_02[2]), .IN4(input_factor_02[30]), .QN(n18) );
  NOR4X0 U25 ( .IN1(input_factor_02[31]), .IN2(input_factor_02[3]), .IN3(
        input_factor_02[4]), .IN4(input_factor_02[5]), .QN(n17) );
  NOR4X0 U26 ( .IN1(input_factor_02[6]), .IN2(input_factor_02[7]), .IN3(
        input_factor_02[8]), .IN4(input_factor_02[9]), .QN(n16) );
  NAND4X0 U27 ( .IN1(n19), .IN2(n18), .IN3(n17), .IN4(n16), .QN(n20) );
  OA22X1 U28 ( .IN1(n23), .IN2(n22), .IN3(n21), .IN4(n20), .Q(n35) );
  INVX0 U29 ( .INP(n35), .ZN(n24) );
  AO22X1 U30 ( .IN1(n2), .IN2(base_multiply_result[23]), .IN3(n32), .IN4(
        base_multiply_result[24]), .Q(N10) );
  AO22X1 U31 ( .IN1(n2), .IN2(base_multiply_result[24]), .IN3(n32), .IN4(
        base_multiply_result[25]), .Q(N11) );
  AO22X1 U32 ( .IN1(n2), .IN2(base_multiply_result[25]), .IN3(n32), .IN4(
        base_multiply_result[26]), .Q(N12) );
  AO22X1 U33 ( .IN1(n2), .IN2(base_multiply_result[26]), .IN3(n32), .IN4(
        base_multiply_result[27]), .Q(N13) );
  AO22X1 U34 ( .IN1(n2), .IN2(base_multiply_result[27]), .IN3(n32), .IN4(
        base_multiply_result[28]), .Q(N14) );
  AO22X1 U35 ( .IN1(n2), .IN2(base_multiply_result[28]), .IN3(n32), .IN4(
        base_multiply_result[29]), .Q(N15) );
  AO22X1 U36 ( .IN1(n2), .IN2(base_multiply_result[29]), .IN3(n32), .IN4(
        base_multiply_result[30]), .Q(N16) );
  AO22X1 U37 ( .IN1(n2), .IN2(base_multiply_result[30]), .IN3(n32), .IN4(
        base_multiply_result[31]), .Q(N17) );
  AO22X1 U38 ( .IN1(n2), .IN2(base_multiply_result[31]), .IN3(n32), .IN4(
        base_multiply_result[32]), .Q(N18) );
  AO22X1 U39 ( .IN1(n2), .IN2(base_multiply_result[32]), .IN3(n32), .IN4(
        base_multiply_result[33]), .Q(N19) );
  AO22X1 U40 ( .IN1(n2), .IN2(base_multiply_result[33]), .IN3(n32), .IN4(
        base_multiply_result[34]), .Q(N20) );
  AO22X1 U41 ( .IN1(n2), .IN2(base_multiply_result[34]), .IN3(n32), .IN4(
        base_multiply_result[35]), .Q(N21) );
  AO22X1 U42 ( .IN1(n2), .IN2(base_multiply_result[35]), .IN3(n32), .IN4(
        base_multiply_result[36]), .Q(N22) );
  AO22X1 U43 ( .IN1(n2), .IN2(base_multiply_result[36]), .IN3(n32), .IN4(
        base_multiply_result[37]), .Q(N23) );
  AO22X1 U44 ( .IN1(n2), .IN2(base_multiply_result[37]), .IN3(n32), .IN4(
        base_multiply_result[38]), .Q(N24) );
  AO22X1 U45 ( .IN1(n2), .IN2(base_multiply_result[38]), .IN3(n32), .IN4(
        base_multiply_result[39]), .Q(N25) );
  AO22X1 U46 ( .IN1(n2), .IN2(base_multiply_result[39]), .IN3(n32), .IN4(
        base_multiply_result[40]), .Q(N26) );
  AO22X1 U47 ( .IN1(n2), .IN2(base_multiply_result[40]), .IN3(n32), .IN4(
        base_multiply_result[41]), .Q(N27) );
  AO22X1 U48 ( .IN1(n2), .IN2(base_multiply_result[41]), .IN3(n32), .IN4(
        base_multiply_result[42]), .Q(N28) );
  AO22X1 U49 ( .IN1(n2), .IN2(base_multiply_result[42]), .IN3(n32), .IN4(
        base_multiply_result[43]), .Q(N29) );
  AO22X1 U50 ( .IN1(n2), .IN2(base_multiply_result[43]), .IN3(n32), .IN4(
        base_multiply_result[44]), .Q(N30) );
  AO22X1 U51 ( .IN1(n2), .IN2(base_multiply_result[44]), .IN3(n32), .IN4(
        base_multiply_result[45]), .Q(N31) );
  AO22X1 U52 ( .IN1(n2), .IN2(base_multiply_result[45]), .IN3(n32), .IN4(
        base_multiply_result[46]), .Q(N32) );
  MUX21X1 U53 ( .IN1(n2), .IN2(n32), .S(pre_mul_output_exponent[0]), .Q(N48)
         );
  AO21X1 U54 ( .IN1(pre_mul_output_exponent[0]), .IN2(n2), .IN3(n32), .Q(n25)
         );
  NOR3X0 U55 ( .IN1(pre_mul_output_exponent[1]), .IN2(
        pre_mul_output_exponent[0]), .IN3(n1), .QN(n27) );
  AO21X1 U56 ( .IN1(pre_mul_output_exponent[1]), .IN2(n25), .IN3(n27), .Q(N49)
         );
  INVX0 U57 ( .INP(input_factor_01[31]), .ZN(n26) );
  OA221X1 U58 ( .IN1(input_factor_01[31]), .IN2(input_factor_02[31]), .IN3(n26), .IN4(n3), .IN5(n35), .Q(N5) );
  AO221X1 U59 ( .IN1(n2), .IN2(pre_mul_output_exponent[1]), .IN3(n2), .IN4(
        pre_mul_output_exponent[0]), .IN5(n32), .Q(n28) );
  MUX21X1 U60 ( .IN1(n27), .IN2(n28), .S(pre_mul_output_exponent[2]), .Q(N50)
         );
  AND2X1 U61 ( .IN1(n2), .IN2(pre_mul_output_exponent[2]), .Q(n29) );
  OR4X1 U62 ( .IN1(pre_mul_output_exponent[1]), .IN2(
        pre_mul_output_exponent[0]), .IN3(pre_mul_output_exponent[3]), .IN4(
        pre_mul_output_exponent[2]), .Q(n34) );
  NOR2X0 U63 ( .IN1(n1), .IN2(n34), .QN(n31) );
  AO221X1 U64 ( .IN1(pre_mul_output_exponent[3]), .IN2(n29), .IN3(
        pre_mul_output_exponent[3]), .IN4(n28), .IN5(n31), .Q(N51) );
  OA21X1 U65 ( .IN1(base_multiply_result[47]), .IN2(n34), .IN3(n35), .Q(n30)
         );
  MUX21X1 U66 ( .IN1(n31), .IN2(n30), .S(pre_mul_output_exponent[4]), .Q(N52)
         );
  AO221X1 U67 ( .IN1(n2), .IN2(pre_mul_output_exponent[4]), .IN3(n2), .IN4(n34), .IN5(n32), .Q(n33) );
  NOR4X0 U68 ( .IN1(pre_mul_output_exponent[5]), .IN2(
        pre_mul_output_exponent[4]), .IN3(n34), .IN4(n1), .QN(n37) );
  AO21X1 U69 ( .IN1(pre_mul_output_exponent[5]), .IN2(n33), .IN3(n37), .Q(N53)
         );
  OR3X1 U70 ( .IN1(pre_mul_output_exponent[5]), .IN2(
        pre_mul_output_exponent[4]), .IN3(n34), .Q(n36) );
  OA21X1 U71 ( .IN1(base_multiply_result[47]), .IN2(n36), .IN3(n35), .Q(n39)
         );
  INVX0 U72 ( .INP(n37), .ZN(n38) );
  NOR2X0 U73 ( .IN1(pre_mul_output_exponent[6]), .IN2(n38), .QN(n41) );
  AO21X1 U74 ( .IN1(pre_mul_output_exponent[6]), .IN2(n39), .IN3(n41), .Q(N54)
         );
  AO21X1 U75 ( .IN1(n2), .IN2(pre_mul_output_exponent[6]), .IN3(n39), .Q(n40)
         );
  MUX21X1 U76 ( .IN1(n41), .IN2(n40), .S(pre_mul_output_exponent[7]), .Q(N55)
         );
endmodule


module sigmoid_function ( clk, rst_n, sigmoid_input, sigmoid_output );
  input [31:0] sigmoid_input;
  output [31:0] sigmoid_output;
  input clk, rst_n;
  wire   SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13;
  wire   [31:0] factor_a;
  wire   [31:0] factor_b;
  wire   [31:0] factor_c;
  wire   [31:0] factor_d;
  wire   [31:0] next_factor_a;
  wire   [31:0] next_factor_b;
  wire   [31:0] next_factor_c;
  wire   [31:0] next_factor_d;
  wire   [31:0] result_mult_b;
  wire   [31:0] next_result_mult_b;
  wire   [31:0] result_adder_b;
  wire   [31:0] next_result_adder_b;
  wire   [31:0] result_mult_c;
  wire   [31:0] next_result_mult_c;
  wire   [31:0] result_adder_c;
  wire   [31:0] next_result_adder_c;
  wire   [31:0] result_mult_d;
  wire   [31:0] next_result_mult_d;
  wire   [31:0] result_adder_d;

  sigmoid_floating_point_compare floating_point_compare_01 ( .clk(clk), 
        .rst_n(rst_n), .factor_input(sigmoid_input), .factor_a({factor_a[31], 
        SYNOPSYS_UNCONNECTED_1, factor_a[29:14], SYNOPSYS_UNCONNECTED_2, 
        factor_a[12:7], SYNOPSYS_UNCONNECTED_3, factor_a[5:0]}), .factor_b({
        factor_b[31], SYNOPSYS_UNCONNECTED_4, factor_b[29:23], 
        SYNOPSYS_UNCONNECTED_5, factor_b[21:20], SYNOPSYS_UNCONNECTED_6, 
        SYNOPSYS_UNCONNECTED_7, factor_b[17:0]}), .factor_c({factor_c[31], 
        SYNOPSYS_UNCONNECTED_8, factor_c[29:21], SYNOPSYS_UNCONNECTED_9, 
        factor_c[19:13], SYNOPSYS_UNCONNECTED_10, factor_c[11:2], 
        SYNOPSYS_UNCONNECTED_11, factor_c[0]}), .factor_d({factor_d[31], 
        SYNOPSYS_UNCONNECTED_12, factor_d[29:15], SYNOPSYS_UNCONNECTED_13, 
        factor_d[13:0]}) );
  floating_point_multiple_6 multiple_01 ( .clk(clk), .rst_n(rst_n), 
        .input_factor_01({next_factor_a[31], 1'b0, next_factor_a[29:14], 1'b0, 
        next_factor_a[12:7], 1'b0, next_factor_a[5:0]}), .input_factor_02(
        sigmoid_input), .output_multiply(result_mult_b) );
  floating_point_adder_6 adder_01 ( .clk(clk), .rst_n(rst_n), 
        .input_factor_01(next_result_mult_b), .input_factor_02({
        next_factor_b[31], 1'b0, next_factor_b[29:23], 1'b0, 
        next_factor_b[21:20], 1'b0, 1'b0, next_factor_b[17:0]}), 
        .output_adder(result_adder_b) );
  floating_point_multiple_5 multiple_02 ( .clk(clk), .rst_n(rst_n), 
        .input_factor_01(next_result_adder_b), .input_factor_02(sigmoid_input), 
        .output_multiply(result_mult_c) );
  floating_point_adder_5 adder_02 ( .clk(clk), .rst_n(rst_n), 
        .input_factor_01(next_result_mult_c), .input_factor_02({
        next_factor_c[31], 1'b0, next_factor_c[29:21], 1'b0, 
        next_factor_c[19:13], 1'b0, next_factor_c[11:2], 1'b0, 
        next_factor_c[0]}), .output_adder(result_adder_c) );
  floating_point_multiple_4 multiple_03 ( .clk(clk), .rst_n(rst_n), 
        .input_factor_01(next_result_adder_c), .input_factor_02(sigmoid_input), 
        .output_multiply(result_mult_d) );
  floating_point_adder_4 adder_03 ( .clk(clk), .rst_n(rst_n), 
        .input_factor_01(next_result_mult_d), .input_factor_02({
        next_factor_d[31], 1'b0, next_factor_d[29:15], 1'b0, 
        next_factor_d[13:0]}), .output_adder(result_adder_d) );
  DFFARX1 next_factor_a_reg_31_ ( .D(factor_a[31]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_a[31]) );
  DFFARX1 next_factor_a_reg_29_ ( .D(factor_a[29]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_a[29]) );
  DFFARX1 next_factor_a_reg_28_ ( .D(factor_a[28]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_a[28]) );
  DFFARX1 next_factor_a_reg_27_ ( .D(factor_a[27]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_a[27]) );
  DFFARX1 next_factor_a_reg_26_ ( .D(factor_a[26]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_a[26]) );
  DFFARX1 next_factor_a_reg_25_ ( .D(factor_a[25]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_a[25]) );
  DFFARX1 next_factor_a_reg_24_ ( .D(factor_a[24]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_a[24]) );
  DFFARX1 next_factor_a_reg_23_ ( .D(factor_a[23]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_a[23]) );
  DFFARX1 next_factor_a_reg_22_ ( .D(factor_a[22]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_a[22]) );
  DFFARX1 next_factor_a_reg_21_ ( .D(factor_a[21]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_a[21]) );
  DFFARX1 next_factor_a_reg_20_ ( .D(factor_a[20]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_a[20]) );
  DFFARX1 next_factor_a_reg_19_ ( .D(factor_a[19]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_a[19]) );
  DFFARX1 next_factor_a_reg_18_ ( .D(factor_a[18]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_a[18]) );
  DFFARX1 next_factor_a_reg_17_ ( .D(factor_a[17]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_a[17]) );
  DFFARX1 next_factor_a_reg_16_ ( .D(factor_a[16]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_a[16]) );
  DFFARX1 next_factor_a_reg_15_ ( .D(factor_a[15]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_a[15]) );
  DFFARX1 next_factor_a_reg_14_ ( .D(factor_a[14]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_a[14]) );
  DFFARX1 next_factor_a_reg_12_ ( .D(factor_a[12]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_a[12]) );
  DFFARX1 next_factor_a_reg_11_ ( .D(factor_a[11]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_a[11]) );
  DFFARX1 next_factor_a_reg_10_ ( .D(factor_a[10]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_a[10]) );
  DFFARX1 next_factor_a_reg_9_ ( .D(factor_a[9]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_a[9]) );
  DFFARX1 next_factor_a_reg_8_ ( .D(factor_a[8]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_a[8]) );
  DFFARX1 next_factor_a_reg_7_ ( .D(factor_a[7]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_a[7]) );
  DFFARX1 next_factor_a_reg_5_ ( .D(factor_a[5]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_a[5]) );
  DFFARX1 next_factor_a_reg_4_ ( .D(factor_a[4]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_a[4]) );
  DFFARX1 next_factor_a_reg_3_ ( .D(factor_a[3]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_a[3]) );
  DFFARX1 next_factor_a_reg_2_ ( .D(factor_a[2]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_a[2]) );
  DFFARX1 next_factor_a_reg_1_ ( .D(factor_a[1]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_a[1]) );
  DFFARX1 next_factor_a_reg_0_ ( .D(factor_a[0]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_a[0]) );
  DFFARX1 next_factor_b_reg_31_ ( .D(factor_b[31]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_b[31]) );
  DFFARX1 next_factor_b_reg_29_ ( .D(factor_b[29]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_b[29]) );
  DFFARX1 next_factor_b_reg_28_ ( .D(factor_b[28]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_b[28]) );
  DFFARX1 next_factor_b_reg_27_ ( .D(factor_b[27]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_b[27]) );
  DFFARX1 next_factor_b_reg_26_ ( .D(factor_b[26]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_b[26]) );
  DFFARX1 next_factor_b_reg_25_ ( .D(factor_b[25]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_b[25]) );
  DFFARX1 next_factor_b_reg_24_ ( .D(factor_b[24]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_b[24]) );
  DFFARX1 next_factor_b_reg_23_ ( .D(factor_b[23]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_b[23]) );
  DFFARX1 next_factor_b_reg_21_ ( .D(factor_b[21]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_b[21]) );
  DFFARX1 next_factor_b_reg_20_ ( .D(factor_b[20]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_b[20]) );
  DFFARX1 next_factor_b_reg_17_ ( .D(factor_b[17]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_b[17]) );
  DFFARX1 next_factor_b_reg_16_ ( .D(factor_b[16]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_b[16]) );
  DFFARX1 next_factor_b_reg_15_ ( .D(factor_b[15]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_b[15]) );
  DFFARX1 next_factor_b_reg_14_ ( .D(factor_b[14]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_b[14]) );
  DFFARX1 next_factor_b_reg_13_ ( .D(factor_b[13]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_b[13]) );
  DFFARX1 next_factor_b_reg_12_ ( .D(factor_b[12]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_b[12]) );
  DFFARX1 next_factor_b_reg_11_ ( .D(factor_b[11]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_b[11]) );
  DFFARX1 next_factor_b_reg_10_ ( .D(factor_b[10]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_b[10]) );
  DFFARX1 next_factor_b_reg_9_ ( .D(factor_b[9]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_b[9]) );
  DFFARX1 next_factor_b_reg_8_ ( .D(factor_b[8]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_b[8]) );
  DFFARX1 next_factor_b_reg_7_ ( .D(factor_b[7]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_b[7]) );
  DFFARX1 next_factor_b_reg_6_ ( .D(factor_b[6]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_b[6]) );
  DFFARX1 next_factor_b_reg_5_ ( .D(factor_b[5]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_b[5]) );
  DFFARX1 next_factor_b_reg_4_ ( .D(factor_b[4]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_b[4]) );
  DFFARX1 next_factor_b_reg_3_ ( .D(factor_b[3]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_b[3]) );
  DFFARX1 next_factor_b_reg_2_ ( .D(factor_b[2]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_b[2]) );
  DFFARX1 next_factor_b_reg_1_ ( .D(factor_b[1]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_b[1]) );
  DFFARX1 next_factor_b_reg_0_ ( .D(factor_b[0]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_b[0]) );
  DFFARX1 next_factor_c_reg_31_ ( .D(factor_c[31]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_c[31]) );
  DFFARX1 next_factor_c_reg_29_ ( .D(factor_c[29]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_c[29]) );
  DFFARX1 next_factor_c_reg_28_ ( .D(factor_c[28]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_c[28]) );
  DFFARX1 next_factor_c_reg_27_ ( .D(factor_c[27]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_c[27]) );
  DFFARX1 next_factor_c_reg_26_ ( .D(factor_c[26]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_c[26]) );
  DFFARX1 next_factor_c_reg_25_ ( .D(factor_c[25]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_c[25]) );
  DFFARX1 next_factor_c_reg_24_ ( .D(factor_c[24]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_c[24]) );
  DFFARX1 next_factor_c_reg_23_ ( .D(factor_c[23]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_c[23]) );
  DFFARX1 next_factor_c_reg_22_ ( .D(factor_c[22]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_c[22]) );
  DFFARX1 next_factor_c_reg_21_ ( .D(factor_c[21]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_c[21]) );
  DFFARX1 next_factor_c_reg_19_ ( .D(factor_c[19]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_c[19]) );
  DFFARX1 next_factor_c_reg_18_ ( .D(factor_c[18]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_c[18]) );
  DFFARX1 next_factor_c_reg_17_ ( .D(factor_c[17]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_c[17]) );
  DFFARX1 next_factor_c_reg_16_ ( .D(factor_c[16]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_c[16]) );
  DFFARX1 next_factor_c_reg_15_ ( .D(factor_c[15]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_c[15]) );
  DFFARX1 next_factor_c_reg_14_ ( .D(factor_c[14]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_c[14]) );
  DFFARX1 next_factor_c_reg_13_ ( .D(factor_c[13]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_c[13]) );
  DFFARX1 next_factor_c_reg_11_ ( .D(factor_c[11]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_c[11]) );
  DFFARX1 next_factor_c_reg_10_ ( .D(factor_c[10]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_c[10]) );
  DFFARX1 next_factor_c_reg_9_ ( .D(factor_c[9]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_c[9]) );
  DFFARX1 next_factor_c_reg_8_ ( .D(factor_c[8]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_c[8]) );
  DFFARX1 next_factor_c_reg_7_ ( .D(factor_c[7]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_c[7]) );
  DFFARX1 next_factor_c_reg_6_ ( .D(factor_c[6]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_c[6]) );
  DFFARX1 next_factor_c_reg_5_ ( .D(factor_c[5]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_c[5]) );
  DFFARX1 next_factor_c_reg_4_ ( .D(factor_c[4]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_c[4]) );
  DFFARX1 next_factor_c_reg_3_ ( .D(factor_c[3]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_c[3]) );
  DFFARX1 next_factor_c_reg_2_ ( .D(factor_c[2]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_c[2]) );
  DFFARX1 next_factor_c_reg_0_ ( .D(factor_c[0]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_c[0]) );
  DFFARX1 next_factor_d_reg_31_ ( .D(factor_d[31]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_d[31]) );
  DFFARX1 next_factor_d_reg_29_ ( .D(factor_d[29]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_d[29]) );
  DFFARX1 next_factor_d_reg_28_ ( .D(factor_d[28]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_d[28]) );
  DFFARX1 next_factor_d_reg_27_ ( .D(factor_d[27]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_d[27]) );
  DFFARX1 next_factor_d_reg_26_ ( .D(factor_d[26]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_d[26]) );
  DFFARX1 next_factor_d_reg_25_ ( .D(factor_d[25]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_d[25]) );
  DFFARX1 next_factor_d_reg_24_ ( .D(factor_d[24]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_d[24]) );
  DFFARX1 next_factor_d_reg_23_ ( .D(factor_d[23]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_d[23]) );
  DFFARX1 next_factor_d_reg_22_ ( .D(factor_d[22]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_d[22]) );
  DFFARX1 next_factor_d_reg_21_ ( .D(factor_d[21]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_d[21]) );
  DFFARX1 next_factor_d_reg_20_ ( .D(factor_d[20]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_d[20]) );
  DFFARX1 next_factor_d_reg_19_ ( .D(factor_d[19]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_d[19]) );
  DFFARX1 next_factor_d_reg_18_ ( .D(factor_d[18]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_d[18]) );
  DFFARX1 next_factor_d_reg_17_ ( .D(factor_d[17]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_d[17]) );
  DFFARX1 next_factor_d_reg_16_ ( .D(factor_d[16]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_d[16]) );
  DFFARX1 next_factor_d_reg_15_ ( .D(factor_d[15]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_d[15]) );
  DFFARX1 next_factor_d_reg_13_ ( .D(factor_d[13]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_d[13]) );
  DFFARX1 next_factor_d_reg_12_ ( .D(factor_d[12]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_d[12]) );
  DFFARX1 next_factor_d_reg_11_ ( .D(factor_d[11]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_d[11]) );
  DFFARX1 next_factor_d_reg_10_ ( .D(factor_d[10]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_d[10]) );
  DFFARX1 next_factor_d_reg_9_ ( .D(factor_d[9]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_d[9]) );
  DFFARX1 next_factor_d_reg_8_ ( .D(factor_d[8]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_d[8]) );
  DFFARX1 next_factor_d_reg_7_ ( .D(factor_d[7]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_d[7]) );
  DFFARX1 next_factor_d_reg_6_ ( .D(factor_d[6]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_d[6]) );
  DFFARX1 next_factor_d_reg_5_ ( .D(factor_d[5]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_d[5]) );
  DFFARX1 next_factor_d_reg_4_ ( .D(factor_d[4]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_d[4]) );
  DFFARX1 next_factor_d_reg_3_ ( .D(factor_d[3]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_d[3]) );
  DFFARX1 next_factor_d_reg_2_ ( .D(factor_d[2]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_d[2]) );
  DFFARX1 next_factor_d_reg_1_ ( .D(factor_d[1]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_d[1]) );
  DFFARX1 next_factor_d_reg_0_ ( .D(factor_d[0]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_d[0]) );
  DFFARX1 next_result_mult_b_reg_31_ ( .D(result_mult_b[31]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_b[31]) );
  DFFARX1 next_result_mult_b_reg_30_ ( .D(result_mult_b[30]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_b[30]) );
  DFFARX1 next_result_mult_b_reg_29_ ( .D(result_mult_b[29]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_b[29]) );
  DFFARX1 next_result_mult_b_reg_28_ ( .D(result_mult_b[28]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_b[28]) );
  DFFARX1 next_result_mult_b_reg_27_ ( .D(result_mult_b[27]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_b[27]) );
  DFFARX1 next_result_mult_b_reg_26_ ( .D(result_mult_b[26]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_b[26]) );
  DFFARX1 next_result_mult_b_reg_25_ ( .D(result_mult_b[25]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_b[25]) );
  DFFARX1 next_result_mult_b_reg_24_ ( .D(result_mult_b[24]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_b[24]) );
  DFFARX1 next_result_mult_b_reg_23_ ( .D(result_mult_b[23]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_b[23]) );
  DFFARX1 next_result_mult_b_reg_22_ ( .D(result_mult_b[22]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_b[22]) );
  DFFARX1 next_result_mult_b_reg_21_ ( .D(result_mult_b[21]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_b[21]) );
  DFFARX1 next_result_mult_b_reg_20_ ( .D(result_mult_b[20]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_b[20]) );
  DFFARX1 next_result_mult_b_reg_19_ ( .D(result_mult_b[19]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_b[19]) );
  DFFARX1 next_result_mult_b_reg_18_ ( .D(result_mult_b[18]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_b[18]) );
  DFFARX1 next_result_mult_b_reg_17_ ( .D(result_mult_b[17]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_b[17]) );
  DFFARX1 next_result_mult_b_reg_16_ ( .D(result_mult_b[16]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_b[16]) );
  DFFARX1 next_result_mult_b_reg_15_ ( .D(result_mult_b[15]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_b[15]) );
  DFFARX1 next_result_mult_b_reg_14_ ( .D(result_mult_b[14]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_b[14]) );
  DFFARX1 next_result_mult_b_reg_13_ ( .D(result_mult_b[13]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_b[13]) );
  DFFARX1 next_result_mult_b_reg_12_ ( .D(result_mult_b[12]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_b[12]) );
  DFFARX1 next_result_mult_b_reg_11_ ( .D(result_mult_b[11]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_b[11]) );
  DFFARX1 next_result_mult_b_reg_10_ ( .D(result_mult_b[10]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_b[10]) );
  DFFARX1 next_result_mult_b_reg_9_ ( .D(result_mult_b[9]), .CLK(clk), .RSTB(
        rst_n), .Q(next_result_mult_b[9]) );
  DFFARX1 next_result_mult_b_reg_8_ ( .D(result_mult_b[8]), .CLK(clk), .RSTB(
        rst_n), .Q(next_result_mult_b[8]) );
  DFFARX1 next_result_mult_b_reg_7_ ( .D(result_mult_b[7]), .CLK(clk), .RSTB(
        rst_n), .Q(next_result_mult_b[7]) );
  DFFARX1 next_result_mult_b_reg_6_ ( .D(result_mult_b[6]), .CLK(clk), .RSTB(
        rst_n), .Q(next_result_mult_b[6]) );
  DFFARX1 next_result_mult_b_reg_5_ ( .D(result_mult_b[5]), .CLK(clk), .RSTB(
        rst_n), .Q(next_result_mult_b[5]) );
  DFFARX1 next_result_mult_b_reg_4_ ( .D(result_mult_b[4]), .CLK(clk), .RSTB(
        rst_n), .Q(next_result_mult_b[4]) );
  DFFARX1 next_result_mult_b_reg_3_ ( .D(result_mult_b[3]), .CLK(clk), .RSTB(
        rst_n), .Q(next_result_mult_b[3]) );
  DFFARX1 next_result_mult_b_reg_2_ ( .D(result_mult_b[2]), .CLK(clk), .RSTB(
        rst_n), .Q(next_result_mult_b[2]) );
  DFFARX1 next_result_mult_b_reg_1_ ( .D(result_mult_b[1]), .CLK(clk), .RSTB(
        rst_n), .Q(next_result_mult_b[1]) );
  DFFARX1 next_result_mult_b_reg_0_ ( .D(result_mult_b[0]), .CLK(clk), .RSTB(
        rst_n), .Q(next_result_mult_b[0]) );
  DFFARX1 next_result_adder_b_reg_31_ ( .D(result_adder_b[31]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[31]) );
  DFFARX1 next_result_adder_b_reg_30_ ( .D(result_adder_b[30]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[30]) );
  DFFARX1 next_result_adder_b_reg_29_ ( .D(result_adder_b[29]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[29]) );
  DFFARX1 next_result_adder_b_reg_28_ ( .D(result_adder_b[28]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[28]) );
  DFFARX1 next_result_adder_b_reg_27_ ( .D(result_adder_b[27]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[27]) );
  DFFARX1 next_result_adder_b_reg_26_ ( .D(result_adder_b[26]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[26]) );
  DFFARX1 next_result_adder_b_reg_25_ ( .D(result_adder_b[25]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[25]) );
  DFFARX1 next_result_adder_b_reg_24_ ( .D(result_adder_b[24]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[24]) );
  DFFARX1 next_result_adder_b_reg_23_ ( .D(result_adder_b[23]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[23]) );
  DFFARX1 next_result_adder_b_reg_22_ ( .D(result_adder_b[22]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[22]) );
  DFFARX1 next_result_adder_b_reg_21_ ( .D(result_adder_b[21]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[21]) );
  DFFARX1 next_result_adder_b_reg_20_ ( .D(result_adder_b[20]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[20]) );
  DFFARX1 next_result_adder_b_reg_19_ ( .D(result_adder_b[19]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[19]) );
  DFFARX1 next_result_adder_b_reg_18_ ( .D(result_adder_b[18]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[18]) );
  DFFARX1 next_result_adder_b_reg_17_ ( .D(result_adder_b[17]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[17]) );
  DFFARX1 next_result_adder_b_reg_16_ ( .D(result_adder_b[16]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[16]) );
  DFFARX1 next_result_adder_b_reg_15_ ( .D(result_adder_b[15]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[15]) );
  DFFARX1 next_result_adder_b_reg_14_ ( .D(result_adder_b[14]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[14]) );
  DFFARX1 next_result_adder_b_reg_13_ ( .D(result_adder_b[13]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[13]) );
  DFFARX1 next_result_adder_b_reg_12_ ( .D(result_adder_b[12]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[12]) );
  DFFARX1 next_result_adder_b_reg_11_ ( .D(result_adder_b[11]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[11]) );
  DFFARX1 next_result_adder_b_reg_10_ ( .D(result_adder_b[10]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[10]) );
  DFFARX1 next_result_adder_b_reg_9_ ( .D(result_adder_b[9]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[9]) );
  DFFARX1 next_result_adder_b_reg_8_ ( .D(result_adder_b[8]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[8]) );
  DFFARX1 next_result_adder_b_reg_7_ ( .D(result_adder_b[7]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[7]) );
  DFFARX1 next_result_adder_b_reg_6_ ( .D(result_adder_b[6]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[6]) );
  DFFARX1 next_result_adder_b_reg_5_ ( .D(result_adder_b[5]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[5]) );
  DFFARX1 next_result_adder_b_reg_4_ ( .D(result_adder_b[4]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[4]) );
  DFFARX1 next_result_adder_b_reg_3_ ( .D(result_adder_b[3]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[3]) );
  DFFARX1 next_result_adder_b_reg_2_ ( .D(result_adder_b[2]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[2]) );
  DFFARX1 next_result_adder_b_reg_1_ ( .D(result_adder_b[1]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[1]) );
  DFFARX1 next_result_adder_b_reg_0_ ( .D(result_adder_b[0]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[0]) );
  DFFARX1 next_result_mult_c_reg_31_ ( .D(result_mult_c[31]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_c[31]) );
  DFFARX1 next_result_mult_c_reg_30_ ( .D(result_mult_c[30]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_c[30]) );
  DFFARX1 next_result_mult_c_reg_29_ ( .D(result_mult_c[29]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_c[29]) );
  DFFARX1 next_result_mult_c_reg_28_ ( .D(result_mult_c[28]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_c[28]) );
  DFFARX1 next_result_mult_c_reg_27_ ( .D(result_mult_c[27]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_c[27]) );
  DFFARX1 next_result_mult_c_reg_26_ ( .D(result_mult_c[26]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_c[26]) );
  DFFARX1 next_result_mult_c_reg_25_ ( .D(result_mult_c[25]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_c[25]) );
  DFFARX1 next_result_mult_c_reg_24_ ( .D(result_mult_c[24]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_c[24]) );
  DFFARX1 next_result_mult_c_reg_23_ ( .D(result_mult_c[23]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_c[23]) );
  DFFARX1 next_result_mult_c_reg_22_ ( .D(result_mult_c[22]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_c[22]) );
  DFFARX1 next_result_mult_c_reg_21_ ( .D(result_mult_c[21]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_c[21]) );
  DFFARX1 next_result_mult_c_reg_20_ ( .D(result_mult_c[20]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_c[20]) );
  DFFARX1 next_result_mult_c_reg_19_ ( .D(result_mult_c[19]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_c[19]) );
  DFFARX1 next_result_mult_c_reg_18_ ( .D(result_mult_c[18]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_c[18]) );
  DFFARX1 next_result_mult_c_reg_17_ ( .D(result_mult_c[17]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_c[17]) );
  DFFARX1 next_result_mult_c_reg_16_ ( .D(result_mult_c[16]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_c[16]) );
  DFFARX1 next_result_mult_c_reg_15_ ( .D(result_mult_c[15]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_c[15]) );
  DFFARX1 next_result_mult_c_reg_14_ ( .D(result_mult_c[14]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_c[14]) );
  DFFARX1 next_result_mult_c_reg_13_ ( .D(result_mult_c[13]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_c[13]) );
  DFFARX1 next_result_mult_c_reg_12_ ( .D(result_mult_c[12]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_c[12]) );
  DFFARX1 next_result_mult_c_reg_11_ ( .D(result_mult_c[11]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_c[11]) );
  DFFARX1 next_result_mult_c_reg_10_ ( .D(result_mult_c[10]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_c[10]) );
  DFFARX1 next_result_mult_c_reg_9_ ( .D(result_mult_c[9]), .CLK(clk), .RSTB(
        rst_n), .Q(next_result_mult_c[9]) );
  DFFARX1 next_result_mult_c_reg_8_ ( .D(result_mult_c[8]), .CLK(clk), .RSTB(
        rst_n), .Q(next_result_mult_c[8]) );
  DFFARX1 next_result_mult_c_reg_7_ ( .D(result_mult_c[7]), .CLK(clk), .RSTB(
        rst_n), .Q(next_result_mult_c[7]) );
  DFFARX1 next_result_mult_c_reg_6_ ( .D(result_mult_c[6]), .CLK(clk), .RSTB(
        rst_n), .Q(next_result_mult_c[6]) );
  DFFARX1 next_result_mult_c_reg_5_ ( .D(result_mult_c[5]), .CLK(clk), .RSTB(
        rst_n), .Q(next_result_mult_c[5]) );
  DFFARX1 next_result_mult_c_reg_4_ ( .D(result_mult_c[4]), .CLK(clk), .RSTB(
        rst_n), .Q(next_result_mult_c[4]) );
  DFFARX1 next_result_mult_c_reg_3_ ( .D(result_mult_c[3]), .CLK(clk), .RSTB(
        rst_n), .Q(next_result_mult_c[3]) );
  DFFARX1 next_result_mult_c_reg_2_ ( .D(result_mult_c[2]), .CLK(clk), .RSTB(
        rst_n), .Q(next_result_mult_c[2]) );
  DFFARX1 next_result_mult_c_reg_1_ ( .D(result_mult_c[1]), .CLK(clk), .RSTB(
        rst_n), .Q(next_result_mult_c[1]) );
  DFFARX1 next_result_mult_c_reg_0_ ( .D(result_mult_c[0]), .CLK(clk), .RSTB(
        rst_n), .Q(next_result_mult_c[0]) );
  DFFARX1 next_result_adder_c_reg_31_ ( .D(result_adder_c[31]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[31]) );
  DFFARX1 next_result_adder_c_reg_30_ ( .D(result_adder_c[30]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[30]) );
  DFFARX1 next_result_adder_c_reg_29_ ( .D(result_adder_c[29]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[29]) );
  DFFARX1 next_result_adder_c_reg_28_ ( .D(result_adder_c[28]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[28]) );
  DFFARX1 next_result_adder_c_reg_27_ ( .D(result_adder_c[27]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[27]) );
  DFFARX1 next_result_adder_c_reg_26_ ( .D(result_adder_c[26]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[26]) );
  DFFARX1 next_result_adder_c_reg_25_ ( .D(result_adder_c[25]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[25]) );
  DFFARX1 next_result_adder_c_reg_24_ ( .D(result_adder_c[24]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[24]) );
  DFFARX1 next_result_adder_c_reg_23_ ( .D(result_adder_c[23]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[23]) );
  DFFARX1 next_result_adder_c_reg_22_ ( .D(result_adder_c[22]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[22]) );
  DFFARX1 next_result_adder_c_reg_21_ ( .D(result_adder_c[21]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[21]) );
  DFFARX1 next_result_adder_c_reg_20_ ( .D(result_adder_c[20]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[20]) );
  DFFARX1 next_result_adder_c_reg_19_ ( .D(result_adder_c[19]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[19]) );
  DFFARX1 next_result_adder_c_reg_18_ ( .D(result_adder_c[18]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[18]) );
  DFFARX1 next_result_adder_c_reg_17_ ( .D(result_adder_c[17]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[17]) );
  DFFARX1 next_result_adder_c_reg_16_ ( .D(result_adder_c[16]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[16]) );
  DFFARX1 next_result_adder_c_reg_15_ ( .D(result_adder_c[15]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[15]) );
  DFFARX1 next_result_adder_c_reg_14_ ( .D(result_adder_c[14]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[14]) );
  DFFARX1 next_result_adder_c_reg_13_ ( .D(result_adder_c[13]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[13]) );
  DFFARX1 next_result_adder_c_reg_12_ ( .D(result_adder_c[12]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[12]) );
  DFFARX1 next_result_adder_c_reg_11_ ( .D(result_adder_c[11]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[11]) );
  DFFARX1 next_result_adder_c_reg_10_ ( .D(result_adder_c[10]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[10]) );
  DFFARX1 next_result_adder_c_reg_9_ ( .D(result_adder_c[9]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[9]) );
  DFFARX1 next_result_adder_c_reg_8_ ( .D(result_adder_c[8]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[8]) );
  DFFARX1 next_result_adder_c_reg_7_ ( .D(result_adder_c[7]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[7]) );
  DFFARX1 next_result_adder_c_reg_6_ ( .D(result_adder_c[6]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[6]) );
  DFFARX1 next_result_adder_c_reg_5_ ( .D(result_adder_c[5]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[5]) );
  DFFARX1 next_result_adder_c_reg_4_ ( .D(result_adder_c[4]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[4]) );
  DFFARX1 next_result_adder_c_reg_3_ ( .D(result_adder_c[3]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[3]) );
  DFFARX1 next_result_adder_c_reg_2_ ( .D(result_adder_c[2]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[2]) );
  DFFARX1 next_result_adder_c_reg_1_ ( .D(result_adder_c[1]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[1]) );
  DFFARX1 next_result_adder_c_reg_0_ ( .D(result_adder_c[0]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[0]) );
  DFFARX1 next_result_mult_d_reg_31_ ( .D(result_mult_d[31]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_d[31]) );
  DFFARX1 next_result_mult_d_reg_30_ ( .D(result_mult_d[30]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_d[30]) );
  DFFARX1 next_result_mult_d_reg_29_ ( .D(result_mult_d[29]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_d[29]) );
  DFFARX1 next_result_mult_d_reg_28_ ( .D(result_mult_d[28]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_d[28]) );
  DFFARX1 next_result_mult_d_reg_27_ ( .D(result_mult_d[27]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_d[27]) );
  DFFARX1 next_result_mult_d_reg_26_ ( .D(result_mult_d[26]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_d[26]) );
  DFFARX1 next_result_mult_d_reg_25_ ( .D(result_mult_d[25]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_d[25]) );
  DFFARX1 next_result_mult_d_reg_24_ ( .D(result_mult_d[24]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_d[24]) );
  DFFARX1 next_result_mult_d_reg_23_ ( .D(result_mult_d[23]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_d[23]) );
  DFFARX1 next_result_mult_d_reg_22_ ( .D(result_mult_d[22]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_d[22]) );
  DFFARX1 next_result_mult_d_reg_21_ ( .D(result_mult_d[21]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_d[21]) );
  DFFARX1 next_result_mult_d_reg_20_ ( .D(result_mult_d[20]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_d[20]) );
  DFFARX1 next_result_mult_d_reg_19_ ( .D(result_mult_d[19]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_d[19]) );
  DFFARX1 next_result_mult_d_reg_18_ ( .D(result_mult_d[18]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_d[18]) );
  DFFARX1 next_result_mult_d_reg_17_ ( .D(result_mult_d[17]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_d[17]) );
  DFFARX1 next_result_mult_d_reg_16_ ( .D(result_mult_d[16]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_d[16]) );
  DFFARX1 next_result_mult_d_reg_15_ ( .D(result_mult_d[15]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_d[15]) );
  DFFARX1 next_result_mult_d_reg_14_ ( .D(result_mult_d[14]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_d[14]) );
  DFFARX1 next_result_mult_d_reg_13_ ( .D(result_mult_d[13]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_d[13]) );
  DFFARX1 next_result_mult_d_reg_12_ ( .D(result_mult_d[12]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_d[12]) );
  DFFARX1 next_result_mult_d_reg_11_ ( .D(result_mult_d[11]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_d[11]) );
  DFFARX1 next_result_mult_d_reg_10_ ( .D(result_mult_d[10]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_d[10]) );
  DFFARX1 next_result_mult_d_reg_9_ ( .D(result_mult_d[9]), .CLK(clk), .RSTB(
        rst_n), .Q(next_result_mult_d[9]) );
  DFFARX1 next_result_mult_d_reg_8_ ( .D(result_mult_d[8]), .CLK(clk), .RSTB(
        rst_n), .Q(next_result_mult_d[8]) );
  DFFARX1 next_result_mult_d_reg_7_ ( .D(result_mult_d[7]), .CLK(clk), .RSTB(
        rst_n), .Q(next_result_mult_d[7]) );
  DFFARX1 next_result_mult_d_reg_6_ ( .D(result_mult_d[6]), .CLK(clk), .RSTB(
        rst_n), .Q(next_result_mult_d[6]) );
  DFFARX1 next_result_mult_d_reg_5_ ( .D(result_mult_d[5]), .CLK(clk), .RSTB(
        rst_n), .Q(next_result_mult_d[5]) );
  DFFARX1 next_result_mult_d_reg_4_ ( .D(result_mult_d[4]), .CLK(clk), .RSTB(
        rst_n), .Q(next_result_mult_d[4]) );
  DFFARX1 next_result_mult_d_reg_3_ ( .D(result_mult_d[3]), .CLK(clk), .RSTB(
        rst_n), .Q(next_result_mult_d[3]) );
  DFFARX1 next_result_mult_d_reg_2_ ( .D(result_mult_d[2]), .CLK(clk), .RSTB(
        rst_n), .Q(next_result_mult_d[2]) );
  DFFARX1 next_result_mult_d_reg_1_ ( .D(result_mult_d[1]), .CLK(clk), .RSTB(
        rst_n), .Q(next_result_mult_d[1]) );
  DFFARX1 next_result_mult_d_reg_0_ ( .D(result_mult_d[0]), .CLK(clk), .RSTB(
        rst_n), .Q(next_result_mult_d[0]) );
  DFFARX1 sigmoid_output_reg_31_ ( .D(result_adder_d[31]), .CLK(clk), .RSTB(
        rst_n), .Q(sigmoid_output[31]) );
  DFFARX1 sigmoid_output_reg_30_ ( .D(result_adder_d[30]), .CLK(clk), .RSTB(
        rst_n), .Q(sigmoid_output[30]) );
  DFFARX1 sigmoid_output_reg_29_ ( .D(result_adder_d[29]), .CLK(clk), .RSTB(
        rst_n), .Q(sigmoid_output[29]) );
  DFFARX1 sigmoid_output_reg_28_ ( .D(result_adder_d[28]), .CLK(clk), .RSTB(
        rst_n), .Q(sigmoid_output[28]) );
  DFFARX1 sigmoid_output_reg_27_ ( .D(result_adder_d[27]), .CLK(clk), .RSTB(
        rst_n), .Q(sigmoid_output[27]) );
  DFFARX1 sigmoid_output_reg_26_ ( .D(result_adder_d[26]), .CLK(clk), .RSTB(
        rst_n), .Q(sigmoid_output[26]) );
  DFFARX1 sigmoid_output_reg_25_ ( .D(result_adder_d[25]), .CLK(clk), .RSTB(
        rst_n), .Q(sigmoid_output[25]) );
  DFFARX1 sigmoid_output_reg_24_ ( .D(result_adder_d[24]), .CLK(clk), .RSTB(
        rst_n), .Q(sigmoid_output[24]) );
  DFFARX1 sigmoid_output_reg_23_ ( .D(result_adder_d[23]), .CLK(clk), .RSTB(
        rst_n), .Q(sigmoid_output[23]) );
  DFFARX1 sigmoid_output_reg_22_ ( .D(result_adder_d[22]), .CLK(clk), .RSTB(
        rst_n), .Q(sigmoid_output[22]) );
  DFFARX1 sigmoid_output_reg_21_ ( .D(result_adder_d[21]), .CLK(clk), .RSTB(
        rst_n), .Q(sigmoid_output[21]) );
  DFFARX1 sigmoid_output_reg_20_ ( .D(result_adder_d[20]), .CLK(clk), .RSTB(
        rst_n), .Q(sigmoid_output[20]) );
  DFFARX1 sigmoid_output_reg_19_ ( .D(result_adder_d[19]), .CLK(clk), .RSTB(
        rst_n), .Q(sigmoid_output[19]) );
  DFFARX1 sigmoid_output_reg_18_ ( .D(result_adder_d[18]), .CLK(clk), .RSTB(
        rst_n), .Q(sigmoid_output[18]) );
  DFFARX1 sigmoid_output_reg_17_ ( .D(result_adder_d[17]), .CLK(clk), .RSTB(
        rst_n), .Q(sigmoid_output[17]) );
  DFFARX1 sigmoid_output_reg_16_ ( .D(result_adder_d[16]), .CLK(clk), .RSTB(
        rst_n), .Q(sigmoid_output[16]) );
  DFFARX1 sigmoid_output_reg_15_ ( .D(result_adder_d[15]), .CLK(clk), .RSTB(
        rst_n), .Q(sigmoid_output[15]) );
  DFFARX1 sigmoid_output_reg_14_ ( .D(result_adder_d[14]), .CLK(clk), .RSTB(
        rst_n), .Q(sigmoid_output[14]) );
  DFFARX1 sigmoid_output_reg_13_ ( .D(result_adder_d[13]), .CLK(clk), .RSTB(
        rst_n), .Q(sigmoid_output[13]) );
  DFFARX1 sigmoid_output_reg_12_ ( .D(result_adder_d[12]), .CLK(clk), .RSTB(
        rst_n), .Q(sigmoid_output[12]) );
  DFFARX1 sigmoid_output_reg_11_ ( .D(result_adder_d[11]), .CLK(clk), .RSTB(
        rst_n), .Q(sigmoid_output[11]) );
  DFFARX1 sigmoid_output_reg_10_ ( .D(result_adder_d[10]), .CLK(clk), .RSTB(
        rst_n), .Q(sigmoid_output[10]) );
  DFFARX1 sigmoid_output_reg_9_ ( .D(result_adder_d[9]), .CLK(clk), .RSTB(
        rst_n), .Q(sigmoid_output[9]) );
  DFFARX1 sigmoid_output_reg_8_ ( .D(result_adder_d[8]), .CLK(clk), .RSTB(
        rst_n), .Q(sigmoid_output[8]) );
  DFFARX1 sigmoid_output_reg_7_ ( .D(result_adder_d[7]), .CLK(clk), .RSTB(
        rst_n), .Q(sigmoid_output[7]) );
  DFFARX1 sigmoid_output_reg_6_ ( .D(result_adder_d[6]), .CLK(clk), .RSTB(
        rst_n), .Q(sigmoid_output[6]) );
  DFFARX1 sigmoid_output_reg_5_ ( .D(result_adder_d[5]), .CLK(clk), .RSTB(
        rst_n), .Q(sigmoid_output[5]) );
  DFFARX1 sigmoid_output_reg_4_ ( .D(result_adder_d[4]), .CLK(clk), .RSTB(
        rst_n), .Q(sigmoid_output[4]) );
  DFFARX1 sigmoid_output_reg_3_ ( .D(result_adder_d[3]), .CLK(clk), .RSTB(
        rst_n), .Q(sigmoid_output[3]) );
  DFFARX1 sigmoid_output_reg_2_ ( .D(result_adder_d[2]), .CLK(clk), .RSTB(
        rst_n), .Q(sigmoid_output[2]) );
  DFFARX1 sigmoid_output_reg_1_ ( .D(result_adder_d[1]), .CLK(clk), .RSTB(
        rst_n), .Q(sigmoid_output[1]) );
  DFFARX1 sigmoid_output_reg_0_ ( .D(result_adder_d[0]), .CLK(clk), .RSTB(
        rst_n), .Q(sigmoid_output[0]) );
endmodule


module tansigmoid_floating_point_compare ( clk, rst_n, factor_input, factor_a, 
        factor_b, factor_c, factor_d );
  input [31:0] factor_input;
  output [31:0] factor_a;
  output [31:0] factor_b;
  output [31:0] factor_c;
  output [31:0] factor_d;
  input clk, rst_n;
  wire   N52, N53, N54, N55, N124, N127, N128, N129, N130, N131, N132, N134,
         N135, N136, N137, N139, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n77, n115, n116, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n76, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155;
  wire   [2:0] case_num;

  DFFARX1 case_num_reg_3_ ( .D(N55), .CLK(clk), .RSTB(rst_n), .Q(n4), .QN(n77)
         );
  DFFARX1 case_num_reg_2_ ( .D(N54), .CLK(clk), .RSTB(rst_n), .Q(case_num[2]), 
        .QN(n1) );
  DFFARX1 case_num_reg_1_ ( .D(N53), .CLK(clk), .RSTB(rst_n), .Q(case_num[1]), 
        .QN(n2) );
  DFFARX1 case_num_reg_0_ ( .D(N52), .CLK(clk), .RSTB(rst_n), .Q(case_num[0]), 
        .QN(n3) );
  DFFARX1 factor_a_reg_31_ ( .D(N136), .CLK(clk), .RSTB(rst_n), .Q(
        factor_a[31]) );
  DFFARX1 factor_a_reg_29_ ( .D(N137), .CLK(clk), .RSTB(rst_n), .Q(
        factor_a[29]) );
  DFFARX1 factor_a_reg_28_ ( .D(N137), .CLK(clk), .RSTB(rst_n), .Q(
        factor_a[28]) );
  DFFARX1 factor_a_reg_27_ ( .D(N137), .CLK(clk), .RSTB(rst_n), .Q(
        factor_a[27]) );
  DFFARX1 factor_a_reg_26_ ( .D(N128), .CLK(clk), .RSTB(rst_n), .Q(
        factor_a[26]) );
  DFFARX1 factor_a_reg_25_ ( .D(N136), .CLK(clk), .RSTB(rst_n), .Q(
        factor_a[25]) );
  DFFARX1 factor_a_reg_24_ ( .D(N134), .CLK(clk), .RSTB(rst_n), .Q(
        factor_a[24]) );
  DFFARX1 factor_a_reg_23_ ( .D(N127), .CLK(clk), .RSTB(rst_n), .Q(
        factor_a[23]) );
  DFFARX1 factor_a_reg_22_ ( .D(N136), .CLK(clk), .RSTB(rst_n), .Q(
        factor_a[22]) );
  DFFARX1 factor_a_reg_21_ ( .D(N135), .CLK(clk), .RSTB(rst_n), .Q(
        factor_a[21]) );
  DFFARX1 factor_a_reg_20_ ( .D(N134), .CLK(clk), .RSTB(rst_n), .Q(
        factor_a[20]) );
  DFFASX1 factor_a_reg_19_ ( .D(n74), .CLK(clk), .SETB(rst_n), .QN(
        factor_a[19]) );
  DFFARX1 factor_a_reg_18_ ( .D(N132), .CLK(clk), .RSTB(rst_n), .Q(
        factor_a[18]) );
  DFFARX1 factor_a_reg_17_ ( .D(N129), .CLK(clk), .RSTB(rst_n), .Q(
        factor_a[17]) );
  DFFARX1 factor_a_reg_16_ ( .D(N130), .CLK(clk), .RSTB(rst_n), .Q(
        factor_a[16]) );
  DFFARX1 factor_a_reg_15_ ( .D(N130), .CLK(clk), .RSTB(rst_n), .Q(
        factor_a[15]) );
  DFFARX1 factor_a_reg_14_ ( .D(N131), .CLK(clk), .RSTB(rst_n), .Q(
        factor_a[14]) );
  DFFASX1 factor_a_reg_12_ ( .D(n75), .CLK(clk), .SETB(rst_n), .QN(
        factor_a[12]) );
  DFFARX1 factor_a_reg_11_ ( .D(N127), .CLK(clk), .RSTB(rst_n), .Q(
        factor_a[11]) );
  DFFARX1 factor_a_reg_10_ ( .D(N130), .CLK(clk), .RSTB(rst_n), .Q(
        factor_a[10]) );
  DFFARX1 factor_a_reg_9_ ( .D(N129), .CLK(clk), .RSTB(rst_n), .Q(factor_a[9])
         );
  DFFARX1 factor_a_reg_8_ ( .D(N128), .CLK(clk), .RSTB(rst_n), .Q(factor_a[8])
         );
  DFFARX1 factor_a_reg_7_ ( .D(N127), .CLK(clk), .RSTB(rst_n), .Q(factor_a[7])
         );
  DFFARX1 factor_a_reg_5_ ( .D(N127), .CLK(clk), .RSTB(rst_n), .Q(factor_a[5])
         );
  DFFASX1 factor_a_reg_4_ ( .D(n75), .CLK(clk), .SETB(rst_n), .QN(factor_a[4])
         );
  DFFASX1 factor_a_reg_3_ ( .D(n116), .CLK(clk), .SETB(rst_n), .QN(factor_a[3]) );
  DFFARX1 factor_a_reg_2_ ( .D(N137), .CLK(clk), .RSTB(rst_n), .Q(factor_a[2])
         );
  DFFARX1 factor_a_reg_1_ ( .D(N124), .CLK(clk), .RSTB(rst_n), .Q(factor_a[1])
         );
  DFFARX1 factor_a_reg_0_ ( .D(N124), .CLK(clk), .RSTB(rst_n), .Q(factor_a[0])
         );
  DFFARX1 factor_b_reg_31_ ( .D(N139), .CLK(clk), .RSTB(rst_n), .Q(
        factor_b[31]) );
  DFFARX1 factor_b_reg_29_ ( .D(N137), .CLK(clk), .RSTB(rst_n), .Q(
        factor_b[29]) );
  DFFARX1 factor_b_reg_28_ ( .D(N137), .CLK(clk), .RSTB(rst_n), .Q(
        factor_b[28]) );
  DFFARX1 factor_b_reg_27_ ( .D(N137), .CLK(clk), .RSTB(rst_n), .Q(
        factor_b[27]) );
  DFFARX1 factor_b_reg_26_ ( .D(N137), .CLK(clk), .RSTB(rst_n), .Q(
        factor_b[26]) );
  DFFARX1 factor_b_reg_25_ ( .D(N124), .CLK(clk), .RSTB(rst_n), .Q(
        factor_b[25]) );
  DFFARX1 factor_b_reg_24_ ( .D(N132), .CLK(clk), .RSTB(rst_n), .Q(
        factor_b[24]) );
  DFFASX1 factor_b_reg_23_ ( .D(n116), .CLK(clk), .SETB(rst_n), .QN(
        factor_b[23]) );
  DFFARX1 factor_b_reg_21_ ( .D(N131), .CLK(clk), .RSTB(rst_n), .Q(
        factor_b[21]) );
  DFFASX1 factor_b_reg_20_ ( .D(n75), .CLK(clk), .SETB(rst_n), .QN(
        factor_b[20]) );
  DFFARX1 factor_b_reg_17_ ( .D(N137), .CLK(clk), .RSTB(rst_n), .Q(
        factor_b[17]) );
  DFFARX1 factor_b_reg_16_ ( .D(N129), .CLK(clk), .RSTB(rst_n), .Q(
        factor_b[16]) );
  DFFARX1 factor_b_reg_15_ ( .D(N131), .CLK(clk), .RSTB(rst_n), .Q(
        factor_b[15]) );
  DFFASX1 factor_b_reg_14_ ( .D(n115), .CLK(clk), .SETB(rst_n), .QN(
        factor_b[14]) );
  DFFARX1 factor_b_reg_13_ ( .D(N131), .CLK(clk), .RSTB(rst_n), .Q(
        factor_b[13]) );
  DFFASX1 factor_b_reg_12_ ( .D(n75), .CLK(clk), .SETB(rst_n), .QN(
        factor_b[12]) );
  DFFARX1 factor_b_reg_11_ ( .D(N127), .CLK(clk), .RSTB(rst_n), .Q(
        factor_b[11]) );
  DFFARX1 factor_b_reg_10_ ( .D(N135), .CLK(clk), .RSTB(rst_n), .Q(
        factor_b[10]) );
  DFFARX1 factor_b_reg_9_ ( .D(N136), .CLK(clk), .RSTB(rst_n), .Q(factor_b[9])
         );
  DFFASX1 factor_b_reg_8_ ( .D(n116), .CLK(clk), .SETB(rst_n), .QN(factor_b[8]) );
  DFFASX1 factor_b_reg_7_ ( .D(n116), .CLK(clk), .SETB(rst_n), .QN(factor_b[7]) );
  DFFARX1 factor_b_reg_6_ ( .D(N124), .CLK(clk), .RSTB(rst_n), .Q(factor_b[6])
         );
  DFFARX1 factor_b_reg_5_ ( .D(N129), .CLK(clk), .RSTB(rst_n), .Q(factor_b[5])
         );
  DFFASX1 factor_b_reg_4_ ( .D(n116), .CLK(clk), .SETB(rst_n), .QN(factor_b[4]) );
  DFFARX1 factor_b_reg_3_ ( .D(N129), .CLK(clk), .RSTB(rst_n), .Q(factor_b[3])
         );
  DFFARX1 factor_b_reg_2_ ( .D(N127), .CLK(clk), .RSTB(rst_n), .Q(factor_b[2])
         );
  DFFARX1 factor_b_reg_1_ ( .D(N129), .CLK(clk), .RSTB(rst_n), .Q(factor_b[1])
         );
  DFFASX1 factor_b_reg_0_ ( .D(n116), .CLK(clk), .SETB(rst_n), .QN(factor_b[0]) );
  DFFX1 factor_c_reg_31_ ( .D(n73), .CLK(clk), .Q(factor_c[31]) );
  DFFX1 factor_c_reg_29_ ( .D(n72), .CLK(clk), .Q(factor_c[29]) );
  DFFX1 factor_c_reg_28_ ( .D(n71), .CLK(clk), .Q(factor_c[28]) );
  DFFX1 factor_c_reg_27_ ( .D(n70), .CLK(clk), .Q(factor_c[27]) );
  DFFX1 factor_c_reg_26_ ( .D(n69), .CLK(clk), .Q(factor_c[26]) );
  DFFX1 factor_c_reg_25_ ( .D(n68), .CLK(clk), .Q(factor_c[25]) );
  DFFX1 factor_c_reg_24_ ( .D(n67), .CLK(clk), .Q(factor_c[24]) );
  DFFX1 factor_c_reg_23_ ( .D(n66), .CLK(clk), .Q(factor_c[23]) );
  DFFX1 factor_c_reg_22_ ( .D(n65), .CLK(clk), .Q(factor_c[22]) );
  DFFX1 factor_c_reg_21_ ( .D(n64), .CLK(clk), .Q(factor_c[21]) );
  DFFX1 factor_c_reg_19_ ( .D(n63), .CLK(clk), .Q(factor_c[19]) );
  DFFX1 factor_c_reg_18_ ( .D(n62), .CLK(clk), .Q(factor_c[18]) );
  DFFX1 factor_c_reg_17_ ( .D(n61), .CLK(clk), .Q(factor_c[17]) );
  DFFX1 factor_c_reg_16_ ( .D(n60), .CLK(clk), .Q(factor_c[16]) );
  DFFX1 factor_c_reg_15_ ( .D(n59), .CLK(clk), .Q(factor_c[15]) );
  DFFX1 factor_c_reg_14_ ( .D(n58), .CLK(clk), .Q(factor_c[14]) );
  DFFX1 factor_c_reg_13_ ( .D(n57), .CLK(clk), .Q(factor_c[13]) );
  DFFX1 factor_c_reg_11_ ( .D(n56), .CLK(clk), .Q(factor_c[11]) );
  DFFX1 factor_c_reg_10_ ( .D(n55), .CLK(clk), .Q(factor_c[10]) );
  DFFX1 factor_c_reg_9_ ( .D(n54), .CLK(clk), .Q(factor_c[9]) );
  DFFX1 factor_c_reg_8_ ( .D(n53), .CLK(clk), .Q(factor_c[8]) );
  DFFX1 factor_c_reg_7_ ( .D(n52), .CLK(clk), .Q(factor_c[7]) );
  DFFX1 factor_c_reg_6_ ( .D(n51), .CLK(clk), .Q(factor_c[6]) );
  DFFX1 factor_c_reg_5_ ( .D(n50), .CLK(clk), .Q(factor_c[5]) );
  DFFX1 factor_c_reg_4_ ( .D(n49), .CLK(clk), .Q(factor_c[4]) );
  DFFX1 factor_c_reg_3_ ( .D(n48), .CLK(clk), .Q(factor_c[3]) );
  DFFX1 factor_c_reg_2_ ( .D(n47), .CLK(clk), .Q(factor_c[2]) );
  DFFX1 factor_c_reg_0_ ( .D(n46), .CLK(clk), .Q(factor_c[0]) );
  DFFX1 factor_d_reg_31_ ( .D(n45), .CLK(clk), .Q(factor_d[31]) );
  DFFX1 factor_d_reg_29_ ( .D(n44), .CLK(clk), .Q(factor_d[29]) );
  DFFX1 factor_d_reg_25_ ( .D(n43), .CLK(clk), .Q(factor_d[25]) );
  DFFX1 factor_d_reg_24_ ( .D(n42), .CLK(clk), .Q(factor_d[24]) );
  DFFX1 factor_d_reg_22_ ( .D(n41), .CLK(clk), .Q(factor_d[22]) );
  DFFX1 factor_d_reg_21_ ( .D(n40), .CLK(clk), .Q(factor_d[21]) );
  DFFX1 factor_d_reg_20_ ( .D(n39), .CLK(clk), .Q(factor_d[20]) );
  DFFX1 factor_d_reg_19_ ( .D(n38), .CLK(clk), .Q(factor_d[19]) );
  DFFX1 factor_d_reg_18_ ( .D(n37), .CLK(clk), .Q(factor_d[18]) );
  DFFX1 factor_d_reg_17_ ( .D(n36), .CLK(clk), .Q(factor_d[17]) );
  DFFX1 factor_d_reg_16_ ( .D(n35), .CLK(clk), .Q(factor_d[16]) );
  DFFX1 factor_d_reg_15_ ( .D(n34), .CLK(clk), .Q(factor_d[15]) );
  DFFX1 factor_d_reg_14_ ( .D(n33), .CLK(clk), .Q(factor_d[14]) );
  DFFX1 factor_d_reg_13_ ( .D(n32), .CLK(clk), .Q(factor_d[13]) );
  DFFX1 factor_d_reg_12_ ( .D(n31), .CLK(clk), .Q(factor_d[12]) );
  DFFX1 factor_d_reg_11_ ( .D(n30), .CLK(clk), .Q(factor_d[11]) );
  DFFX1 factor_d_reg_10_ ( .D(n29), .CLK(clk), .Q(factor_d[10]) );
  DFFX1 factor_d_reg_9_ ( .D(n28), .CLK(clk), .Q(factor_d[9]) );
  DFFX1 factor_d_reg_8_ ( .D(n27), .CLK(clk), .Q(factor_d[8]) );
  DFFX1 factor_d_reg_7_ ( .D(n26), .CLK(clk), .Q(factor_d[7]) );
  DFFX1 factor_d_reg_6_ ( .D(n25), .CLK(clk), .Q(factor_d[6]) );
  DFFX1 factor_d_reg_5_ ( .D(n24), .CLK(clk), .Q(factor_d[5]) );
  DFFX1 factor_d_reg_4_ ( .D(n23), .CLK(clk), .Q(factor_d[4]) );
  DFFX1 factor_d_reg_3_ ( .D(n22), .CLK(clk), .Q(factor_d[3]) );
  DFFX1 factor_d_reg_2_ ( .D(n21), .CLK(clk), .Q(factor_d[2]) );
  DFFX1 factor_d_reg_1_ ( .D(n20), .CLK(clk), .Q(factor_d[1]) );
  DFFX1 factor_d_reg_0_ ( .D(n19), .CLK(clk), .Q(factor_d[0]) );
  INVX1 U3 ( .INP(rst_n), .ZN(n18) );
  NAND2X0 U4 ( .IN1(n9), .IN2(n10), .QN(n84) );
  NAND2X0 U5 ( .IN1(n5), .IN2(n6), .QN(n102) );
  NAND2X0 U6 ( .IN1(n119), .IN2(n132), .QN(n12) );
  NAND2X0 U7 ( .IN1(n89), .IN2(n136), .QN(n132) );
  NAND2X0 U8 ( .IN1(n7), .IN2(n8), .QN(n136) );
  NAND2X0 U9 ( .IN1(n141), .IN2(n130), .QN(n138) );
  NAND2X0 U10 ( .IN1(n124), .IN2(n123), .QN(n125) );
  NAND2X0 U11 ( .IN1(n74), .IN2(n115), .QN(N131) );
  NAND2X0 U12 ( .IN1(n116), .IN2(n74), .QN(N130) );
  NAND2X0 U13 ( .IN1(n78), .IN2(n115), .QN(N129) );
  NAND2X0 U14 ( .IN1(n80), .IN2(n115), .QN(N132) );
  NAND2X0 U15 ( .IN1(n79), .IN2(N124), .QN(n74) );
  NAND2X0 U16 ( .IN1(n75), .IN2(n115), .QN(N135) );
  NAND2X0 U17 ( .IN1(n116), .IN2(n145), .QN(N127) );
  NAND2X0 U18 ( .IN1(n116), .IN2(n75), .QN(N134) );
  NAND2X0 U19 ( .IN1(n116), .IN2(n115), .QN(N136) );
  NAND2X0 U20 ( .IN1(n127), .IN2(n126), .QN(n128) );
  NAND2X0 U21 ( .IN1(n131), .IN2(n130), .QN(n134) );
  NAND2X0 U22 ( .IN1(n135), .IN2(n17), .QN(n139) );
  NAND2X0 U23 ( .IN1(n143), .IN2(n142), .QN(N55) );
  NAND2X0 U24 ( .IN1(n141), .IN2(n140), .QN(n143) );
  NAND2X0 U25 ( .IN1(n1), .IN2(n3), .QN(n144) );
  NOR2X0 U26 ( .IN1(n18), .IN2(n75), .QN(n154) );
  INVX0 U27 ( .INP(n145), .ZN(N124) );
  NAND2X0 U28 ( .IN1(case_num[1]), .IN2(n77), .QN(n145) );
  NOR2X0 U29 ( .IN1(n18), .IN2(n116), .QN(n155) );
  NAND3X0 U30 ( .IN1(n151), .IN2(case_num[0]), .IN3(n77), .QN(n116) );
  NOR2X0 U31 ( .IN1(n11), .IN2(n12), .QN(n120) );
  NAND2X0 U32 ( .IN1(factor_input[1]), .IN2(n101), .QN(n6) );
  NOR2X0 U33 ( .IN1(factor_input[6]), .IN2(n100), .QN(n5) );
  NOR2X0 U34 ( .IN1(n133), .IN2(n127), .QN(n11) );
  NOR2X0 U35 ( .IN1(n13), .IN2(n14), .QN(n127) );
  NAND2X0 U36 ( .IN1(n96), .IN2(factor_input[19]), .QN(n14) );
  NOR2X0 U37 ( .IN1(n97), .IN2(factor_input[18]), .QN(n13) );
  NAND2X0 U38 ( .IN1(factor_input[20]), .IN2(n87), .QN(n8) );
  NAND2X0 U39 ( .IN1(factor_input[7]), .IN2(n83), .QN(n10) );
  NOR2X0 U40 ( .IN1(factor_input[9]), .IN2(factor_input[8]), .QN(n9) );
  NOR2X0 U41 ( .IN1(factor_input[22]), .IN2(factor_input[21]), .QN(n7) );
  OA21X1 U42 ( .IN1(case_num[1]), .IN2(n144), .IN3(n77), .Q(N137) );
  INVX0 U43 ( .INP(factor_input[15]), .ZN(n15) );
  INVX0 U44 ( .INP(factor_input[16]), .ZN(n16) );
  INVX0 U45 ( .INP(factor_input[30]), .ZN(n17) );
  INVX0 U46 ( .INP(factor_input[31]), .ZN(n76) );
  MUX21X1 U47 ( .IN1(n1), .IN2(case_num[2]), .S(case_num[0]), .Q(n79) );
  NAND3X0 U48 ( .IN1(case_num[2]), .IN2(n77), .IN3(n2), .QN(n115) );
  NOR2X0 U49 ( .IN1(case_num[2]), .IN2(case_num[1]), .QN(n151) );
  INVX0 U50 ( .INP(N130), .ZN(n78) );
  OR2X1 U51 ( .IN1(n79), .IN2(n145), .Q(n75) );
  INVX0 U52 ( .INP(N134), .ZN(n80) );
  OA221X1 U53 ( .IN1(case_num[1]), .IN2(case_num[0]), .IN3(n2), .IN4(
        case_num[2]), .IN5(n77), .Q(N139) );
  OR4X1 U54 ( .IN1(factor_input[24]), .IN2(factor_input[25]), .IN3(
        factor_input[23]), .IN4(factor_input[27]), .Q(n81) );
  NOR4X0 U55 ( .IN1(factor_input[26]), .IN2(factor_input[28]), .IN3(
        factor_input[29]), .IN4(n81), .QN(n124) );
  NAND2X0 U56 ( .IN1(n124), .IN2(factor_input[30]), .QN(n122) );
  INVX0 U57 ( .INP(n122), .ZN(n131) );
  AND4X1 U58 ( .IN1(factor_input[28]), .IN2(factor_input[29]), .IN3(
        factor_input[24]), .IN4(factor_input[25]), .Q(n82) );
  NAND4X0 U59 ( .IN1(factor_input[27]), .IN2(factor_input[26]), .IN3(n82), 
        .IN4(n17), .QN(n135) );
  INVX0 U60 ( .INP(n135), .ZN(n98) );
  NOR2X0 U61 ( .IN1(factor_input[23]), .IN2(n135), .QN(n89) );
  INVX0 U62 ( .INP(n89), .ZN(n88) );
  NOR3X0 U63 ( .IN1(factor_input[12]), .IN2(factor_input[13]), .IN3(
        factor_input[14]), .QN(n112) );
  AO221X1 U64 ( .IN1(factor_input[5]), .IN2(factor_input[3]), .IN3(
        factor_input[5]), .IN4(factor_input[4]), .IN5(factor_input[6]), .Q(n83) );
  NAND3X0 U65 ( .IN1(factor_input[10]), .IN2(factor_input[11]), .IN3(n84), 
        .QN(n85) );
  NAND4X0 U66 ( .IN1(n112), .IN2(n16), .IN3(n15), .IN4(n85), .QN(n86) );
  AO221X1 U67 ( .IN1(factor_input[18]), .IN2(factor_input[17]), .IN3(
        factor_input[18]), .IN4(n86), .IN5(factor_input[19]), .Q(n87) );
  OA22X1 U68 ( .IN1(n131), .IN2(n98), .IN3(n88), .IN4(n136), .Q(n121) );
  OA21X1 U69 ( .IN1(factor_input[9]), .IN2(factor_input[10]), .IN3(
        factor_input[11]), .Q(n93) );
  NAND4X0 U70 ( .IN1(factor_input[5]), .IN2(factor_input[2]), .IN3(
        factor_input[3]), .IN4(factor_input[4]), .QN(n99) );
  NAND2X0 U71 ( .IN1(factor_input[6]), .IN2(factor_input[7]), .QN(n108) );
  NOR2X0 U72 ( .IN1(n99), .IN2(n108), .QN(n90) );
  AO221X1 U73 ( .IN1(n90), .IN2(factor_input[1]), .IN3(n90), .IN4(
        factor_input[0]), .IN5(factor_input[10]), .Q(n92) );
  OR3X1 U74 ( .IN1(factor_input[12]), .IN2(factor_input[13]), .IN3(
        factor_input[15]), .Q(n91) );
  AO221X1 U75 ( .IN1(n93), .IN2(factor_input[8]), .IN3(n93), .IN4(n92), .IN5(
        n91), .Q(n95) );
  OR2X1 U76 ( .IN1(factor_input[14]), .IN2(factor_input[15]), .Q(n94) );
  AND4X1 U77 ( .IN1(factor_input[16]), .IN2(factor_input[17]), .IN3(n95), 
        .IN4(n94), .Q(n97) );
  AND3X1 U78 ( .IN1(factor_input[20]), .IN2(factor_input[21]), .IN3(
        factor_input[22]), .Q(n96) );
  NAND2X0 U79 ( .IN1(factor_input[23]), .IN2(n98), .QN(n133) );
  OR4X1 U80 ( .IN1(factor_input[13]), .IN2(factor_input[16]), .IN3(
        factor_input[14]), .IN4(factor_input[15]), .Q(n104) );
  INVX0 U81 ( .INP(n99), .ZN(n101) );
  OR2X1 U82 ( .IN1(factor_input[7]), .IN2(factor_input[8]), .Q(n100) );
  AO221X1 U83 ( .IN1(factor_input[10]), .IN2(factor_input[9]), .IN3(
        factor_input[10]), .IN4(n102), .IN5(factor_input[11]), .Q(n103) );
  OA221X1 U84 ( .IN1(n104), .IN2(n103), .IN3(n104), .IN4(factor_input[12]), 
        .IN5(factor_input[17]), .Q(n105) );
  AO221X1 U85 ( .IN1(factor_input[19]), .IN2(factor_input[18]), .IN3(
        factor_input[19]), .IN4(n105), .IN5(factor_input[21]), .Q(n106) );
  OA21X1 U86 ( .IN1(factor_input[20]), .IN2(n106), .IN3(factor_input[22]), .Q(
        n140) );
  AND3X1 U87 ( .IN1(factor_input[2]), .IN2(factor_input[1]), .IN3(
        factor_input[0]), .Q(n107) );
  NOR4X0 U88 ( .IN1(factor_input[5]), .IN2(factor_input[3]), .IN3(
        factor_input[4]), .IN4(n107), .QN(n109) );
  NOR2X0 U89 ( .IN1(n109), .IN2(n108), .QN(n111) );
  OR4X1 U90 ( .IN1(factor_input[11]), .IN2(factor_input[10]), .IN3(
        factor_input[13]), .IN4(factor_input[14]), .Q(n110) );
  AOI221X1 U91 ( .IN1(factor_input[9]), .IN2(factor_input[8]), .IN3(
        factor_input[9]), .IN4(n111), .IN5(n110), .QN(n113) );
  NOR3X0 U92 ( .IN1(n15), .IN2(n113), .IN3(n112), .QN(n114) );
  OA21X1 U93 ( .IN1(factor_input[16]), .IN2(n114), .IN3(factor_input[17]), .Q(
        n117) );
  AO21X1 U94 ( .IN1(factor_input[18]), .IN2(n117), .IN3(factor_input[19]), .Q(
        n118) );
  NAND4X0 U95 ( .IN1(factor_input[21]), .IN2(factor_input[20]), .IN3(
        factor_input[22]), .IN4(n118), .QN(n123) );
  NAND3X0 U96 ( .IN1(n131), .IN2(n140), .IN3(n123), .QN(n119) );
  MUX21X1 U97 ( .IN1(n121), .IN2(n120), .S(factor_input[31]), .Q(n129) );
  NOR2X0 U98 ( .IN1(factor_input[31]), .IN2(n122), .QN(n141) );
  INVX0 U99 ( .INP(n140), .ZN(n130) );
  NAND3X0 U100 ( .IN1(n125), .IN2(n76), .IN3(factor_input[30]), .QN(n142) );
  NOR2X0 U101 ( .IN1(factor_input[31]), .IN2(n133), .QN(n126) );
  NAND4X0 U102 ( .IN1(n129), .IN2(n138), .IN3(n142), .IN4(n128), .QN(N52) );
  NAND3X0 U103 ( .IN1(n134), .IN2(n133), .IN3(n132), .QN(N53) );
  AO221X1 U104 ( .IN1(factor_input[31]), .IN2(factor_input[23]), .IN3(
        factor_input[31]), .IN4(n136), .IN5(n135), .Q(n137) );
  NAND3X0 U105 ( .IN1(n139), .IN2(n138), .IN3(n137), .QN(N54) );
  MUX21X1 U106 ( .IN1(N130), .IN2(factor_d[4]), .S(n18), .Q(n23) );
  MUX21X1 U107 ( .IN1(N134), .IN2(factor_d[6]), .S(n18), .Q(n25) );
  MUX21X1 U108 ( .IN1(N134), .IN2(factor_d[16]), .S(n18), .Q(n35) );
  MUX21X1 U109 ( .IN1(N130), .IN2(factor_d[19]), .S(n18), .Q(n38) );
  MUX21X1 U110 ( .IN1(n115), .IN2(factor_d[29]), .S(n18), .Q(n44) );
  MUX21X1 U111 ( .IN1(N134), .IN2(factor_c[0]), .S(n18), .Q(n46) );
  MUX21X1 U112 ( .IN1(N130), .IN2(factor_c[5]), .S(n18), .Q(n50) );
  MUX21X1 U113 ( .IN1(N130), .IN2(factor_c[8]), .S(n18), .Q(n53) );
  MUX21X1 U114 ( .IN1(N130), .IN2(factor_c[11]), .S(n18), .Q(n56) );
  MUX21X1 U115 ( .IN1(N134), .IN2(factor_c[13]), .S(n18), .Q(n57) );
  MUX21X1 U116 ( .IN1(N134), .IN2(factor_c[14]), .S(n18), .Q(n58) );
  MUX21X1 U117 ( .IN1(N130), .IN2(factor_c[15]), .S(n18), .Q(n59) );
  MUX21X1 U118 ( .IN1(N134), .IN2(factor_c[18]), .S(n18), .Q(n62) );
  MUX21X1 U119 ( .IN1(N137), .IN2(factor_c[25]), .S(n18), .Q(n68) );
  MUX21X1 U120 ( .IN1(N137), .IN2(factor_c[26]), .S(n18), .Q(n69) );
  MUX21X1 U121 ( .IN1(N137), .IN2(factor_c[27]), .S(n18), .Q(n70) );
  MUX21X1 U122 ( .IN1(N137), .IN2(factor_c[28]), .S(n18), .Q(n71) );
  MUX21X1 U123 ( .IN1(N137), .IN2(factor_c[29]), .S(n18), .Q(n72) );
  MUX21X1 U124 ( .IN1(N124), .IN2(factor_d[0]), .S(n18), .Q(n19) );
  AO21X1 U125 ( .IN1(n18), .IN2(factor_d[1]), .IN3(n155), .Q(n20) );
  AO21X1 U126 ( .IN1(n18), .IN2(factor_d[2]), .IN3(n155), .Q(n21) );
  MUX21X1 U127 ( .IN1(N127), .IN2(factor_d[3]), .S(n18), .Q(n22) );
  NOR2X0 U128 ( .IN1(n18), .IN2(n74), .QN(n153) );
  AO21X1 U129 ( .IN1(n18), .IN2(factor_d[5]), .IN3(n153), .Q(n24) );
  MUX21X1 U130 ( .IN1(N124), .IN2(factor_d[7]), .S(n18), .Q(n26) );
  AO21X1 U131 ( .IN1(n18), .IN2(factor_d[8]), .IN3(n153), .Q(n27) );
  MUX21X1 U132 ( .IN1(N124), .IN2(factor_d[9]), .S(n18), .Q(n28) );
  AO21X1 U133 ( .IN1(n18), .IN2(factor_d[10]), .IN3(n155), .Q(n29) );
  AO21X1 U134 ( .IN1(n18), .IN2(factor_d[11]), .IN3(n154), .Q(n30) );
  AO21X1 U135 ( .IN1(n18), .IN2(factor_d[12]), .IN3(n153), .Q(n31) );
  AO21X1 U136 ( .IN1(n18), .IN2(factor_d[13]), .IN3(n154), .Q(n32) );
  MUX21X1 U137 ( .IN1(N127), .IN2(factor_d[14]), .S(n18), .Q(n33) );
  AO21X1 U138 ( .IN1(n18), .IN2(factor_d[15]), .IN3(n153), .Q(n34) );
  AO21X1 U139 ( .IN1(n18), .IN2(factor_d[17]), .IN3(n154), .Q(n36) );
  AO21X1 U140 ( .IN1(n18), .IN2(factor_d[18]), .IN3(n154), .Q(n37) );
  AO21X1 U141 ( .IN1(n18), .IN2(factor_d[20]), .IN3(n155), .Q(n39) );
  MUX21X1 U142 ( .IN1(N124), .IN2(factor_d[21]), .S(n18), .Q(n40) );
  MUX21X1 U143 ( .IN1(N124), .IN2(factor_d[22]), .S(n18), .Q(n41) );
  NOR2X0 U144 ( .IN1(case_num[0]), .IN2(n2), .QN(n150) );
  NOR2X0 U145 ( .IN1(n151), .IN2(n4), .QN(N128) );
  INVX0 U146 ( .INP(N128), .ZN(n147) );
  AO221X1 U147 ( .IN1(case_num[2]), .IN2(n150), .IN3(n1), .IN4(case_num[0]), 
        .IN5(n147), .Q(n146) );
  MUX21X1 U148 ( .IN1(n146), .IN2(factor_d[24]), .S(n18), .Q(n42) );
  NOR2X0 U149 ( .IN1(n3), .IN2(n1), .QN(n148) );
  AO221X1 U150 ( .IN1(n1), .IN2(n3), .IN3(n148), .IN4(case_num[1]), .IN5(n147), 
        .Q(n149) );
  MUX21X1 U151 ( .IN1(n149), .IN2(factor_d[25]), .S(n18), .Q(n43) );
  OA21X1 U152 ( .IN1(n151), .IN2(n150), .IN3(rst_n), .Q(n152) );
  AO22X1 U153 ( .IN1(n18), .IN2(factor_d[31]), .IN3(n77), .IN4(n152), .Q(n45)
         );
  MUX21X1 U154 ( .IN1(N127), .IN2(factor_c[2]), .S(n18), .Q(n47) );
  AO21X1 U155 ( .IN1(n18), .IN2(factor_c[3]), .IN3(n154), .Q(n48) );
  AO21X1 U156 ( .IN1(n18), .IN2(factor_c[4]), .IN3(n154), .Q(n49) );
  AO21X1 U157 ( .IN1(n18), .IN2(factor_c[6]), .IN3(n155), .Q(n51) );
  AO21X1 U158 ( .IN1(n18), .IN2(factor_c[7]), .IN3(n154), .Q(n52) );
  MUX21X1 U159 ( .IN1(N127), .IN2(factor_c[9]), .S(n18), .Q(n54) );
  AO21X1 U160 ( .IN1(n18), .IN2(factor_c[10]), .IN3(n154), .Q(n55) );
  AO21X1 U161 ( .IN1(n18), .IN2(factor_c[16]), .IN3(n153), .Q(n60) );
  AO21X1 U162 ( .IN1(n18), .IN2(factor_c[17]), .IN3(n154), .Q(n61) );
  AO21X1 U163 ( .IN1(n18), .IN2(factor_c[19]), .IN3(n155), .Q(n63) );
  AO21X1 U164 ( .IN1(n18), .IN2(factor_c[21]), .IN3(n154), .Q(n64) );
  AO21X1 U165 ( .IN1(n18), .IN2(factor_c[22]), .IN3(n155), .Q(n65) );
  MUX21X1 U166 ( .IN1(N135), .IN2(factor_c[23]), .S(n18), .Q(n66) );
  MUX21X1 U167 ( .IN1(N128), .IN2(factor_c[24]), .S(n18), .Q(n67) );
  AO21X1 U168 ( .IN1(n18), .IN2(factor_c[31]), .IN3(n155), .Q(n73) );
endmodule


module add_33 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_34 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_35 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_36 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_37 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_38 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_39 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_40 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_41 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_42 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_43 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_44 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_45 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_46 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_47 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_48 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_49 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_50 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_51 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_52 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_53 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_54 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_55 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_56 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(b), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(b), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module adder24_1 ( clk, rst_n, a, b, cin, out );
  input [23:0] a;
  input [23:0] b;
  output [24:0] out;
  input clk, rst_n, cin;
  wire   c_tmp;
  wire   [24:0] s;
  wire   [22:0] c;

  add_56 add_01 ( .s(s[0]), .a(a[0]), .b(b[0]), .ci(1'b0), .co(c[0]) );
  add_55 add_02 ( .s(s[1]), .a(a[1]), .b(b[1]), .ci(c[0]), .co(c[1]) );
  add_54 add_03 ( .s(s[2]), .a(a[2]), .b(b[2]), .ci(c[1]), .co(c[2]) );
  add_53 add_04 ( .s(s[3]), .a(a[3]), .b(b[3]), .ci(c[2]), .co(c[3]) );
  add_52 add_05 ( .s(s[4]), .a(a[4]), .b(b[4]), .ci(c[3]), .co(c[4]) );
  add_51 add_06 ( .s(s[5]), .a(a[5]), .b(b[5]), .ci(c[4]), .co(c[5]) );
  add_50 add_07 ( .s(s[6]), .a(a[6]), .b(b[6]), .ci(c[5]), .co(c[6]) );
  add_49 add_08 ( .s(s[7]), .a(a[7]), .b(b[7]), .ci(c[6]), .co(c[7]) );
  add_48 add_09 ( .s(s[8]), .a(a[8]), .b(b[8]), .ci(c[7]), .co(c[8]) );
  add_47 add_10 ( .s(s[9]), .a(a[9]), .b(b[9]), .ci(c[8]), .co(c[9]) );
  add_46 add_11 ( .s(s[10]), .a(a[10]), .b(b[10]), .ci(c[9]), .co(c[10]) );
  add_45 add_12 ( .s(s[11]), .a(a[11]), .b(b[11]), .ci(c_tmp), .co(c[11]) );
  add_44 add_13 ( .s(s[12]), .a(a[12]), .b(b[12]), .ci(c[11]), .co(c[12]) );
  add_43 add_14 ( .s(s[13]), .a(a[13]), .b(b[13]), .ci(c[12]), .co(c[13]) );
  add_42 add_15 ( .s(s[14]), .a(a[14]), .b(b[14]), .ci(c[13]), .co(c[14]) );
  add_41 add_16 ( .s(s[15]), .a(a[15]), .b(b[15]), .ci(c[14]), .co(c[15]) );
  add_40 add_17 ( .s(s[16]), .a(a[16]), .b(b[16]), .ci(c[15]), .co(c[16]) );
  add_39 add_18 ( .s(s[17]), .a(a[17]), .b(b[17]), .ci(c[16]), .co(c[17]) );
  add_38 add_19 ( .s(s[18]), .a(a[18]), .b(b[18]), .ci(c[17]), .co(c[18]) );
  add_37 add_20 ( .s(s[19]), .a(a[19]), .b(b[19]), .ci(c[18]), .co(c[19]) );
  add_36 add_21 ( .s(s[20]), .a(a[20]), .b(b[20]), .ci(c[19]), .co(c[20]) );
  add_35 add_22 ( .s(s[21]), .a(a[21]), .b(b[21]), .ci(c[20]), .co(c[21]) );
  add_34 add_23 ( .s(s[22]), .a(a[22]), .b(b[22]), .ci(c[21]), .co(c[22]) );
  add_33 add_24 ( .s(s[23]), .a(a[23]), .b(b[23]), .ci(c[22]), .co(s[24]) );
  DFFARX1 out_reg_10_ ( .D(s[10]), .CLK(clk), .RSTB(rst_n), .Q(out[10]) );
  DFFARX1 out_reg_9_ ( .D(s[9]), .CLK(clk), .RSTB(rst_n), .Q(out[9]) );
  DFFARX1 out_reg_8_ ( .D(s[8]), .CLK(clk), .RSTB(rst_n), .Q(out[8]) );
  DFFARX1 out_reg_7_ ( .D(s[7]), .CLK(clk), .RSTB(rst_n), .Q(out[7]) );
  DFFARX1 out_reg_6_ ( .D(s[6]), .CLK(clk), .RSTB(rst_n), .Q(out[6]) );
  DFFARX1 out_reg_5_ ( .D(s[5]), .CLK(clk), .RSTB(rst_n), .Q(out[5]) );
  DFFARX1 out_reg_4_ ( .D(s[4]), .CLK(clk), .RSTB(rst_n), .Q(out[4]) );
  DFFARX1 out_reg_3_ ( .D(s[3]), .CLK(clk), .RSTB(rst_n), .Q(out[3]) );
  DFFARX1 out_reg_2_ ( .D(s[2]), .CLK(clk), .RSTB(rst_n), .Q(out[2]) );
  DFFARX1 out_reg_1_ ( .D(s[1]), .CLK(clk), .RSTB(rst_n), .Q(out[1]) );
  DFFARX1 out_reg_0_ ( .D(s[0]), .CLK(clk), .RSTB(rst_n), .Q(out[0]) );
  DFFARX1 c_tmp_reg ( .D(c[10]), .CLK(clk), .RSTB(rst_n), .Q(c_tmp) );
  DFFARX1 out_reg_24_ ( .D(s[24]), .CLK(clk), .RSTB(rst_n), .Q(out[24]) );
  DFFARX1 out_reg_23_ ( .D(s[23]), .CLK(clk), .RSTB(rst_n), .Q(out[23]) );
  DFFARX1 out_reg_22_ ( .D(s[22]), .CLK(clk), .RSTB(rst_n), .Q(out[22]) );
  DFFARX1 out_reg_21_ ( .D(s[21]), .CLK(clk), .RSTB(rst_n), .Q(out[21]) );
  DFFARX1 out_reg_20_ ( .D(s[20]), .CLK(clk), .RSTB(rst_n), .Q(out[20]) );
  DFFARX1 out_reg_19_ ( .D(s[19]), .CLK(clk), .RSTB(rst_n), .Q(out[19]) );
  DFFARX1 out_reg_18_ ( .D(s[18]), .CLK(clk), .RSTB(rst_n), .Q(out[18]) );
  DFFARX1 out_reg_17_ ( .D(s[17]), .CLK(clk), .RSTB(rst_n), .Q(out[17]) );
  DFFARX1 out_reg_16_ ( .D(s[16]), .CLK(clk), .RSTB(rst_n), .Q(out[16]) );
  DFFARX1 out_reg_15_ ( .D(s[15]), .CLK(clk), .RSTB(rst_n), .Q(out[15]) );
  DFFARX1 out_reg_14_ ( .D(s[14]), .CLK(clk), .RSTB(rst_n), .Q(out[14]) );
  DFFARX1 out_reg_13_ ( .D(s[13]), .CLK(clk), .RSTB(rst_n), .Q(out[13]) );
  DFFARX1 out_reg_12_ ( .D(s[12]), .CLK(clk), .RSTB(rst_n), .Q(out[12]) );
  DFFARX1 out_reg_11_ ( .D(s[11]), .CLK(clk), .RSTB(rst_n), .Q(out[11]) );
endmodule


module add_57 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_58 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_59 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_60 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_61 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_62 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_63 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_64 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_65 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_66 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_67 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_68 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_69 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_70 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_71 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_72 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_73 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_74 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_75 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_76 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_77 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_78 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_79 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_80 ( s, a, ci, co, b_BAR );
  input a, ci, b_BAR;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(b_BAR), .IN2(n1), .QN(co) );
  INVX0 U2 ( .INP(a), .ZN(n1) );
  MUX21X1 U3 ( .IN1(a), .IN2(n1), .S(b_BAR), .Q(s) );
endmodule


module adder24_2 ( clk, rst_n, a, b, cin, out );
  input [23:0] a;
  input [23:0] b;
  output [24:0] out;
  input clk, rst_n, cin;
  wire   c_tmp, n_1_net_, n_2_net_, n_3_net_, n_4_net_, n_5_net_, n_6_net_,
         n_7_net_, n_8_net_, n_9_net_, n_10_net_, n_11_net_, n_12_net_,
         n_13_net_, n_14_net_, n_15_net_, n_16_net_, n_17_net_, n_18_net_,
         n_19_net_, n_20_net_, n_21_net_, n_22_net_, n_23_net_;
  wire   [24:0] s;
  wire   [23:0] c;

  add_80 add_01 ( .s(s[0]), .a(a[0]), .ci(1'b1), .co(c[0]), .b_BAR(b[0]) );
  add_79 add_02 ( .s(s[1]), .a(a[1]), .b(n_1_net_), .ci(c[0]), .co(c[1]) );
  add_78 add_03 ( .s(s[2]), .a(a[2]), .b(n_2_net_), .ci(c[1]), .co(c[2]) );
  add_77 add_04 ( .s(s[3]), .a(a[3]), .b(n_3_net_), .ci(c[2]), .co(c[3]) );
  add_76 add_05 ( .s(s[4]), .a(a[4]), .b(n_4_net_), .ci(c[3]), .co(c[4]) );
  add_75 add_06 ( .s(s[5]), .a(a[5]), .b(n_5_net_), .ci(c[4]), .co(c[5]) );
  add_74 add_07 ( .s(s[6]), .a(a[6]), .b(n_6_net_), .ci(c[5]), .co(c[6]) );
  add_73 add_08 ( .s(s[7]), .a(a[7]), .b(n_7_net_), .ci(c[6]), .co(c[7]) );
  add_72 add_09 ( .s(s[8]), .a(a[8]), .b(n_8_net_), .ci(c[7]), .co(c[8]) );
  add_71 add_10 ( .s(s[9]), .a(a[9]), .b(n_9_net_), .ci(c[8]), .co(c[9]) );
  add_70 add_11 ( .s(s[10]), .a(a[10]), .b(n_10_net_), .ci(c[9]), .co(c[10])
         );
  add_69 add_12 ( .s(s[11]), .a(a[11]), .b(n_11_net_), .ci(c_tmp), .co(c[11])
         );
  add_68 add_13 ( .s(s[12]), .a(a[12]), .b(n_12_net_), .ci(c[11]), .co(c[12])
         );
  add_67 add_14 ( .s(s[13]), .a(a[13]), .b(n_13_net_), .ci(c[12]), .co(c[13])
         );
  add_66 add_15 ( .s(s[14]), .a(a[14]), .b(n_14_net_), .ci(c[13]), .co(c[14])
         );
  add_65 add_16 ( .s(s[15]), .a(a[15]), .b(n_15_net_), .ci(c[14]), .co(c[15])
         );
  add_64 add_17 ( .s(s[16]), .a(a[16]), .b(n_16_net_), .ci(c[15]), .co(c[16])
         );
  add_63 add_18 ( .s(s[17]), .a(a[17]), .b(n_17_net_), .ci(c[16]), .co(c[17])
         );
  add_62 add_19 ( .s(s[18]), .a(a[18]), .b(n_18_net_), .ci(c[17]), .co(c[18])
         );
  add_61 add_20 ( .s(s[19]), .a(a[19]), .b(n_19_net_), .ci(c[18]), .co(c[19])
         );
  add_60 add_21 ( .s(s[20]), .a(a[20]), .b(n_20_net_), .ci(c[19]), .co(c[20])
         );
  add_59 add_22 ( .s(s[21]), .a(a[21]), .b(n_21_net_), .ci(c[20]), .co(c[21])
         );
  add_58 add_23 ( .s(s[22]), .a(a[22]), .b(n_22_net_), .ci(c[21]), .co(c[22])
         );
  add_57 add_24 ( .s(s[23]), .a(a[23]), .b(n_23_net_), .ci(c[22]), .co(c[23])
         );
  DFFARX1 out_reg_10_ ( .D(s[10]), .CLK(clk), .RSTB(rst_n), .Q(out[10]) );
  DFFARX1 out_reg_9_ ( .D(s[9]), .CLK(clk), .RSTB(rst_n), .Q(out[9]) );
  DFFARX1 out_reg_8_ ( .D(s[8]), .CLK(clk), .RSTB(rst_n), .Q(out[8]) );
  DFFARX1 out_reg_7_ ( .D(s[7]), .CLK(clk), .RSTB(rst_n), .Q(out[7]) );
  DFFARX1 out_reg_6_ ( .D(s[6]), .CLK(clk), .RSTB(rst_n), .Q(out[6]) );
  DFFARX1 out_reg_5_ ( .D(s[5]), .CLK(clk), .RSTB(rst_n), .Q(out[5]) );
  DFFARX1 out_reg_4_ ( .D(s[4]), .CLK(clk), .RSTB(rst_n), .Q(out[4]) );
  DFFARX1 out_reg_3_ ( .D(s[3]), .CLK(clk), .RSTB(rst_n), .Q(out[3]) );
  DFFARX1 out_reg_2_ ( .D(s[2]), .CLK(clk), .RSTB(rst_n), .Q(out[2]) );
  DFFARX1 out_reg_1_ ( .D(s[1]), .CLK(clk), .RSTB(rst_n), .Q(out[1]) );
  DFFARX1 out_reg_0_ ( .D(s[0]), .CLK(clk), .RSTB(rst_n), .Q(out[0]) );
  DFFARX1 c_tmp_reg ( .D(c[10]), .CLK(clk), .RSTB(rst_n), .Q(c_tmp) );
  DFFARX1 out_reg_24_ ( .D(s[24]), .CLK(clk), .RSTB(rst_n), .Q(out[24]) );
  DFFARX1 out_reg_23_ ( .D(s[23]), .CLK(clk), .RSTB(rst_n), .Q(out[23]) );
  DFFARX1 out_reg_22_ ( .D(s[22]), .CLK(clk), .RSTB(rst_n), .Q(out[22]) );
  DFFARX1 out_reg_21_ ( .D(s[21]), .CLK(clk), .RSTB(rst_n), .Q(out[21]) );
  DFFARX1 out_reg_20_ ( .D(s[20]), .CLK(clk), .RSTB(rst_n), .Q(out[20]) );
  DFFARX1 out_reg_19_ ( .D(s[19]), .CLK(clk), .RSTB(rst_n), .Q(out[19]) );
  DFFARX1 out_reg_18_ ( .D(s[18]), .CLK(clk), .RSTB(rst_n), .Q(out[18]) );
  DFFARX1 out_reg_17_ ( .D(s[17]), .CLK(clk), .RSTB(rst_n), .Q(out[17]) );
  DFFARX1 out_reg_16_ ( .D(s[16]), .CLK(clk), .RSTB(rst_n), .Q(out[16]) );
  DFFARX1 out_reg_15_ ( .D(s[15]), .CLK(clk), .RSTB(rst_n), .Q(out[15]) );
  DFFARX1 out_reg_14_ ( .D(s[14]), .CLK(clk), .RSTB(rst_n), .Q(out[14]) );
  DFFARX1 out_reg_13_ ( .D(s[13]), .CLK(clk), .RSTB(rst_n), .Q(out[13]) );
  DFFARX1 out_reg_12_ ( .D(s[12]), .CLK(clk), .RSTB(rst_n), .Q(out[12]) );
  DFFARX1 out_reg_11_ ( .D(s[11]), .CLK(clk), .RSTB(rst_n), .Q(out[11]) );
  INVX0 U3 ( .INP(b[1]), .ZN(n_1_net_) );
  INVX0 U4 ( .INP(b[2]), .ZN(n_2_net_) );
  INVX0 U5 ( .INP(b[3]), .ZN(n_3_net_) );
  INVX0 U6 ( .INP(b[4]), .ZN(n_4_net_) );
  INVX0 U7 ( .INP(b[5]), .ZN(n_5_net_) );
  INVX0 U8 ( .INP(b[6]), .ZN(n_6_net_) );
  INVX0 U9 ( .INP(b[7]), .ZN(n_7_net_) );
  INVX0 U10 ( .INP(b[8]), .ZN(n_8_net_) );
  INVX0 U11 ( .INP(b[9]), .ZN(n_9_net_) );
  INVX0 U12 ( .INP(b[10]), .ZN(n_10_net_) );
  INVX0 U13 ( .INP(c[23]), .ZN(s[24]) );
  INVX0 U14 ( .INP(b[11]), .ZN(n_11_net_) );
  INVX0 U15 ( .INP(b[12]), .ZN(n_12_net_) );
  INVX0 U16 ( .INP(b[13]), .ZN(n_13_net_) );
  INVX0 U17 ( .INP(b[14]), .ZN(n_14_net_) );
  INVX0 U18 ( .INP(b[15]), .ZN(n_15_net_) );
  INVX0 U19 ( .INP(b[16]), .ZN(n_16_net_) );
  INVX0 U20 ( .INP(b[17]), .ZN(n_17_net_) );
  INVX0 U21 ( .INP(b[18]), .ZN(n_18_net_) );
  INVX0 U22 ( .INP(b[19]), .ZN(n_19_net_) );
  INVX0 U23 ( .INP(b[20]), .ZN(n_20_net_) );
  INVX0 U24 ( .INP(b[21]), .ZN(n_21_net_) );
  INVX0 U25 ( .INP(b[22]), .ZN(n_22_net_) );
  INVX0 U26 ( .INP(b[23]), .ZN(n_23_net_) );
endmodule


module add_1 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  XNOR2X1 U1 ( .IN1(ci), .IN2(a), .Q(s) );
endmodule


module add_2 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_3 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_4 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_5 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_6 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_7 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_8 ( s, a, ci, co, b_BAR );
  input a, ci, b_BAR;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(b_BAR), .IN2(n1), .QN(co) );
  INVX0 U2 ( .INP(a), .ZN(n1) );
  MUX21X1 U3 ( .IN1(a), .IN2(n1), .S(b_BAR), .Q(s) );
endmodule


module adder8_1 ( out, a, b, cin );
  output [7:0] out;
  input [7:0] a;
  input [7:0] b;
  input cin;
  wire   n_1_net_, n_2_net_, n_4_net_;
  wire   [6:0] c;

  add_8 add_01 ( .s(out[0]), .a(a[0]), .ci(1'b1), .co(c[0]), .b_BAR(b[0]) );
  add_7 add_02 ( .s(out[1]), .a(a[1]), .b(n_1_net_), .ci(c[0]), .co(c[1]) );
  add_6 add_03 ( .s(out[2]), .a(a[2]), .b(n_2_net_), .ci(c[1]), .co(c[2]) );
  add_5 add_04 ( .s(out[3]), .a(a[3]), .b(1'b1), .ci(c[2]), .co(c[3]) );
  add_4 add_05 ( .s(out[4]), .a(a[4]), .b(n_4_net_), .ci(c[3]), .co(c[4]) );
  add_3 add_06 ( .s(out[5]), .a(a[5]), .b(1'b1), .ci(c[4]), .co(c[5]) );
  add_2 add_07 ( .s(out[6]), .a(a[6]), .b(1'b1), .ci(c[5]), .co(c[6]) );
  add_1 add_08 ( .s(out[7]), .a(a[7]), .b(1'b1), .ci(c[6]) );
  INVX0 U1 ( .INP(b[4]), .ZN(n_4_net_) );
  INVX0 U2 ( .INP(b[1]), .ZN(n_1_net_) );
  INVX0 U3 ( .INP(b[2]), .ZN(n_2_net_) );
endmodule


module add_9 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  XNOR2X1 U1 ( .IN1(ci), .IN2(a), .Q(s) );
endmodule


module add_10 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_11 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_12 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_13 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_14 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_15 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_16 ( s, a, ci, co, b_BAR );
  input a, ci, b_BAR;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(b_BAR), .IN2(n1), .QN(co) );
  INVX0 U2 ( .INP(a), .ZN(n1) );
  MUX21X1 U3 ( .IN1(a), .IN2(n1), .S(b_BAR), .Q(s) );
endmodule


module adder8_2 ( out, a, b, cin );
  output [7:0] out;
  input [7:0] a;
  input [7:0] b;
  input cin;
  wire   n_1_net_, n_2_net_, n_3_net_;
  wire   [6:0] c;

  add_16 add_01 ( .s(out[0]), .a(a[0]), .ci(1'b1), .co(c[0]), .b_BAR(b[0]) );
  add_15 add_02 ( .s(out[1]), .a(a[1]), .b(n_1_net_), .ci(c[0]), .co(c[1]) );
  add_14 add_03 ( .s(out[2]), .a(a[2]), .b(n_2_net_), .ci(c[1]), .co(c[2]) );
  add_13 add_04 ( .s(out[3]), .a(a[3]), .b(n_3_net_), .ci(c[2]), .co(c[3]) );
  add_12 add_05 ( .s(out[4]), .a(a[4]), .b(1'b1), .ci(c[3]), .co(c[4]) );
  add_11 add_06 ( .s(out[5]), .a(a[5]), .b(1'b1), .ci(c[4]), .co(c[5]) );
  add_10 add_07 ( .s(out[6]), .a(a[6]), .b(1'b1), .ci(c[5]), .co(c[6]) );
  add_9 add_08 ( .s(out[7]), .a(a[7]), .b(1'b1), .ci(c[6]) );
  INVX0 U1 ( .INP(b[1]), .ZN(n_1_net_) );
  INVX0 U2 ( .INP(b[2]), .ZN(n_2_net_) );
  INVX0 U3 ( .INP(b[3]), .ZN(n_3_net_) );
endmodule


module add_17 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  XNOR2X1 U1 ( .IN1(ci), .IN2(a), .Q(s) );
endmodule


module add_18 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_19 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_20 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_21 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_22 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_23 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_24 ( s, a, ci, co, b_BAR );
  input a, ci, b_BAR;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(b_BAR), .IN2(n1), .QN(co) );
  INVX0 U2 ( .INP(a), .ZN(n1) );
  MUX21X1 U3 ( .IN1(a), .IN2(n1), .S(b_BAR), .Q(s) );
endmodule


module adder8_3 ( out, a, b, cin );
  output [7:0] out;
  input [7:0] a;
  input [7:0] b;
  input cin;
  wire   n_1_net_, n_2_net_, n_3_net_;
  wire   [6:0] c;

  add_24 add_01 ( .s(out[0]), .a(a[0]), .ci(1'b1), .co(c[0]), .b_BAR(b[0]) );
  add_23 add_02 ( .s(out[1]), .a(a[1]), .b(n_1_net_), .ci(c[0]), .co(c[1]) );
  add_22 add_03 ( .s(out[2]), .a(a[2]), .b(n_2_net_), .ci(c[1]), .co(c[2]) );
  add_21 add_04 ( .s(out[3]), .a(a[3]), .b(n_3_net_), .ci(c[2]), .co(c[3]) );
  add_20 add_05 ( .s(out[4]), .a(a[4]), .b(1'b1), .ci(c[3]), .co(c[4]) );
  add_19 add_06 ( .s(out[5]), .a(a[5]), .b(1'b1), .ci(c[4]), .co(c[5]) );
  add_18 add_07 ( .s(out[6]), .a(a[6]), .b(1'b1), .ci(c[5]), .co(c[6]) );
  add_17 add_08 ( .s(out[7]), .a(a[7]), .b(1'b1), .ci(c[6]) );
  INVX0 U1 ( .INP(b[1]), .ZN(n_1_net_) );
  INVX0 U2 ( .INP(b[2]), .ZN(n_2_net_) );
  INVX0 U3 ( .INP(b[3]), .ZN(n_3_net_) );
endmodule


module add_25 ( s, a, b, co, ci_BAR );
  input a, b, ci_BAR;
  output s, co;


  XNOR2X1 U1 ( .IN1(a), .IN2(ci_BAR), .Q(s) );
endmodule


module add_26 ( s, a, b, ci, co_BAR );
  input a, b, ci;
  output s, co_BAR;


  NAND2X0 U1 ( .IN1(ci), .IN2(a), .QN(co_BAR) );
  OA21X1 U2 ( .IN1(ci), .IN2(a), .IN3(co_BAR), .Q(s) );
endmodule


module add_27 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_28 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_29 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_30 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_31 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_32 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(b), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(b), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module adder8_4 ( out, a, b, cin );
  output [7:0] out;
  input [7:0] a;
  input [7:0] b;
  input cin;

  wire   [6:0] c;

  add_32 add_01 ( .s(out[0]), .a(a[0]), .b(b[0]), .ci(1'b0), .co(c[0]) );
  add_31 add_02 ( .s(out[1]), .a(a[1]), .b(1'b0), .ci(c[0]), .co(c[1]) );
  add_30 add_03 ( .s(out[2]), .a(a[2]), .b(1'b0), .ci(c[1]), .co(c[2]) );
  add_29 add_04 ( .s(out[3]), .a(a[3]), .b(1'b0), .ci(c[2]), .co(c[3]) );
  add_28 add_05 ( .s(out[4]), .a(a[4]), .b(1'b0), .ci(c[3]), .co(c[4]) );
  add_27 add_06 ( .s(out[5]), .a(a[5]), .b(1'b0), .ci(c[4]), .co(c[5]) );
  add_26 add_07 ( .s(out[6]), .a(a[6]), .b(1'b0), .ci(c[5]), .co_BAR(c[6]) );
  add_25 add_08 ( .s(out[7]), .a(a[7]), .b(1'b0), .ci_BAR(c[6]) );
endmodule


module add_81 ( s, a, ci, co, b_BAR );
  input a, ci, b_BAR;
  output s, co;


  XNOR2X1 U1 ( .IN1(ci), .IN2(a), .Q(s) );
endmodule


module add_82 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_83 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_84 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_85 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_86 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_87 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_88 ( s, a, ci, co, b_BAR );
  input a, ci, b_BAR;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(b_BAR), .IN2(n1), .QN(co) );
  INVX0 U2 ( .INP(a), .ZN(n1) );
  MUX21X1 U3 ( .IN1(a), .IN2(n1), .S(b_BAR), .Q(s) );
endmodule


module adder8_5 ( out, a, b, cin );
  output [7:0] out;
  input [7:0] a;
  input [7:0] b;
  input cin;
  wire   n_1_net_, n_2_net_, n_3_net_;
  wire   [6:0] c;

  add_88 add_01 ( .s(out[0]), .a(a[0]), .ci(1'b1), .co(c[0]), .b_BAR(b[0]) );
  add_87 add_02 ( .s(out[1]), .a(a[1]), .b(n_1_net_), .ci(c[0]), .co(c[1]) );
  add_86 add_03 ( .s(out[2]), .a(a[2]), .b(n_2_net_), .ci(c[1]), .co(c[2]) );
  add_85 add_04 ( .s(out[3]), .a(a[3]), .b(n_3_net_), .ci(c[2]), .co(c[3]) );
  add_84 add_05 ( .s(out[4]), .a(a[4]), .b(n_3_net_), .ci(c[3]), .co(c[4]) );
  add_83 add_06 ( .s(out[5]), .a(a[5]), .b(n_3_net_), .ci(c[4]), .co(c[5]) );
  add_82 add_07 ( .s(out[6]), .a(a[6]), .b(n_3_net_), .ci(c[5]), .co(c[6]) );
  add_81 add_08 ( .s(out[7]), .a(a[7]), .ci(c[6]), .b_BAR(1'b0) );
  INVX0 U1 ( .INP(b[3]), .ZN(n_3_net_) );
  INVX0 U2 ( .INP(b[1]), .ZN(n_1_net_) );
  INVX0 U3 ( .INP(b[2]), .ZN(n_2_net_) );
endmodule


module add_89 ( s, a, ci, co, b_BAR );
  input a, ci, b_BAR;
  output s, co;


  XNOR2X1 U1 ( .IN1(b_BAR), .IN2(ci), .Q(s) );
endmodule


module add_90 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_91 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_92 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_93 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_94 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_95 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_96 ( s, a, ci, co, b_BAR );
  input a, ci, b_BAR;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(b_BAR), .IN2(n1), .QN(co) );
  INVX0 U2 ( .INP(a), .ZN(n1) );
  MUX21X1 U3 ( .IN1(a), .IN2(n1), .S(b_BAR), .Q(s) );
endmodule


module adder8_6 ( out, a, b, cin );
  output [7:0] out;
  input [7:0] a;
  input [7:0] b;
  input cin;
  wire   n_1_net_, n_2_net_, n_3_net_, n_4_net_, n_5_net_, n_6_net_;
  wire   [6:0] c;

  add_96 add_01 ( .s(out[0]), .a(a[0]), .ci(1'b1), .co(c[0]), .b_BAR(b[0]) );
  add_95 add_02 ( .s(out[1]), .a(a[1]), .b(n_1_net_), .ci(c[0]), .co(c[1]) );
  add_94 add_03 ( .s(out[2]), .a(a[2]), .b(n_2_net_), .ci(c[1]), .co(c[2]) );
  add_93 add_04 ( .s(out[3]), .a(a[3]), .b(n_3_net_), .ci(c[2]), .co(c[3]) );
  add_92 add_05 ( .s(out[4]), .a(a[4]), .b(n_4_net_), .ci(c[3]), .co(c[4]) );
  add_91 add_06 ( .s(out[5]), .a(a[5]), .b(n_5_net_), .ci(c[4]), .co(c[5]) );
  add_90 add_07 ( .s(out[6]), .a(a[6]), .b(n_6_net_), .ci(c[5]), .co(c[6]) );
  add_89 add_08 ( .s(out[7]), .a(1'b0), .ci(c[6]), .b_BAR(b[7]) );
  INVX0 U1 ( .INP(b[1]), .ZN(n_1_net_) );
  INVX0 U2 ( .INP(b[2]), .ZN(n_2_net_) );
  INVX0 U3 ( .INP(b[3]), .ZN(n_3_net_) );
  INVX0 U4 ( .INP(b[4]), .ZN(n_4_net_) );
  INVX0 U5 ( .INP(b[5]), .ZN(n_5_net_) );
  INVX0 U6 ( .INP(b[6]), .ZN(n_6_net_) );
endmodule


module floating_point_adder_1 ( clk, rst_n, input_factor_01, input_factor_02, 
        output_adder );
  input [31:0] input_factor_01;
  input [31:0] input_factor_02;
  output [31:0] output_adder;
  input clk, rst_n;
  wire   N34, N35, N36, N37, N38, N39, N40, N41, N152, N153, N154, N155, N156,
         N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, N167,
         N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178,
         N179, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189,
         N190, N191, N192, N193, N194, N195, N196, N197, N198,
         add_sub_result_24_, N211, shift_temp_01_0_, N226, N227, N228, N229,
         N230, N231, N232, N233, N234, N235, N236, N237, N238, N239, N240,
         N241, N242, N243, N244, N245, N246, N247, N248, N256, N257, N258,
         N260, N261, N262, N263, N264, N265, N266, N267, N268, N269, N270,
         N271, N272, N273, N274, N275, N276, N277, N278, N279, N280, N281,
         N306, N307, N308, N346, N347, N348, N349, N350, N351, N352, N353,
         N354, N355, N380, N381, N382, N383, N384, N385, N386, N387, N388,
         N389, N390, N391, N392, N393, N394, N395, N396, N397, N398, N399,
         N400, N401, N402, N403, N404, N405, N406, N407, N408, N409, N410, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862;
  wire   [7:0] exp_diff_value;
  wire   [7:0] exponent_factor_21;
  wire   [7:0] exponent_factor_12;
  wire   [23:0] shift_smaller_factor;
  wire   [22:0] larger_factor;
  wire   [7:0] larger_exponent;
  wire   [24:0] add_result;
  wire   [24:0] sub_result;
  wire   [22:0] pre_sig_res_01;
  wire   [3:0] shift_temp_02;
  wire   [22:1] pre_sig_res_02;
  wire   [2:0] shift_temp_03;
  wire   [22:9] pre_sig_res_03;
  wire   [4:0] shift_temp_04;
  wire   [22:16] pre_sig_res_04;
  wire   [7:0] add_output_exponent_w1;
  wire   [7:0] add_output_exponent_w2;
  wire   [7:0] add_output_exponent_w3;
  wire   [7:0] add_output_exponent_w4;

  adder8_6 adder8_01 ( .out(exponent_factor_21), .a({1'b0, 
        input_factor_02[29:23]}), .b(input_factor_01[30:23]), .cin(1'b1) );
  adder8_5 adder8_02 ( .out(exponent_factor_12), .a(input_factor_01[30:23]), 
        .b({1'b0, 1'b0, 1'b0, 1'b0, input_factor_02[26:23]}), .cin(1'b1) );
  adder24_2 adder24_01 ( .clk(clk), .rst_n(rst_n), .a({shift_temp_04[4], 
        larger_factor}), .b(shift_smaller_factor), .cin(1'b1), .out(sub_result) );
  adder24_1 adder24_02 ( .clk(clk), .rst_n(rst_n), .a({shift_temp_04[4], 
        larger_factor}), .b(shift_smaller_factor), .cin(1'b0), .out(add_result) );
  adder8_4 adder8_03 ( .out(add_output_exponent_w1), .a(larger_exponent), .b({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, shift_temp_01_0_}), .cin(
        1'b0) );
  adder8_3 adder8_04 ( .out(add_output_exponent_w2), .a(larger_exponent), .b({
        1'b0, 1'b0, 1'b0, 1'b0, shift_temp_02}), .cin(1'b1) );
  adder8_2 adder8_05 ( .out(add_output_exponent_w3), .a(larger_exponent), .b({
        1'b0, 1'b0, 1'b0, 1'b0, shift_temp_04[4], shift_temp_03}), .cin(1'b1)
         );
  adder8_1 adder8_06 ( .out(add_output_exponent_w4), .a(larger_exponent), .b({
        1'b0, 1'b0, 1'b0, shift_temp_04[4], 1'b0, shift_temp_04[2:0]}), .cin(
        1'b1) );
  DFFARX1 exp_diff_value_reg_7_ ( .D(N41), .CLK(clk), .RSTB(rst_n), .Q(
        exp_diff_value[7]) );
  DFFARX1 exp_diff_value_reg_6_ ( .D(N40), .CLK(clk), .RSTB(rst_n), .Q(
        exp_diff_value[6]) );
  DFFARX1 exp_diff_value_reg_5_ ( .D(N39), .CLK(clk), .RSTB(rst_n), .Q(
        exp_diff_value[5]) );
  DFFARX1 exp_diff_value_reg_4_ ( .D(N38), .CLK(clk), .RSTB(rst_n), .Q(
        exp_diff_value[4]) );
  DFFARX1 exp_diff_value_reg_3_ ( .D(N37), .CLK(clk), .RSTB(rst_n), .Q(
        exp_diff_value[3]), .QN(n6) );
  DFFARX1 exp_diff_value_reg_2_ ( .D(N36), .CLK(clk), .RSTB(rst_n), .Q(
        exp_diff_value[2]), .QN(n5) );
  DFFARX1 exp_diff_value_reg_1_ ( .D(N35), .CLK(clk), .RSTB(rst_n), .Q(
        exp_diff_value[1]), .QN(n7) );
  DFFARX1 exp_diff_value_reg_0_ ( .D(N34), .CLK(clk), .RSTB(rst_n), .Q(
        exp_diff_value[0]), .QN(n4) );
  DFFARX1 larger_factor_reg_22_ ( .D(N198), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[22]) );
  DFFARX1 larger_factor_reg_21_ ( .D(N197), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[21]) );
  DFFARX1 larger_factor_reg_20_ ( .D(N196), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[20]) );
  DFFARX1 larger_factor_reg_19_ ( .D(N195), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[19]) );
  DFFARX1 larger_factor_reg_18_ ( .D(N194), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[18]) );
  DFFARX1 larger_factor_reg_17_ ( .D(N193), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[17]) );
  DFFARX1 larger_factor_reg_16_ ( .D(N192), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[16]) );
  DFFARX1 larger_factor_reg_15_ ( .D(N191), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[15]) );
  DFFARX1 larger_factor_reg_14_ ( .D(N190), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[14]) );
  DFFARX1 larger_factor_reg_13_ ( .D(N189), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[13]) );
  DFFARX1 larger_factor_reg_12_ ( .D(N188), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[12]) );
  DFFARX1 larger_factor_reg_11_ ( .D(N187), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[11]) );
  DFFARX1 larger_factor_reg_10_ ( .D(N186), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[10]) );
  DFFARX1 larger_factor_reg_9_ ( .D(N185), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[9]) );
  DFFARX1 larger_factor_reg_8_ ( .D(N184), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[8]) );
  DFFARX1 larger_factor_reg_7_ ( .D(N183), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[7]) );
  DFFARX1 larger_factor_reg_6_ ( .D(N182), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[6]) );
  DFFARX1 larger_factor_reg_5_ ( .D(N181), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[5]) );
  DFFARX1 larger_factor_reg_4_ ( .D(N180), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[4]) );
  DFFARX1 larger_factor_reg_3_ ( .D(N179), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[3]) );
  DFFARX1 larger_factor_reg_2_ ( .D(N178), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[2]) );
  DFFARX1 larger_factor_reg_1_ ( .D(N177), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[1]) );
  DFFARX1 larger_factor_reg_0_ ( .D(N176), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[0]) );
  DFFARX1 shift_smaller_factor_reg_23_ ( .D(N175), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[23]) );
  DFFARX1 shift_smaller_factor_reg_22_ ( .D(N174), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[22]) );
  DFFARX1 shift_smaller_factor_reg_21_ ( .D(N173), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[21]) );
  DFFARX1 shift_smaller_factor_reg_20_ ( .D(N172), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[20]) );
  DFFARX1 shift_smaller_factor_reg_19_ ( .D(N171), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[19]) );
  DFFARX1 shift_smaller_factor_reg_18_ ( .D(N170), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[18]) );
  DFFARX1 shift_smaller_factor_reg_17_ ( .D(N169), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[17]) );
  DFFARX1 shift_smaller_factor_reg_16_ ( .D(N168), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[16]) );
  DFFARX1 shift_smaller_factor_reg_15_ ( .D(N167), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[15]) );
  DFFARX1 shift_smaller_factor_reg_14_ ( .D(N166), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[14]) );
  DFFARX1 shift_smaller_factor_reg_13_ ( .D(N165), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[13]) );
  DFFARX1 shift_smaller_factor_reg_12_ ( .D(N164), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[12]) );
  DFFARX1 shift_smaller_factor_reg_11_ ( .D(N163), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[11]) );
  DFFARX1 shift_smaller_factor_reg_10_ ( .D(N162), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[10]) );
  DFFARX1 shift_smaller_factor_reg_9_ ( .D(N161), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[9]) );
  DFFARX1 shift_smaller_factor_reg_8_ ( .D(N160), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[8]) );
  DFFARX1 shift_smaller_factor_reg_7_ ( .D(N159), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[7]) );
  DFFARX1 shift_smaller_factor_reg_6_ ( .D(N158), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[6]) );
  DFFARX1 shift_smaller_factor_reg_5_ ( .D(N157), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[5]) );
  DFFARX1 shift_smaller_factor_reg_4_ ( .D(N156), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[4]) );
  DFFARX1 shift_smaller_factor_reg_3_ ( .D(N155), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[3]) );
  DFFARX1 shift_smaller_factor_reg_2_ ( .D(N154), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[2]) );
  DFFARX1 shift_smaller_factor_reg_1_ ( .D(N153), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[1]) );
  DFFARX1 shift_smaller_factor_reg_0_ ( .D(N152), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[0]) );
  DFFX1 larger_exponent_reg_7_ ( .D(n840), .CLK(clk), .Q(larger_exponent[7])
         );
  DFFX1 larger_exponent_reg_6_ ( .D(n841), .CLK(clk), .Q(larger_exponent[6])
         );
  DFFX1 larger_exponent_reg_5_ ( .D(n842), .CLK(clk), .Q(larger_exponent[5])
         );
  DFFX1 larger_exponent_reg_4_ ( .D(n843), .CLK(clk), .Q(larger_exponent[4])
         );
  DFFX1 larger_exponent_reg_3_ ( .D(n844), .CLK(clk), .Q(larger_exponent[3])
         );
  DFFX1 larger_exponent_reg_2_ ( .D(n845), .CLK(clk), .Q(larger_exponent[2])
         );
  DFFX1 larger_exponent_reg_1_ ( .D(n846), .CLK(clk), .Q(larger_exponent[1])
         );
  DFFX1 larger_exponent_reg_0_ ( .D(n847), .CLK(clk), .Q(larger_exponent[0])
         );
  DFFARX1 shift_temp_04_reg_4_ ( .D(1'b1), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_04[4]) );
  DFFARX1 shift_temp_01_reg_0_ ( .D(add_sub_result_24_), .CLK(clk), .RSTB(
        rst_n), .Q(shift_temp_01_0_) );
  DFFARX1 pre_sig_res_02_reg_1_ ( .D(N260), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[1]) );
  DFFARX1 pre_sig_res_02_reg_2_ ( .D(N261), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[2]) );
  DFFARX1 pre_sig_res_02_reg_3_ ( .D(N262), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[3]) );
  DFFARX1 pre_sig_res_02_reg_4_ ( .D(N263), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[4]) );
  DFFARX1 pre_sig_res_02_reg_5_ ( .D(N264), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[5]) );
  DFFARX1 pre_sig_res_02_reg_6_ ( .D(N265), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[6]) );
  DFFARX1 pre_sig_res_02_reg_7_ ( .D(N266), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[7]) );
  DFFARX1 shift_temp_02_reg_2_ ( .D(N258), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_02[2]) );
  DFFASX1 shift_temp_02_reg_3_ ( .D(n839), .CLK(clk), .SETB(rst_n), .QN(
        shift_temp_02[3]) );
  DFFARX1 pre_sig_res_02_reg_8_ ( .D(N267), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[8]) );
  DFFARX1 pre_sig_res_02_reg_9_ ( .D(N268), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[9]) );
  DFFARX1 pre_sig_res_02_reg_10_ ( .D(N269), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[10]) );
  DFFARX1 pre_sig_res_02_reg_11_ ( .D(N270), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[11]) );
  DFFARX1 pre_sig_res_02_reg_12_ ( .D(N271), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[12]) );
  DFFARX1 pre_sig_res_02_reg_13_ ( .D(N272), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[13]) );
  DFFARX1 pre_sig_res_02_reg_14_ ( .D(N273), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[14]) );
  DFFARX1 pre_sig_res_02_reg_15_ ( .D(N274), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[15]) );
  DFFARX1 pre_sig_res_02_reg_16_ ( .D(N275), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[16]) );
  DFFARX1 pre_sig_res_02_reg_17_ ( .D(N276), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[17]) );
  DFFARX1 pre_sig_res_02_reg_18_ ( .D(N277), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[18]) );
  DFFARX1 pre_sig_res_02_reg_19_ ( .D(N278), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[19]) );
  DFFARX1 pre_sig_res_02_reg_20_ ( .D(N279), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[20]) );
  DFFARX1 pre_sig_res_02_reg_21_ ( .D(N280), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[21]) );
  DFFARX1 pre_sig_res_02_reg_22_ ( .D(N281), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[22]) );
  DFFARX1 shift_temp_02_reg_1_ ( .D(N257), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_02[1]) );
  DFFARX1 shift_temp_02_reg_0_ ( .D(N256), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_02[0]) );
  DFFX1 pre_sig_res_03_reg_9_ ( .D(n848), .CLK(clk), .Q(pre_sig_res_03[9]) );
  DFFX1 pre_sig_res_03_reg_10_ ( .D(n849), .CLK(clk), .Q(pre_sig_res_03[10])
         );
  DFFX1 pre_sig_res_03_reg_12_ ( .D(n850), .CLK(clk), .Q(pre_sig_res_03[12])
         );
  DFFX1 pre_sig_res_03_reg_11_ ( .D(n851), .CLK(clk), .Q(pre_sig_res_03[11])
         );
  DFFX1 pre_sig_res_03_reg_13_ ( .D(n852), .CLK(clk), .Q(pre_sig_res_03[13])
         );
  DFFX1 pre_sig_res_03_reg_14_ ( .D(n853), .CLK(clk), .Q(pre_sig_res_03[14])
         );
  DFFARX1 shift_temp_03_reg_2_ ( .D(N308), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_03[2]) );
  DFFARX1 shift_temp_03_reg_0_ ( .D(N306), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_03[0]) );
  DFFARX1 shift_temp_03_reg_1_ ( .D(N307), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_03[1]) );
  DFFX1 pre_sig_res_03_reg_15_ ( .D(n854), .CLK(clk), .Q(pre_sig_res_03[15])
         );
  DFFX1 pre_sig_res_03_reg_16_ ( .D(n855), .CLK(clk), .Q(pre_sig_res_03[16])
         );
  DFFX1 pre_sig_res_03_reg_17_ ( .D(n856), .CLK(clk), .Q(pre_sig_res_03[17])
         );
  DFFX1 pre_sig_res_03_reg_18_ ( .D(n857), .CLK(clk), .Q(pre_sig_res_03[18])
         );
  DFFX1 pre_sig_res_03_reg_19_ ( .D(n858), .CLK(clk), .Q(pre_sig_res_03[19])
         );
  DFFX1 pre_sig_res_03_reg_20_ ( .D(n859), .CLK(clk), .Q(pre_sig_res_03[20])
         );
  DFFX1 pre_sig_res_03_reg_21_ ( .D(n860), .CLK(clk), .Q(pre_sig_res_03[21])
         );
  DFFX1 pre_sig_res_03_reg_22_ ( .D(n861), .CLK(clk), .Q(pre_sig_res_03[22])
         );
  DFFARX1 pre_sig_res_04_reg_16_ ( .D(N349), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_04[16]) );
  DFFARX1 pre_sig_res_04_reg_17_ ( .D(N350), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_04[17]) );
  DFFARX1 pre_sig_res_04_reg_18_ ( .D(N351), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_04[18]) );
  DFFARX1 pre_sig_res_04_reg_19_ ( .D(N352), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_04[19]) );
  DFFARX1 pre_sig_res_04_reg_20_ ( .D(N353), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_04[20]) );
  DFFARX1 pre_sig_res_04_reg_21_ ( .D(N354), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_04[21]) );
  DFFARX1 pre_sig_res_04_reg_22_ ( .D(N355), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_04[22]) );
  DFFARX1 add_output_sign_reg ( .D(N211), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[31]) );
  DFFARX1 pre_sig_res_01_reg_0_ ( .D(N226), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[0]) );
  DFFARX1 pre_sig_res_01_reg_1_ ( .D(N227), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[1]) );
  DFFARX1 pre_sig_res_01_reg_2_ ( .D(N228), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[2]) );
  DFFARX1 pre_sig_res_01_reg_3_ ( .D(N229), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[3]) );
  DFFARX1 pre_sig_res_01_reg_4_ ( .D(N230), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[4]) );
  DFFARX1 pre_sig_res_01_reg_5_ ( .D(N231), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[5]) );
  DFFARX1 pre_sig_res_01_reg_6_ ( .D(N232), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[6]) );
  DFFARX1 pre_sig_res_01_reg_7_ ( .D(N233), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[7]) );
  DFFARX1 pre_sig_res_01_reg_8_ ( .D(N234), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[8]) );
  DFFARX1 pre_sig_res_01_reg_9_ ( .D(N235), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[9]) );
  DFFARX1 pre_sig_res_01_reg_10_ ( .D(N236), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[10]) );
  DFFARX1 pre_sig_res_01_reg_11_ ( .D(N237), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[11]) );
  DFFARX1 pre_sig_res_01_reg_12_ ( .D(N238), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[12]) );
  DFFARX1 pre_sig_res_01_reg_13_ ( .D(N239), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[13]) );
  DFFARX1 pre_sig_res_01_reg_14_ ( .D(N240), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[14]) );
  DFFARX1 pre_sig_res_01_reg_15_ ( .D(N241), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[15]) );
  DFFARX1 pre_sig_res_01_reg_16_ ( .D(N242), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[16]) );
  DFFARX1 pre_sig_res_01_reg_17_ ( .D(N243), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[17]) );
  DFFARX1 pre_sig_res_01_reg_18_ ( .D(N244), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[18]) );
  DFFARX1 pre_sig_res_01_reg_19_ ( .D(N245), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[19]) );
  DFFARX1 pre_sig_res_01_reg_20_ ( .D(N246), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[20]) );
  DFFARX1 pre_sig_res_01_reg_21_ ( .D(N247), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[21]) );
  DFFARX1 pre_sig_res_01_reg_22_ ( .D(N248), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[22]) );
  DFFARX1 shift_temp_04_reg_2_ ( .D(N348), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_04[2]) );
  DFFARX1 shift_temp_04_reg_1_ ( .D(N347), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_04[1]) );
  DFFARX1 shift_temp_04_reg_0_ ( .D(N346), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_04[0]) );
  DFFARX1 add_output_exponent_reg_7_ ( .D(N387), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[30]) );
  DFFARX1 add_output_exponent_reg_6_ ( .D(N386), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[29]) );
  DFFARX1 add_output_exponent_reg_5_ ( .D(N385), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[28]) );
  DFFARX1 add_output_exponent_reg_4_ ( .D(N384), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[27]) );
  DFFARX1 add_output_exponent_reg_3_ ( .D(N383), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[26]) );
  DFFARX1 add_output_exponent_reg_2_ ( .D(N382), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[25]) );
  DFFARX1 add_output_exponent_reg_1_ ( .D(N381), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[24]) );
  DFFARX1 add_output_exponent_reg_0_ ( .D(N380), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[23]) );
  DFFARX1 add_output_significands_reg_22_ ( .D(N410), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[22]) );
  DFFARX1 add_output_significands_reg_21_ ( .D(N409), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[21]) );
  DFFARX1 add_output_significands_reg_20_ ( .D(N408), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[20]) );
  DFFARX1 add_output_significands_reg_19_ ( .D(N407), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[19]) );
  DFFARX1 add_output_significands_reg_18_ ( .D(N406), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[18]) );
  DFFARX1 add_output_significands_reg_17_ ( .D(N405), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[17]) );
  DFFARX1 add_output_significands_reg_16_ ( .D(N404), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[16]) );
  DFFARX1 add_output_significands_reg_15_ ( .D(N403), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[15]) );
  DFFARX1 add_output_significands_reg_14_ ( .D(N402), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[14]) );
  DFFARX1 add_output_significands_reg_13_ ( .D(N401), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[13]) );
  DFFARX1 add_output_significands_reg_12_ ( .D(N400), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[12]) );
  DFFARX1 add_output_significands_reg_11_ ( .D(N399), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[11]) );
  DFFARX1 add_output_significands_reg_10_ ( .D(N398), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[10]) );
  DFFARX1 add_output_significands_reg_9_ ( .D(N397), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[9]) );
  DFFARX1 add_output_significands_reg_8_ ( .D(N396), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[8]) );
  DFFARX1 add_output_significands_reg_7_ ( .D(N395), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[7]) );
  DFFARX1 add_output_significands_reg_6_ ( .D(N394), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[6]) );
  DFFARX1 add_output_significands_reg_5_ ( .D(N393), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[5]) );
  DFFARX1 add_output_significands_reg_4_ ( .D(N392), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[4]) );
  DFFARX1 add_output_significands_reg_3_ ( .D(N391), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[3]) );
  DFFARX1 add_output_significands_reg_2_ ( .D(N390), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[2]) );
  DFFARX1 add_output_significands_reg_1_ ( .D(N389), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[1]) );
  DFFARX1 add_output_significands_reg_0_ ( .D(N388), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[0]) );
  INVX1 U5 ( .INP(rst_n), .ZN(n862) );
  NAND2X0 U3 ( .IN1(input_factor_01[0]), .IN2(n76), .QN(n42) );
  NAND2X0 U4 ( .IN1(n492), .IN2(n405), .QN(n564) );
  NAND2X0 U6 ( .IN1(n38), .IN2(n20), .QN(n22) );
  NAND2X0 U7 ( .IN1(input_factor_01[24]), .IN2(n32), .QN(n19) );
  NAND2X0 U8 ( .IN1(input_factor_01[23]), .IN2(n390), .QN(n18) );
  NAND2X0 U9 ( .IN1(n811), .IN2(n532), .QN(n388) );
  NAND2X0 U10 ( .IN1(n781), .IN2(n524), .QN(n387) );
  NAND2X0 U11 ( .IN1(n774), .IN2(n525), .QN(n386) );
  NAND2X0 U12 ( .IN1(n750), .IN2(n724), .QN(n567) );
  NAND2X0 U13 ( .IN1(n409), .IN2(n502), .QN(n384) );
  NAND2X0 U14 ( .IN1(n500), .IN2(n412), .QN(n383) );
  NAND2X0 U15 ( .IN1(n382), .IN2(n570), .QN(n411) );
  NAND2X0 U16 ( .IN1(n69), .IN2(n68), .QN(n222) );
  NAND2X0 U17 ( .IN1(n81), .IN2(n80), .QN(n221) );
  NAND2X0 U18 ( .IN1(n124), .IN2(n123), .QN(n238) );
  NAND2X0 U19 ( .IN1(n134), .IN2(n133), .QN(n237) );
  NAND2X0 U20 ( .IN1(n154), .IN2(n153), .QN(n254) );
  NAND2X0 U21 ( .IN1(n164), .IN2(n163), .QN(n253) );
  NAND2X0 U22 ( .IN1(n825), .IN2(n275), .QN(n255) );
  NAND2X0 U23 ( .IN1(n275), .IN2(n709), .QN(n256) );
  NAND2X0 U24 ( .IN1(n188), .IN2(n187), .QN(n274) );
  NAND2X0 U25 ( .IN1(n198), .IN2(n197), .QN(n273) );
  NAND2X0 U26 ( .IN1(n73), .IN2(n72), .QN(n215) );
  NAND2X0 U27 ( .IN1(n85), .IN2(n84), .QN(n218) );
  NAND2X0 U28 ( .IN1(n128), .IN2(n127), .QN(n231) );
  NAND2X0 U29 ( .IN1(n139), .IN2(n137), .QN(n234) );
  NAND2X0 U30 ( .IN1(n158), .IN2(n157), .QN(n247) );
  NAND2X0 U31 ( .IN1(n168), .IN2(n167), .QN(n250) );
  NAND2X0 U32 ( .IN1(n192), .IN2(n191), .QN(n267) );
  NAND2X0 U33 ( .IN1(n205), .IN2(n204), .QN(n270) );
  NAND2X0 U34 ( .IN1(n28), .IN2(n29), .QN(n12) );
  NAND2X0 U35 ( .IN1(input_factor_01[16]), .IN2(n332), .QN(n28) );
  NAND2X0 U36 ( .IN1(input_factor_01[25]), .IN2(n390), .QN(n38) );
  NAND2X0 U37 ( .IN1(n379), .IN2(n377), .QN(n827) );
  NAND2X0 U38 ( .IN1(n716), .IN2(pre_sig_res_01[9]), .QN(n635) );
  NAND2X0 U39 ( .IN1(n716), .IN2(pre_sig_res_01[10]), .QN(n641) );
  NAND2X0 U40 ( .IN1(n716), .IN2(pre_sig_res_01[11]), .QN(n647) );
  NAND2X0 U41 ( .IN1(n716), .IN2(pre_sig_res_01[12]), .QN(n653) );
  NAND2X0 U42 ( .IN1(n716), .IN2(pre_sig_res_01[13]), .QN(n659) );
  NAND2X0 U43 ( .IN1(n716), .IN2(pre_sig_res_01[14]), .QN(n665) );
  NAND2X0 U44 ( .IN1(n716), .IN2(pre_sig_res_01[15]), .QN(n671) );
  NAND2X0 U45 ( .IN1(n716), .IN2(pre_sig_res_01[16]), .QN(n675) );
  NAND2X0 U46 ( .IN1(n716), .IN2(pre_sig_res_01[17]), .QN(n681) );
  NAND2X0 U47 ( .IN1(n716), .IN2(pre_sig_res_01[18]), .QN(n687) );
  NAND2X0 U48 ( .IN1(n716), .IN2(pre_sig_res_01[19]), .QN(n693) );
  NAND2X0 U49 ( .IN1(n716), .IN2(pre_sig_res_01[20]), .QN(n699) );
  NAND2X0 U50 ( .IN1(n716), .IN2(pre_sig_res_01[21]), .QN(n705) );
  NAND2X0 U51 ( .IN1(n716), .IN2(pre_sig_res_01[22]), .QN(n717) );
  NAND2X0 U52 ( .IN1(n716), .IN2(add_output_exponent_w1[1]), .QN(n576) );
  NAND2X0 U53 ( .IN1(n526), .IN2(n821), .QN(n544) );
  NAND2X0 U54 ( .IN1(n523), .IN2(n532), .QN(n529) );
  NAND2X0 U55 ( .IN1(n524), .IN2(n794), .QN(n542) );
  NAND2X0 U56 ( .IN1(n525), .IN2(n761), .QN(n543) );
  NAND2X0 U57 ( .IN1(n766), .IN2(n750), .QN(n725) );
  NAND2X0 U58 ( .IN1(n724), .IN2(n737), .QN(n799) );
  NAND2X0 U59 ( .IN1(n522), .IN2(n510), .QN(n728) );
  NAND2X0 U60 ( .IN1(n522), .IN2(n514), .QN(n721) );
  NAND2X0 U61 ( .IN1(n405), .IN2(n404), .QN(n504) );
  NAND2X0 U62 ( .IN1(n422), .IN2(n823), .QN(n419) );
  NAND2X0 U63 ( .IN1(n409), .IN2(n406), .QN(n493) );
  NAND2X0 U64 ( .IN1(n412), .IN2(n407), .QN(n497) );
  NAND2X0 U65 ( .IN1(n408), .IN2(n570), .QN(n495) );
  NAND2X0 U66 ( .IN1(n67), .IN2(n66), .QN(n74) );
  NAND2X0 U67 ( .IN1(n79), .IN2(n77), .QN(n86) );
  NAND2X0 U68 ( .IN1(input_factor_01[0]), .IN2(n184), .QN(n90) );
  NAND2X0 U69 ( .IN1(n122), .IN2(n121), .QN(n129) );
  NAND2X0 U70 ( .IN1(n132), .IN2(n131), .QN(n140) );
  NAND2X0 U71 ( .IN1(input_factor_01[1]), .IN2(n184), .QN(n144) );
  NAND2X0 U72 ( .IN1(n152), .IN2(n151), .QN(n159) );
  NAND2X0 U73 ( .IN1(n162), .IN2(n161), .QN(n169) );
  NAND2X0 U74 ( .IN1(input_factor_01[2]), .IN2(n184), .QN(n173) );
  NAND2X0 U75 ( .IN1(n275), .IN2(n6), .QN(n182) );
  NAND2X0 U76 ( .IN1(n186), .IN2(n185), .QN(n193) );
  NAND2X0 U77 ( .IN1(n196), .IN2(n195), .QN(n206) );
  NAND2X0 U78 ( .IN1(input_factor_01[3]), .IN2(n184), .QN(n210) );
  NAND2X0 U79 ( .IN1(n83), .IN2(n82), .QN(n214) );
  NAND2X0 U80 ( .IN1(n71), .IN2(n70), .QN(n213) );
  NAND2X0 U81 ( .IN1(n136), .IN2(n135), .QN(n230) );
  NAND2X0 U82 ( .IN1(n126), .IN2(n125), .QN(n229) );
  NAND2X0 U83 ( .IN1(n166), .IN2(n165), .QN(n246) );
  NAND2X0 U84 ( .IN1(n156), .IN2(n155), .QN(n245) );
  NAND2X0 U85 ( .IN1(n379), .IN2(n366), .QN(n276) );
  NAND2X0 U86 ( .IN1(n200), .IN2(n199), .QN(n265) );
  NAND2X0 U87 ( .IN1(n190), .IN2(n189), .QN(n263) );
  NAND2X0 U88 ( .IN1(exp_diff_value[3]), .IN2(n357), .QN(n330) );
  NAND2X0 U89 ( .IN1(exp_diff_value[3]), .IN2(n355), .QN(n331) );
  NAND2X0 U90 ( .IN1(n331), .IN2(n330), .QN(n333) );
  NAND2X0 U91 ( .IN1(n357), .IN2(n6), .QN(n351) );
  NAND2X0 U92 ( .IN1(n355), .IN2(n6), .QN(n349) );
  NAND2X0 U93 ( .IN1(n366), .IN2(n65), .QN(n378) );
  NAND2X0 U94 ( .IN1(n357), .IN2(n356), .QN(n367) );
  NAND2X0 U95 ( .IN1(n356), .IN2(n355), .QN(n369) );
  NAND2X0 U96 ( .IN1(input_factor_01[27]), .IN2(n389), .QN(n37) );
  NAND2X0 U97 ( .IN1(n380), .IN2(n379), .QN(n399) );
  NAND2X0 U98 ( .IN1(n827), .IN2(n378), .QN(n401) );
  NAND2X0 U99 ( .IN1(n602), .IN2(n601), .QN(N389) );
  NAND2X0 U100 ( .IN1(n606), .IN2(n605), .QN(N390) );
  NAND2X0 U101 ( .IN1(n610), .IN2(n609), .QN(N391) );
  NAND2X0 U102 ( .IN1(n614), .IN2(n613), .QN(N392) );
  NAND2X0 U103 ( .IN1(n618), .IN2(n617), .QN(N393) );
  NAND2X0 U104 ( .IN1(n622), .IN2(n621), .QN(N394) );
  NAND2X0 U105 ( .IN1(n626), .IN2(n625), .QN(N395) );
  NAND2X0 U106 ( .IN1(n630), .IN2(n629), .QN(N396) );
  NAND2X0 U107 ( .IN1(n714), .IN2(pre_sig_res_03[9]), .QN(n633) );
  NAND2X0 U108 ( .IN1(n713), .IN2(pre_sig_res_02[9]), .QN(n634) );
  NAND2X0 U109 ( .IN1(n714), .IN2(pre_sig_res_03[10]), .QN(n639) );
  NAND2X0 U110 ( .IN1(n713), .IN2(pre_sig_res_02[10]), .QN(n640) );
  NAND2X0 U111 ( .IN1(n714), .IN2(pre_sig_res_03[11]), .QN(n645) );
  NAND2X0 U112 ( .IN1(n713), .IN2(pre_sig_res_02[11]), .QN(n646) );
  NAND2X0 U113 ( .IN1(n714), .IN2(pre_sig_res_03[12]), .QN(n651) );
  NAND2X0 U114 ( .IN1(n713), .IN2(pre_sig_res_02[12]), .QN(n652) );
  NAND2X0 U115 ( .IN1(n714), .IN2(pre_sig_res_03[13]), .QN(n657) );
  NAND2X0 U116 ( .IN1(n713), .IN2(pre_sig_res_02[13]), .QN(n658) );
  NAND2X0 U117 ( .IN1(n714), .IN2(pre_sig_res_03[14]), .QN(n663) );
  NAND2X0 U118 ( .IN1(n713), .IN2(pre_sig_res_02[14]), .QN(n664) );
  NAND2X0 U119 ( .IN1(n714), .IN2(pre_sig_res_03[15]), .QN(n669) );
  NAND2X0 U120 ( .IN1(n713), .IN2(pre_sig_res_02[15]), .QN(n670) );
  NAND2X0 U121 ( .IN1(n715), .IN2(pre_sig_res_04[16]), .QN(n676) );
  NAND2X0 U122 ( .IN1(n715), .IN2(pre_sig_res_04[17]), .QN(n682) );
  NAND2X0 U123 ( .IN1(n715), .IN2(pre_sig_res_04[18]), .QN(n688) );
  NAND2X0 U124 ( .IN1(n715), .IN2(pre_sig_res_04[19]), .QN(n694) );
  NAND2X0 U125 ( .IN1(n715), .IN2(pre_sig_res_04[20]), .QN(n700) );
  NAND2X0 U126 ( .IN1(n715), .IN2(pre_sig_res_04[21]), .QN(n706) );
  NAND2X0 U127 ( .IN1(n715), .IN2(pre_sig_res_04[22]), .QN(n718) );
  NAND2X0 U128 ( .IN1(n714), .IN2(add_output_exponent_w3[0]), .QN(n573) );
  NAND2X0 U129 ( .IN1(n715), .IN2(add_output_exponent_w4[1]), .QN(n577) );
  NAND2X0 U130 ( .IN1(n715), .IN2(add_output_exponent_w4[2]), .QN(n580) );
  NAND2X0 U131 ( .IN1(n714), .IN2(add_output_exponent_w3[3]), .QN(n584) );
  NAND2X0 U132 ( .IN1(n714), .IN2(add_output_exponent_w3[4]), .QN(n587) );
  NAND2X0 U133 ( .IN1(n714), .IN2(add_output_exponent_w3[5]), .QN(n590) );
  NAND2X0 U134 ( .IN1(n715), .IN2(add_output_exponent_w4[6]), .QN(n593) );
  NAND2X0 U135 ( .IN1(n9), .IN2(n10), .QN(N387) );
  NAND2X0 U136 ( .IN1(n715), .IN2(add_output_exponent_w4[7]), .QN(n10) );
  NAND2X0 U137 ( .IN1(n529), .IN2(n528), .QN(N348) );
  NAND2X0 U138 ( .IN1(n546), .IN2(n801), .QN(n547) );
  NAND2X0 U139 ( .IN1(n546), .IN2(n821), .QN(n537) );
  NAND2X0 U140 ( .IN1(n546), .IN2(n823), .QN(n533) );
  NAND2X0 U141 ( .IN1(n531), .IN2(n530), .QN(N352) );
  NAND2X0 U142 ( .IN1(pre_sig_res_03[22]), .IN2(n826), .QN(n730) );
  NAND2X0 U143 ( .IN1(n814), .IN2(n729), .QN(n731) );
  NAND2X0 U144 ( .IN1(pre_sig_res_03[21]), .IN2(n826), .QN(n738) );
  NAND2X0 U145 ( .IN1(n814), .IN2(n737), .QN(n739) );
  NAND2X0 U146 ( .IN1(pre_sig_res_03[20]), .IN2(n826), .QN(n746) );
  NAND2X0 U147 ( .IN1(n814), .IN2(n745), .QN(n747) );
  NAND2X0 U148 ( .IN1(pre_sig_res_03[19]), .IN2(n826), .QN(n754) );
  NAND2X0 U149 ( .IN1(n814), .IN2(n753), .QN(n755) );
  NAND2X0 U150 ( .IN1(pre_sig_res_03[18]), .IN2(n826), .QN(n762) );
  NAND2X0 U151 ( .IN1(n814), .IN2(n761), .QN(n763) );
  NAND2X0 U152 ( .IN1(pre_sig_res_03[17]), .IN2(n826), .QN(n770) );
  NAND2X0 U153 ( .IN1(n814), .IN2(n769), .QN(n771) );
  NAND2X0 U154 ( .IN1(pre_sig_res_03[16]), .IN2(n826), .QN(n777) );
  NAND2X0 U155 ( .IN1(n814), .IN2(n794), .QN(n778) );
  NAND2X0 U156 ( .IN1(pre_sig_res_03[15]), .IN2(n826), .QN(n786) );
  NAND2X0 U157 ( .IN1(n814), .IN2(n802), .QN(n787) );
  NAND2X0 U158 ( .IN1(n721), .IN2(n728), .QN(n515) );
  NAND2X0 U159 ( .IN1(pre_sig_res_03[14]), .IN2(n862), .QN(n796) );
  NAND2X0 U160 ( .IN1(n824), .IN2(n794), .QN(n795) );
  NAND2X0 U161 ( .IN1(n814), .IN2(n793), .QN(n797) );
  NAND2X0 U162 ( .IN1(pre_sig_res_03[13]), .IN2(n826), .QN(n804) );
  NAND2X0 U163 ( .IN1(n824), .IN2(n802), .QN(n803) );
  NAND2X0 U164 ( .IN1(n814), .IN2(n801), .QN(n805) );
  NAND2X0 U165 ( .IN1(n809), .IN2(n808), .QN(n851) );
  NAND2X0 U166 ( .IN1(pre_sig_res_03[12]), .IN2(n826), .QN(n817) );
  NAND2X0 U167 ( .IN1(n814), .IN2(n821), .QN(n819) );
  NAND2X0 U168 ( .IN1(n422), .IN2(n821), .QN(n423) );
  NAND2X0 U169 ( .IN1(n427), .IN2(n802), .QN(n418) );
  NAND2X0 U170 ( .IN1(n428), .IN2(n801), .QN(n415) );
  NAND2X0 U171 ( .IN1(n414), .IN2(n413), .QN(N263) );
  NAND2X0 U172 ( .IN1(n828), .IN2(n829), .QN(n847) );
  NAND2X0 U173 ( .IN1(n830), .IN2(n829), .QN(n845) );
  NAND2X0 U174 ( .IN1(n832), .IN2(n836), .QN(n844) );
  NAND2X0 U175 ( .IN1(n833), .IN2(n836), .QN(n843) );
  NAND2X0 U176 ( .IN1(n834), .IN2(n836), .QN(n842) );
  NAND2X0 U177 ( .IN1(n837), .IN2(n836), .QN(n841) );
  NAND2X0 U178 ( .IN1(n355), .IN2(n87), .QN(n88) );
  NAND2X0 U179 ( .IN1(n357), .IN2(n75), .QN(n89) );
  NAND2X0 U180 ( .IN1(n355), .IN2(n141), .QN(n142) );
  NAND2X0 U181 ( .IN1(n357), .IN2(n130), .QN(n143) );
  NAND2X0 U182 ( .IN1(n355), .IN2(n170), .QN(n171) );
  NAND2X0 U183 ( .IN1(n357), .IN2(n160), .QN(n172) );
  NAND2X0 U184 ( .IN1(n355), .IN2(n207), .QN(n208) );
  NAND2X0 U185 ( .IN1(n357), .IN2(n194), .QN(n209) );
  NAND2X0 U186 ( .IN1(n340), .IN2(n339), .QN(N168) );
  NAND2X0 U187 ( .IN1(n344), .IN2(n343), .QN(N169) );
  NAND2X0 U188 ( .IN1(n348), .IN2(n347), .QN(N170) );
  NAND2X0 U189 ( .IN1(n354), .IN2(n353), .QN(N171) );
  NAND2X0 U190 ( .IN1(n361), .IN2(n360), .QN(N172) );
  NAND2X0 U191 ( .IN1(n365), .IN2(n364), .QN(N173) );
  NAND2X0 U192 ( .IN1(n372), .IN2(n371), .QN(N174) );
  NAND2X0 U193 ( .IN1(n377), .IN2(n376), .QN(N175) );
  NAND2X0 U197 ( .IN1(input_factor_02[29]), .IN2(n831), .QN(n836) );
  INVX0 U198 ( .INP(n563), .ZN(n839) );
  INVX0 U199 ( .INP(n427), .ZN(n499) );
  NOR2X0 U200 ( .IN1(n728), .IN2(n826), .QN(n814) );
  INVX0 U201 ( .INP(n822), .ZN(n812) );
  INVX0 U202 ( .INP(n801), .ZN(n813) );
  INVX0 U203 ( .INP(n802), .ZN(n791) );
  INVX0 U204 ( .INP(n769), .ZN(n782) );
  NAND2X0 U205 ( .IN1(input_factor_02[29]), .IN2(n16), .QN(n594) );
  NOR2X0 U206 ( .IN1(n572), .IN2(n571), .QN(n714) );
  INVX0 U207 ( .INP(n745), .ZN(n758) );
  INVX0 U208 ( .INP(n564), .ZN(n522) );
  INVX0 U209 ( .INP(n753), .ZN(n766) );
  NOR2X0 U210 ( .IN1(n568), .IN2(n571), .QN(n713) );
  INVX0 U211 ( .INP(n464), .ZN(n565) );
  NOR2X0 U212 ( .IN1(n570), .IN2(n571), .QN(n716) );
  NAND4X0 U213 ( .IN1(n561), .IN2(n560), .IN3(n559), .IN4(n558), .QN(n711) );
  INVX0 U214 ( .INP(n8), .ZN(n15) );
  INVX0 U215 ( .INP(n379), .ZN(n709) );
  INVX0 U216 ( .INP(n827), .ZN(n825) );
  INVX0 U217 ( .INP(n178), .ZN(n202) );
  INVX0 U218 ( .INP(n179), .ZN(n203) );
  INVX0 U219 ( .INP(n332), .ZN(n374) );
  INVX0 U220 ( .INP(n177), .ZN(n201) );
  OR2X1 U221 ( .IN1(n65), .IN2(n377), .Q(n380) );
  INVX0 U222 ( .INP(input_factor_01[22]), .ZN(n710) );
  NOR3X0 U223 ( .IN1(input_factor_01[30]), .IN2(n25), .IN3(n24), .QN(n379) );
  INVX0 U224 ( .INP(input_factor_02[23]), .ZN(n390) );
  INVX0 U225 ( .INP(input_factor_02[29]), .ZN(n389) );
  INVX0 U226 ( .INP(n406), .ZN(n502) );
  NOR2X0 U227 ( .IN1(add_sub_result_24_), .IN2(n403), .QN(n570) );
  MUX21X1 U228 ( .IN1(sub_result[24]), .IN2(add_result[24]), .S(n13), .Q(
        add_sub_result_24_) );
  INVX0 U229 ( .INP(n404), .ZN(n492) );
  INVX0 U230 ( .INP(n14), .ZN(n13) );
  INVX0 U231 ( .INP(n511), .ZN(n14) );
  INVX0 U232 ( .INP(n737), .ZN(n750) );
  INVX0 U233 ( .INP(n761), .ZN(n774) );
  INVX0 U234 ( .INP(n794), .ZN(n781) );
  INVX0 U235 ( .INP(n793), .ZN(n811) );
  INVX0 U236 ( .INP(n821), .ZN(n807) );
  INVX0 U237 ( .INP(n823), .ZN(n815) );
  MUX21X1 U238 ( .IN1(n381), .IN2(input_factor_01[31]), .S(input_factor_02[31]), .Q(n511) );
  INVX0 U239 ( .INP(input_factor_01[31]), .ZN(n381) );
  INVX0 U240 ( .INP(n455), .ZN(n723) );
  INVX0 U241 ( .INP(n729), .ZN(n742) );
  INVX0 U242 ( .INP(n824), .ZN(n810) );
  INVX0 U243 ( .INP(n450), .ZN(n734) );
  NOR2X0 U244 ( .IN1(n598), .IN2(n597), .QN(n9) );
  AND4X1 U245 ( .IN1(n570), .IN2(n569), .IN3(n572), .IN4(n568), .Q(n715) );
  OR2X1 U246 ( .IN1(n567), .IN2(n758), .Q(n790) );
  NAND3X0 U247 ( .IN1(n502), .IN2(n409), .IN3(n473), .QN(n491) );
  NOR2X0 U248 ( .IN1(n11), .IN2(n12), .QN(n216) );
  NOR2X0 U249 ( .IN1(n691), .IN2(n203), .QN(n11) );
  NOR2X0 U250 ( .IN1(exp_diff_value[3]), .IN2(exp_diff_value[2]), .QN(n356) );
  NOR2X0 U251 ( .IN1(n827), .IN2(n375), .QN(n357) );
  NOR2X0 U252 ( .IN1(exp_diff_value[1]), .IN2(n4), .QN(n178) );
  NOR2X0 U253 ( .IN1(exp_diff_value[1]), .IN2(exp_diff_value[0]), .QN(n332) );
  NOR2X0 U254 ( .IN1(exp_diff_value[0]), .IN2(n7), .QN(n177) );
  NOR2X0 U255 ( .IN1(n379), .IN2(n375), .QN(n355) );
  NOR2X0 U256 ( .IN1(exp_diff_value[3]), .IN2(n5), .QN(n212) );
  INVX0 U257 ( .INP(input_factor_01[15]), .ZN(n667) );
  INVX0 U258 ( .INP(input_factor_01[14]), .ZN(n661) );
  INVX0 U259 ( .INP(input_factor_01[13]), .ZN(n655) );
  INVX0 U260 ( .INP(input_factor_01[12]), .ZN(n649) );
  INVX0 U261 ( .INP(input_factor_01[11]), .ZN(n643) );
  INVX0 U262 ( .INP(input_factor_01[10]), .ZN(n637) );
  INVX0 U263 ( .INP(input_factor_01[9]), .ZN(n631) );
  INVX0 U264 ( .INP(input_factor_01[8]), .ZN(n627) );
  INVX0 U265 ( .INP(input_factor_01[7]), .ZN(n623) );
  INVX0 U266 ( .INP(input_factor_01[6]), .ZN(n619) );
  INVX0 U267 ( .INP(input_factor_01[5]), .ZN(n615) );
  INVX0 U268 ( .INP(input_factor_01[4]), .ZN(n611) );
  MUX21X1 U269 ( .IN1(sub_result[1]), .IN2(add_result[1]), .S(n511), .Q(n821)
         );
  INVX0 U270 ( .INP(n711), .ZN(n16) );
  AND4X1 U271 ( .IN1(n398), .IN2(n397), .IN3(n396), .IN4(n395), .Q(n8) );
  AO22X1 U272 ( .IN1(input_factor_01[30]), .IN2(rst_n), .IN3(n862), .IN4(
        larger_exponent[7]), .Q(n840) );
  INVX0 U274 ( .INP(input_factor_02[24]), .ZN(n32) );
  NOR2X0 U275 ( .IN1(input_factor_01[24]), .IN2(n32), .QN(n36) );
  NOR2X0 U276 ( .IN1(input_factor_01[25]), .IN2(n390), .QN(n17) );
  AO221X1 U277 ( .IN1(n19), .IN2(n36), .IN3(n19), .IN4(n18), .IN5(n17), .Q(n20) );
  OA221X1 U278 ( .IN1(n389), .IN2(input_factor_01[26]), .IN3(n389), .IN4(n22), 
        .IN5(input_factor_01[27]), .Q(n21) );
  OA221X1 U279 ( .IN1(n389), .IN2(input_factor_01[28]), .IN3(n389), .IN4(n21), 
        .IN5(input_factor_01[29]), .Q(n25) );
  OR2X1 U280 ( .IN1(input_factor_01[28]), .IN2(input_factor_01[26]), .Q(n552)
         );
  NOR3X0 U281 ( .IN1(n552), .IN2(input_factor_01[27]), .IN3(n22), .QN(n23) );
  NOR2X0 U282 ( .IN1(n23), .IN2(input_factor_02[29]), .QN(n24) );
  AO22X1 U283 ( .IN1(input_factor_02[18]), .IN2(n177), .IN3(
        input_factor_02[16]), .IN4(n332), .Q(n27) );
  NOR2X0 U284 ( .IN1(n7), .IN2(n4), .QN(n179) );
  AO22X1 U285 ( .IN1(input_factor_02[19]), .IN2(n179), .IN3(
        input_factor_02[17]), .IN4(n178), .Q(n26) );
  NOR2X0 U286 ( .IN1(n27), .IN2(n26), .QN(n219) );
  INVX0 U287 ( .INP(input_factor_02[22]), .ZN(n712) );
  INVX0 U288 ( .INP(input_factor_02[21]), .ZN(n704) );
  INVX0 U289 ( .INP(input_factor_02[20]), .ZN(n698) );
  AO222X1 U290 ( .IN1(n177), .IN2(n712), .IN3(n178), .IN4(n704), .IN5(n332), 
        .IN6(n698), .Q(n359) );
  MUX21X1 U291 ( .IN1(n219), .IN2(n359), .S(exp_diff_value[2]), .Q(n337) );
  INVX0 U292 ( .INP(input_factor_01[18]), .ZN(n685) );
  INVX0 U293 ( .INP(input_factor_01[17]), .ZN(n679) );
  OA22X1 U294 ( .IN1(n685), .IN2(n201), .IN3(n679), .IN4(n202), .Q(n29) );
  INVX0 U295 ( .INP(input_factor_01[19]), .ZN(n691) );
  INVX0 U296 ( .INP(input_factor_01[21]), .ZN(n703) );
  INVX0 U297 ( .INP(input_factor_01[20]), .ZN(n697) );
  AO222X1 U298 ( .IN1(n710), .IN2(n177), .IN3(n703), .IN4(n178), .IN5(n697), 
        .IN6(n332), .Q(n358) );
  MUX21X1 U299 ( .IN1(n216), .IN2(n358), .S(exp_diff_value[2]), .Q(n338) );
  OA22X1 U300 ( .IN1(input_factor_01[25]), .IN2(n390), .IN3(
        input_factor_01[28]), .IN4(n389), .Q(n40) );
  INVX0 U301 ( .INP(input_factor_01[29]), .ZN(n31) );
  NAND2X0 U302 ( .IN1(input_factor_01[27]), .IN2(input_factor_01[26]), .QN(n30) );
  AO222X1 U303 ( .IN1(input_factor_02[29]), .IN2(n31), .IN3(n389), .IN4(
        input_factor_01[29]), .IN5(n552), .IN6(n30), .Q(n35) );
  INVX0 U304 ( .INP(input_factor_01[23]), .ZN(n33) );
  AO222X1 U305 ( .IN1(input_factor_01[23]), .IN2(n390), .IN3(n33), .IN4(
        input_factor_02[23]), .IN5(input_factor_01[24]), .IN6(n32), .Q(n34) );
  NOR4X0 U306 ( .IN1(input_factor_01[30]), .IN2(n36), .IN3(n35), .IN4(n34), 
        .QN(n39) );
  NAND4X0 U307 ( .IN1(n40), .IN2(n39), .IN3(n38), .IN4(n37), .QN(n377) );
  OA22X1 U308 ( .IN1(n379), .IN2(n337), .IN3(n338), .IN4(n827), .Q(n64) );
  NOR3X0 U309 ( .IN1(exp_diff_value[5]), .IN2(exp_diff_value[6]), .IN3(
        exp_diff_value[7]), .QN(n41) );
  AND2X1 U310 ( .IN1(exp_diff_value[4]), .IN2(n41), .Q(n275) );
  INVX0 U311 ( .INP(input_factor_02[0]), .ZN(n76) );
  INVX0 U312 ( .INP(input_factor_01[1]), .ZN(n599) );
  AO222X1 U313 ( .IN1(input_factor_02[1]), .IN2(n599), .IN3(input_factor_02[1]), .IN4(n42), .IN5(n599), .IN6(n42), .Q(n43) );
  INVX0 U314 ( .INP(input_factor_01[2]), .ZN(n603) );
  AO222X1 U315 ( .IN1(input_factor_02[2]), .IN2(n43), .IN3(input_factor_02[2]), 
        .IN4(n603), .IN5(n43), .IN6(n603), .Q(n44) );
  INVX0 U316 ( .INP(input_factor_01[3]), .ZN(n607) );
  AO222X1 U317 ( .IN1(input_factor_02[3]), .IN2(n44), .IN3(input_factor_02[3]), 
        .IN4(n607), .IN5(n44), .IN6(n607), .Q(n45) );
  AO222X1 U318 ( .IN1(input_factor_02[4]), .IN2(n45), .IN3(input_factor_02[4]), 
        .IN4(n611), .IN5(n45), .IN6(n611), .Q(n46) );
  AO222X1 U319 ( .IN1(input_factor_02[5]), .IN2(n46), .IN3(input_factor_02[5]), 
        .IN4(n615), .IN5(n46), .IN6(n615), .Q(n47) );
  AO222X1 U320 ( .IN1(input_factor_02[6]), .IN2(n47), .IN3(input_factor_02[6]), 
        .IN4(n619), .IN5(n47), .IN6(n619), .Q(n48) );
  AO222X1 U321 ( .IN1(input_factor_02[7]), .IN2(n48), .IN3(input_factor_02[7]), 
        .IN4(n623), .IN5(n48), .IN6(n623), .Q(n49) );
  AO222X1 U322 ( .IN1(input_factor_02[8]), .IN2(n49), .IN3(input_factor_02[8]), 
        .IN4(n627), .IN5(n49), .IN6(n627), .Q(n50) );
  AO222X1 U323 ( .IN1(input_factor_02[9]), .IN2(n50), .IN3(input_factor_02[9]), 
        .IN4(n631), .IN5(n50), .IN6(n631), .Q(n51) );
  AO222X1 U324 ( .IN1(input_factor_02[10]), .IN2(n51), .IN3(
        input_factor_02[10]), .IN4(n637), .IN5(n51), .IN6(n637), .Q(n52) );
  AO222X1 U325 ( .IN1(input_factor_02[11]), .IN2(n52), .IN3(
        input_factor_02[11]), .IN4(n643), .IN5(n52), .IN6(n643), .Q(n53) );
  AO222X1 U326 ( .IN1(input_factor_02[12]), .IN2(n53), .IN3(
        input_factor_02[12]), .IN4(n649), .IN5(n53), .IN6(n649), .Q(n54) );
  AO222X1 U327 ( .IN1(input_factor_02[13]), .IN2(n54), .IN3(
        input_factor_02[13]), .IN4(n655), .IN5(n54), .IN6(n655), .Q(n55) );
  AO222X1 U328 ( .IN1(input_factor_02[14]), .IN2(n55), .IN3(
        input_factor_02[14]), .IN4(n661), .IN5(n55), .IN6(n661), .Q(n56) );
  AO222X1 U329 ( .IN1(input_factor_02[15]), .IN2(n56), .IN3(
        input_factor_02[15]), .IN4(n667), .IN5(n56), .IN6(n667), .Q(n57) );
  INVX0 U330 ( .INP(input_factor_01[16]), .ZN(n673) );
  AO222X1 U331 ( .IN1(input_factor_02[16]), .IN2(n57), .IN3(
        input_factor_02[16]), .IN4(n673), .IN5(n57), .IN6(n673), .Q(n58) );
  AO222X1 U332 ( .IN1(input_factor_02[17]), .IN2(n58), .IN3(
        input_factor_02[17]), .IN4(n679), .IN5(n58), .IN6(n679), .Q(n59) );
  AO222X1 U333 ( .IN1(input_factor_02[18]), .IN2(n59), .IN3(
        input_factor_02[18]), .IN4(n685), .IN5(n59), .IN6(n685), .Q(n60) );
  AO222X1 U334 ( .IN1(input_factor_02[19]), .IN2(n60), .IN3(
        input_factor_02[19]), .IN4(n691), .IN5(n60), .IN6(n691), .Q(n61) );
  AO222X1 U335 ( .IN1(input_factor_02[20]), .IN2(n61), .IN3(
        input_factor_02[20]), .IN4(n697), .IN5(n61), .IN6(n697), .Q(n62) );
  AO222X1 U336 ( .IN1(input_factor_02[21]), .IN2(n62), .IN3(
        input_factor_02[21]), .IN4(n703), .IN5(n62), .IN6(n703), .Q(n63) );
  AO222X1 U337 ( .IN1(input_factor_02[22]), .IN2(n63), .IN3(
        input_factor_02[22]), .IN4(n710), .IN5(n63), .IN6(n710), .Q(n65) );
  OA22X1 U338 ( .IN1(n64), .IN2(n182), .IN3(n76), .IN4(n380), .Q(n91) );
  INVX0 U339 ( .INP(n377), .ZN(n366) );
  INVX0 U340 ( .INP(n378), .ZN(n184) );
  OR4X1 U341 ( .IN1(exp_diff_value[4]), .IN2(exp_diff_value[5]), .IN3(
        exp_diff_value[6]), .IN4(exp_diff_value[7]), .Q(n375) );
  INVX0 U342 ( .INP(input_factor_01[0]), .ZN(n553) );
  OA22X1 U343 ( .IN1(n603), .IN2(n201), .IN3(n553), .IN4(n374), .Q(n67) );
  OA22X1 U344 ( .IN1(n607), .IN2(n203), .IN3(n599), .IN4(n202), .Q(n66) );
  OA22X1 U345 ( .IN1(n619), .IN2(n201), .IN3(n611), .IN4(n374), .Q(n69) );
  OA22X1 U346 ( .IN1(n623), .IN2(n203), .IN3(n615), .IN4(n202), .Q(n68) );
  OA22X1 U347 ( .IN1(n637), .IN2(n201), .IN3(n627), .IN4(n374), .Q(n71) );
  OA22X1 U348 ( .IN1(n643), .IN2(n203), .IN3(n631), .IN4(n202), .Q(n70) );
  OA22X1 U349 ( .IN1(n661), .IN2(n201), .IN3(n649), .IN4(n374), .Q(n73) );
  OA22X1 U350 ( .IN1(n667), .IN2(n203), .IN3(n655), .IN4(n202), .Q(n72) );
  MUX21X1 U351 ( .IN1(n213), .IN2(n215), .S(exp_diff_value[2]), .Q(n285) );
  AO222X1 U352 ( .IN1(n74), .IN2(n356), .IN3(n222), .IN4(n212), .IN5(n285), 
        .IN6(exp_diff_value[3]), .Q(n75) );
  INVX0 U353 ( .INP(input_factor_02[2]), .ZN(n604) );
  OA22X1 U354 ( .IN1(n604), .IN2(n201), .IN3(n76), .IN4(n374), .Q(n79) );
  INVX0 U355 ( .INP(input_factor_02[3]), .ZN(n608) );
  INVX0 U356 ( .INP(input_factor_02[1]), .ZN(n600) );
  OA22X1 U357 ( .IN1(n608), .IN2(n203), .IN3(n600), .IN4(n202), .Q(n77) );
  INVX0 U358 ( .INP(input_factor_02[6]), .ZN(n620) );
  INVX0 U359 ( .INP(input_factor_02[4]), .ZN(n612) );
  OA22X1 U360 ( .IN1(n620), .IN2(n201), .IN3(n612), .IN4(n374), .Q(n81) );
  INVX0 U361 ( .INP(input_factor_02[7]), .ZN(n624) );
  INVX0 U362 ( .INP(input_factor_02[5]), .ZN(n616) );
  OA22X1 U363 ( .IN1(n624), .IN2(n203), .IN3(n616), .IN4(n202), .Q(n80) );
  INVX0 U364 ( .INP(input_factor_02[10]), .ZN(n638) );
  INVX0 U365 ( .INP(input_factor_02[8]), .ZN(n628) );
  OA22X1 U366 ( .IN1(n638), .IN2(n201), .IN3(n628), .IN4(n374), .Q(n83) );
  INVX0 U367 ( .INP(input_factor_02[11]), .ZN(n644) );
  INVX0 U368 ( .INP(input_factor_02[9]), .ZN(n632) );
  OA22X1 U369 ( .IN1(n644), .IN2(n203), .IN3(n632), .IN4(n202), .Q(n82) );
  INVX0 U370 ( .INP(input_factor_02[14]), .ZN(n662) );
  INVX0 U371 ( .INP(input_factor_02[12]), .ZN(n650) );
  OA22X1 U372 ( .IN1(n662), .IN2(n201), .IN3(n650), .IN4(n374), .Q(n85) );
  INVX0 U373 ( .INP(input_factor_02[15]), .ZN(n668) );
  INVX0 U374 ( .INP(input_factor_02[13]), .ZN(n656) );
  OA22X1 U375 ( .IN1(n668), .IN2(n203), .IN3(n656), .IN4(n202), .Q(n84) );
  MUX21X1 U376 ( .IN1(n214), .IN2(n218), .S(exp_diff_value[2]), .Q(n283) );
  AO222X1 U377 ( .IN1(n86), .IN2(n356), .IN3(n221), .IN4(n212), .IN5(n283), 
        .IN6(exp_diff_value[3]), .Q(n87) );
  NAND4X0 U378 ( .IN1(n91), .IN2(n90), .IN3(n89), .IN4(n88), .QN(N152) );
  AO22X1 U379 ( .IN1(input_factor_02[19]), .IN2(n177), .IN3(
        input_factor_02[17]), .IN4(n332), .Q(n93) );
  AO22X1 U380 ( .IN1(input_factor_02[20]), .IN2(n179), .IN3(
        input_factor_02[18]), .IN4(n178), .Q(n92) );
  NOR2X0 U381 ( .IN1(n93), .IN2(n92), .QN(n235) );
  AO22X1 U382 ( .IN1(input_factor_02[22]), .IN2(n178), .IN3(
        input_factor_02[21]), .IN4(n4), .Q(n116) );
  NOR2X0 U383 ( .IN1(n177), .IN2(n116), .QN(n362) );
  MUX21X1 U384 ( .IN1(n235), .IN2(n362), .S(exp_diff_value[2]), .Q(n342) );
  AO22X1 U385 ( .IN1(input_factor_01[19]), .IN2(n177), .IN3(
        input_factor_01[17]), .IN4(n332), .Q(n118) );
  AO22X1 U386 ( .IN1(input_factor_01[20]), .IN2(n179), .IN3(
        input_factor_01[18]), .IN4(n178), .Q(n117) );
  NOR2X0 U387 ( .IN1(n118), .IN2(n117), .QN(n232) );
  AO22X1 U388 ( .IN1(input_factor_01[22]), .IN2(n178), .IN3(
        input_factor_01[21]), .IN4(n4), .Q(n119) );
  NOR2X0 U389 ( .IN1(n177), .IN2(n119), .QN(n363) );
  MUX21X1 U390 ( .IN1(n232), .IN2(n363), .S(exp_diff_value[2]), .Q(n341) );
  OA22X1 U391 ( .IN1(n379), .IN2(n342), .IN3(n341), .IN4(n827), .Q(n120) );
  OA22X1 U392 ( .IN1(n120), .IN2(n182), .IN3(n600), .IN4(n380), .Q(n145) );
  OA22X1 U393 ( .IN1(n607), .IN2(n201), .IN3(n599), .IN4(n374), .Q(n122) );
  OA22X1 U394 ( .IN1(n611), .IN2(n203), .IN3(n603), .IN4(n202), .Q(n121) );
  OA22X1 U395 ( .IN1(n623), .IN2(n201), .IN3(n615), .IN4(n374), .Q(n124) );
  OA22X1 U396 ( .IN1(n627), .IN2(n203), .IN3(n619), .IN4(n202), .Q(n123) );
  OA22X1 U397 ( .IN1(n643), .IN2(n201), .IN3(n631), .IN4(n374), .Q(n126) );
  OA22X1 U398 ( .IN1(n649), .IN2(n203), .IN3(n637), .IN4(n202), .Q(n125) );
  OA22X1 U399 ( .IN1(n667), .IN2(n201), .IN3(n655), .IN4(n374), .Q(n128) );
  OA22X1 U400 ( .IN1(n673), .IN2(n203), .IN3(n661), .IN4(n202), .Q(n127) );
  MUX21X1 U401 ( .IN1(n229), .IN2(n231), .S(exp_diff_value[2]), .Q(n292) );
  AO222X1 U402 ( .IN1(n129), .IN2(n356), .IN3(n238), .IN4(n212), .IN5(n292), 
        .IN6(exp_diff_value[3]), .Q(n130) );
  OA22X1 U403 ( .IN1(n608), .IN2(n201), .IN3(n600), .IN4(n374), .Q(n132) );
  OA22X1 U404 ( .IN1(n612), .IN2(n203), .IN3(n604), .IN4(n202), .Q(n131) );
  OA22X1 U405 ( .IN1(n624), .IN2(n201), .IN3(n616), .IN4(n374), .Q(n134) );
  OA22X1 U406 ( .IN1(n628), .IN2(n203), .IN3(n620), .IN4(n202), .Q(n133) );
  OA22X1 U407 ( .IN1(n644), .IN2(n201), .IN3(n632), .IN4(n374), .Q(n136) );
  OA22X1 U408 ( .IN1(n650), .IN2(n203), .IN3(n638), .IN4(n202), .Q(n135) );
  OA22X1 U409 ( .IN1(n668), .IN2(n201), .IN3(n656), .IN4(n374), .Q(n139) );
  INVX0 U410 ( .INP(input_factor_02[16]), .ZN(n674) );
  OA22X1 U411 ( .IN1(n674), .IN2(n203), .IN3(n662), .IN4(n202), .Q(n137) );
  MUX21X1 U412 ( .IN1(n230), .IN2(n234), .S(exp_diff_value[2]), .Q(n290) );
  AO222X1 U413 ( .IN1(n140), .IN2(n356), .IN3(n237), .IN4(n212), .IN5(n290), 
        .IN6(exp_diff_value[3]), .Q(n141) );
  NAND4X0 U414 ( .IN1(n145), .IN2(n144), .IN3(n143), .IN4(n142), .QN(N153) );
  AO22X1 U415 ( .IN1(input_factor_02[20]), .IN2(n177), .IN3(
        input_factor_02[18]), .IN4(n332), .Q(n147) );
  AO22X1 U416 ( .IN1(input_factor_02[21]), .IN2(n179), .IN3(
        input_factor_02[19]), .IN4(n178), .Q(n146) );
  NOR2X0 U417 ( .IN1(n147), .IN2(n146), .QN(n251) );
  AO21X1 U418 ( .IN1(n712), .IN2(n4), .IN3(exp_diff_value[1]), .Q(n370) );
  MUX21X1 U419 ( .IN1(n251), .IN2(n370), .S(exp_diff_value[2]), .Q(n345) );
  AO22X1 U420 ( .IN1(input_factor_01[20]), .IN2(n177), .IN3(
        input_factor_01[18]), .IN4(n332), .Q(n149) );
  AO22X1 U421 ( .IN1(input_factor_01[21]), .IN2(n179), .IN3(
        input_factor_01[19]), .IN4(n178), .Q(n148) );
  NOR2X0 U422 ( .IN1(n149), .IN2(n148), .QN(n248) );
  AO21X1 U423 ( .IN1(n710), .IN2(n4), .IN3(exp_diff_value[1]), .Q(n368) );
  MUX21X1 U424 ( .IN1(n248), .IN2(n368), .S(exp_diff_value[2]), .Q(n346) );
  OA22X1 U425 ( .IN1(n379), .IN2(n345), .IN3(n346), .IN4(n827), .Q(n150) );
  OA22X1 U426 ( .IN1(n150), .IN2(n182), .IN3(n604), .IN4(n380), .Q(n174) );
  OA22X1 U427 ( .IN1(n611), .IN2(n201), .IN3(n603), .IN4(n374), .Q(n152) );
  OA22X1 U428 ( .IN1(n615), .IN2(n203), .IN3(n607), .IN4(n202), .Q(n151) );
  OA22X1 U429 ( .IN1(n627), .IN2(n201), .IN3(n619), .IN4(n374), .Q(n154) );
  OA22X1 U430 ( .IN1(n631), .IN2(n203), .IN3(n623), .IN4(n202), .Q(n153) );
  OA22X1 U431 ( .IN1(n649), .IN2(n201), .IN3(n637), .IN4(n374), .Q(n156) );
  OA22X1 U432 ( .IN1(n655), .IN2(n203), .IN3(n643), .IN4(n202), .Q(n155) );
  OA22X1 U433 ( .IN1(n673), .IN2(n201), .IN3(n661), .IN4(n374), .Q(n158) );
  OA22X1 U434 ( .IN1(n679), .IN2(n203), .IN3(n667), .IN4(n202), .Q(n157) );
  MUX21X1 U435 ( .IN1(n245), .IN2(n247), .S(exp_diff_value[2]), .Q(n299) );
  AO222X1 U436 ( .IN1(n159), .IN2(n356), .IN3(n254), .IN4(n212), .IN5(n299), 
        .IN6(exp_diff_value[3]), .Q(n160) );
  OA22X1 U437 ( .IN1(n612), .IN2(n201), .IN3(n604), .IN4(n374), .Q(n162) );
  OA22X1 U438 ( .IN1(n616), .IN2(n203), .IN3(n608), .IN4(n202), .Q(n161) );
  OA22X1 U439 ( .IN1(n628), .IN2(n201), .IN3(n620), .IN4(n374), .Q(n164) );
  OA22X1 U440 ( .IN1(n632), .IN2(n203), .IN3(n624), .IN4(n202), .Q(n163) );
  OA22X1 U441 ( .IN1(n650), .IN2(n201), .IN3(n638), .IN4(n374), .Q(n166) );
  OA22X1 U442 ( .IN1(n656), .IN2(n203), .IN3(n644), .IN4(n202), .Q(n165) );
  OA22X1 U443 ( .IN1(n674), .IN2(n201), .IN3(n662), .IN4(n374), .Q(n168) );
  INVX0 U444 ( .INP(input_factor_02[17]), .ZN(n680) );
  OA22X1 U445 ( .IN1(n680), .IN2(n203), .IN3(n668), .IN4(n202), .Q(n167) );
  MUX21X1 U446 ( .IN1(n246), .IN2(n250), .S(exp_diff_value[2]), .Q(n297) );
  AO222X1 U447 ( .IN1(n169), .IN2(n356), .IN3(n253), .IN4(n212), .IN5(n297), 
        .IN6(exp_diff_value[3]), .Q(n170) );
  NAND4X0 U448 ( .IN1(n174), .IN2(n173), .IN3(n172), .IN4(n171), .QN(N154) );
  AO22X1 U449 ( .IN1(input_factor_02[21]), .IN2(n177), .IN3(
        input_factor_02[19]), .IN4(n332), .Q(n176) );
  AO22X1 U450 ( .IN1(input_factor_02[22]), .IN2(n179), .IN3(
        input_factor_02[20]), .IN4(n178), .Q(n175) );
  NOR2X0 U451 ( .IN1(n176), .IN2(n175), .QN(n271) );
  MUX21X1 U452 ( .IN1(n271), .IN2(n374), .S(exp_diff_value[2]), .Q(n350) );
  AO22X1 U453 ( .IN1(input_factor_01[21]), .IN2(n177), .IN3(
        input_factor_01[19]), .IN4(n332), .Q(n181) );
  AO22X1 U454 ( .IN1(input_factor_01[22]), .IN2(n179), .IN3(
        input_factor_01[20]), .IN4(n178), .Q(n180) );
  NOR2X0 U455 ( .IN1(n181), .IN2(n180), .QN(n268) );
  MUX21X1 U456 ( .IN1(n268), .IN2(n374), .S(exp_diff_value[2]), .Q(n352) );
  OA22X1 U457 ( .IN1(n379), .IN2(n350), .IN3(n352), .IN4(n827), .Q(n183) );
  OA22X1 U458 ( .IN1(n183), .IN2(n182), .IN3(n608), .IN4(n380), .Q(n211) );
  OA22X1 U459 ( .IN1(n615), .IN2(n201), .IN3(n607), .IN4(n374), .Q(n186) );
  OA22X1 U460 ( .IN1(n619), .IN2(n203), .IN3(n611), .IN4(n202), .Q(n185) );
  OA22X1 U461 ( .IN1(n631), .IN2(n201), .IN3(n623), .IN4(n374), .Q(n188) );
  OA22X1 U462 ( .IN1(n637), .IN2(n203), .IN3(n627), .IN4(n202), .Q(n187) );
  OA22X1 U463 ( .IN1(n655), .IN2(n201), .IN3(n643), .IN4(n374), .Q(n190) );
  OA22X1 U464 ( .IN1(n661), .IN2(n203), .IN3(n649), .IN4(n202), .Q(n189) );
  OA22X1 U465 ( .IN1(n679), .IN2(n201), .IN3(n667), .IN4(n374), .Q(n192) );
  OA22X1 U466 ( .IN1(n685), .IN2(n203), .IN3(n673), .IN4(n202), .Q(n191) );
  MUX21X1 U467 ( .IN1(n263), .IN2(n267), .S(exp_diff_value[2]), .Q(n306) );
  AO222X1 U468 ( .IN1(n193), .IN2(n356), .IN3(n274), .IN4(n212), .IN5(n306), 
        .IN6(exp_diff_value[3]), .Q(n194) );
  OA22X1 U469 ( .IN1(n616), .IN2(n201), .IN3(n608), .IN4(n374), .Q(n196) );
  OA22X1 U470 ( .IN1(n620), .IN2(n203), .IN3(n612), .IN4(n202), .Q(n195) );
  OA22X1 U471 ( .IN1(n632), .IN2(n201), .IN3(n624), .IN4(n374), .Q(n198) );
  OA22X1 U472 ( .IN1(n638), .IN2(n203), .IN3(n628), .IN4(n202), .Q(n197) );
  OA22X1 U473 ( .IN1(n656), .IN2(n201), .IN3(n644), .IN4(n374), .Q(n200) );
  OA22X1 U474 ( .IN1(n662), .IN2(n203), .IN3(n650), .IN4(n202), .Q(n199) );
  OA22X1 U475 ( .IN1(n680), .IN2(n201), .IN3(n668), .IN4(n374), .Q(n205) );
  INVX0 U476 ( .INP(input_factor_02[18]), .ZN(n686) );
  OA22X1 U477 ( .IN1(n686), .IN2(n203), .IN3(n674), .IN4(n202), .Q(n204) );
  MUX21X1 U478 ( .IN1(n265), .IN2(n270), .S(exp_diff_value[2]), .Q(n304) );
  AO222X1 U479 ( .IN1(n206), .IN2(n356), .IN3(n273), .IN4(n212), .IN5(n304), 
        .IN6(exp_diff_value[3]), .Q(n207) );
  NAND4X0 U480 ( .IN1(n211), .IN2(n210), .IN3(n209), .IN4(n208), .QN(N155) );
  AND2X1 U481 ( .IN1(n212), .IN2(n355), .Q(n266) );
  AND2X1 U482 ( .IN1(n357), .IN2(n212), .Q(n264) );
  AOI22X1 U483 ( .IN1(n266), .IN2(n214), .IN3(n264), .IN4(n213), .QN(n228) );
  INVX0 U484 ( .INP(n215), .ZN(n217) );
  MUX21X1 U485 ( .IN1(n217), .IN2(n216), .S(exp_diff_value[2]), .Q(n312) );
  INVX0 U486 ( .INP(n218), .ZN(n220) );
  MUX21X1 U487 ( .IN1(n220), .IN2(n219), .S(exp_diff_value[2]), .Q(n311) );
  OA22X1 U488 ( .IN1(n330), .IN2(n312), .IN3(n331), .IN4(n311), .Q(n227) );
  OA22X1 U489 ( .IN1(n612), .IN2(n380), .IN3(n611), .IN4(n378), .Q(n226) );
  AOI22X1 U490 ( .IN1(n357), .IN2(n222), .IN3(n355), .IN4(n221), .QN(n224) );
  OA22X1 U491 ( .IN1(n359), .IN2(n256), .IN3(n358), .IN4(n255), .Q(n223) );
  INVX0 U492 ( .INP(n356), .ZN(n373) );
  AO21X1 U493 ( .IN1(n224), .IN2(n223), .IN3(n373), .Q(n225) );
  NAND4X0 U494 ( .IN1(n228), .IN2(n227), .IN3(n226), .IN4(n225), .QN(N156) );
  AOI22X1 U495 ( .IN1(n266), .IN2(n230), .IN3(n264), .IN4(n229), .QN(n244) );
  INVX0 U496 ( .INP(n231), .ZN(n233) );
  MUX21X1 U497 ( .IN1(n233), .IN2(n232), .S(exp_diff_value[2]), .Q(n317) );
  INVX0 U498 ( .INP(n234), .ZN(n236) );
  MUX21X1 U499 ( .IN1(n236), .IN2(n235), .S(exp_diff_value[2]), .Q(n316) );
  OA22X1 U500 ( .IN1(n330), .IN2(n317), .IN3(n331), .IN4(n316), .Q(n243) );
  OA22X1 U501 ( .IN1(n616), .IN2(n380), .IN3(n615), .IN4(n378), .Q(n242) );
  AOI22X1 U502 ( .IN1(n357), .IN2(n238), .IN3(n355), .IN4(n237), .QN(n240) );
  OA22X1 U503 ( .IN1(n363), .IN2(n255), .IN3(n362), .IN4(n256), .Q(n239) );
  AO21X1 U504 ( .IN1(n240), .IN2(n239), .IN3(n373), .Q(n241) );
  NAND4X0 U505 ( .IN1(n244), .IN2(n243), .IN3(n242), .IN4(n241), .QN(N157) );
  AOI22X1 U506 ( .IN1(n266), .IN2(n246), .IN3(n264), .IN4(n245), .QN(n262) );
  INVX0 U507 ( .INP(n247), .ZN(n249) );
  MUX21X1 U508 ( .IN1(n249), .IN2(n248), .S(exp_diff_value[2]), .Q(n322) );
  INVX0 U509 ( .INP(n250), .ZN(n252) );
  MUX21X1 U510 ( .IN1(n252), .IN2(n251), .S(exp_diff_value[2]), .Q(n321) );
  OA22X1 U511 ( .IN1(n330), .IN2(n322), .IN3(n331), .IN4(n321), .Q(n261) );
  OA22X1 U512 ( .IN1(n620), .IN2(n380), .IN3(n619), .IN4(n378), .Q(n260) );
  AOI22X1 U513 ( .IN1(n357), .IN2(n254), .IN3(n355), .IN4(n253), .QN(n258) );
  OA22X1 U514 ( .IN1(n370), .IN2(n256), .IN3(n368), .IN4(n255), .Q(n257) );
  AO21X1 U515 ( .IN1(n258), .IN2(n257), .IN3(n373), .Q(n259) );
  NAND4X0 U516 ( .IN1(n262), .IN2(n261), .IN3(n260), .IN4(n259), .QN(N158) );
  AOI22X1 U517 ( .IN1(n266), .IN2(n265), .IN3(n264), .IN4(n263), .QN(n282) );
  INVX0 U518 ( .INP(n267), .ZN(n269) );
  MUX21X1 U519 ( .IN1(n269), .IN2(n268), .S(exp_diff_value[2]), .Q(n329) );
  INVX0 U520 ( .INP(n270), .ZN(n272) );
  MUX21X1 U521 ( .IN1(n272), .IN2(n271), .S(exp_diff_value[2]), .Q(n328) );
  OA22X1 U522 ( .IN1(n330), .IN2(n329), .IN3(n331), .IN4(n328), .Q(n281) );
  OA22X1 U523 ( .IN1(n624), .IN2(n380), .IN3(n623), .IN4(n378), .Q(n280) );
  AOI22X1 U524 ( .IN1(n357), .IN2(n274), .IN3(n355), .IN4(n273), .QN(n278) );
  NAND3X0 U525 ( .IN1(n276), .IN2(n332), .IN3(n275), .QN(n277) );
  AO21X1 U526 ( .IN1(n278), .IN2(n277), .IN3(n373), .Q(n279) );
  NAND4X0 U527 ( .IN1(n282), .IN2(n281), .IN3(n280), .IN4(n279), .QN(N159) );
  INVX0 U528 ( .INP(n283), .ZN(n284) );
  OA22X1 U529 ( .IN1(n337), .IN2(n331), .IN3(n349), .IN4(n284), .Q(n289) );
  INVX0 U530 ( .INP(n285), .ZN(n286) );
  OA22X1 U531 ( .IN1(n338), .IN2(n330), .IN3(n351), .IN4(n286), .Q(n288) );
  OA22X1 U532 ( .IN1(n628), .IN2(n380), .IN3(n627), .IN4(n378), .Q(n287) );
  NAND3X0 U533 ( .IN1(n289), .IN2(n288), .IN3(n287), .QN(N160) );
  INVX0 U534 ( .INP(n290), .ZN(n291) );
  OA22X1 U535 ( .IN1(n342), .IN2(n331), .IN3(n291), .IN4(n349), .Q(n296) );
  INVX0 U536 ( .INP(n292), .ZN(n293) );
  OA22X1 U537 ( .IN1(n341), .IN2(n330), .IN3(n293), .IN4(n351), .Q(n295) );
  OA22X1 U538 ( .IN1(n632), .IN2(n380), .IN3(n631), .IN4(n378), .Q(n294) );
  NAND3X0 U539 ( .IN1(n296), .IN2(n295), .IN3(n294), .QN(N161) );
  INVX0 U540 ( .INP(n297), .ZN(n298) );
  OA22X1 U541 ( .IN1(n345), .IN2(n331), .IN3(n349), .IN4(n298), .Q(n303) );
  INVX0 U542 ( .INP(n299), .ZN(n300) );
  OA22X1 U543 ( .IN1(n346), .IN2(n330), .IN3(n351), .IN4(n300), .Q(n302) );
  OA22X1 U544 ( .IN1(n638), .IN2(n380), .IN3(n637), .IN4(n378), .Q(n301) );
  NAND3X0 U545 ( .IN1(n303), .IN2(n302), .IN3(n301), .QN(N162) );
  INVX0 U546 ( .INP(n304), .ZN(n305) );
  OA22X1 U547 ( .IN1(n350), .IN2(n331), .IN3(n349), .IN4(n305), .Q(n310) );
  INVX0 U548 ( .INP(n306), .ZN(n307) );
  OA22X1 U549 ( .IN1(n352), .IN2(n330), .IN3(n351), .IN4(n307), .Q(n309) );
  OA22X1 U550 ( .IN1(n644), .IN2(n380), .IN3(n643), .IN4(n378), .Q(n308) );
  NAND3X0 U551 ( .IN1(n310), .IN2(n309), .IN3(n308), .QN(N163) );
  OA22X1 U552 ( .IN1(n312), .IN2(n351), .IN3(n311), .IN4(n349), .Q(n315) );
  OR2X1 U553 ( .IN1(n331), .IN2(exp_diff_value[2]), .Q(n324) );
  OR2X1 U554 ( .IN1(n330), .IN2(exp_diff_value[2]), .Q(n323) );
  OA22X1 U555 ( .IN1(n359), .IN2(n324), .IN3(n358), .IN4(n323), .Q(n314) );
  OA22X1 U556 ( .IN1(n650), .IN2(n380), .IN3(n649), .IN4(n378), .Q(n313) );
  NAND3X0 U557 ( .IN1(n315), .IN2(n314), .IN3(n313), .QN(N164) );
  OA22X1 U558 ( .IN1(n317), .IN2(n351), .IN3(n316), .IN4(n349), .Q(n320) );
  OA22X1 U559 ( .IN1(n363), .IN2(n323), .IN3(n362), .IN4(n324), .Q(n319) );
  OA22X1 U560 ( .IN1(n656), .IN2(n380), .IN3(n655), .IN4(n378), .Q(n318) );
  NAND3X0 U561 ( .IN1(n320), .IN2(n319), .IN3(n318), .QN(N165) );
  OA22X1 U562 ( .IN1(n322), .IN2(n351), .IN3(n321), .IN4(n349), .Q(n327) );
  OA22X1 U563 ( .IN1(n370), .IN2(n324), .IN3(n368), .IN4(n323), .Q(n326) );
  OA22X1 U564 ( .IN1(n662), .IN2(n380), .IN3(n661), .IN4(n378), .Q(n325) );
  NAND3X0 U565 ( .IN1(n327), .IN2(n326), .IN3(n325), .QN(N166) );
  OA22X1 U566 ( .IN1(n329), .IN2(n351), .IN3(n328), .IN4(n349), .Q(n336) );
  OA22X1 U567 ( .IN1(n668), .IN2(n380), .IN3(n667), .IN4(n378), .Q(n335) );
  NAND3X0 U568 ( .IN1(n333), .IN2(n5), .IN3(n332), .QN(n334) );
  NAND3X0 U569 ( .IN1(n336), .IN2(n335), .IN3(n334), .QN(N167) );
  OA22X1 U570 ( .IN1(n338), .IN2(n351), .IN3(n337), .IN4(n349), .Q(n340) );
  OA22X1 U571 ( .IN1(n674), .IN2(n380), .IN3(n673), .IN4(n378), .Q(n339) );
  OA22X1 U572 ( .IN1(n342), .IN2(n349), .IN3(n341), .IN4(n351), .Q(n344) );
  OA22X1 U573 ( .IN1(n680), .IN2(n380), .IN3(n679), .IN4(n378), .Q(n343) );
  OA22X1 U574 ( .IN1(n346), .IN2(n351), .IN3(n345), .IN4(n349), .Q(n348) );
  OA22X1 U575 ( .IN1(n686), .IN2(n380), .IN3(n685), .IN4(n378), .Q(n347) );
  OA22X1 U576 ( .IN1(n352), .IN2(n351), .IN3(n350), .IN4(n349), .Q(n354) );
  INVX0 U577 ( .INP(input_factor_02[19]), .ZN(n692) );
  OA22X1 U578 ( .IN1(n692), .IN2(n380), .IN3(n691), .IN4(n378), .Q(n353) );
  OA22X1 U579 ( .IN1(n359), .IN2(n369), .IN3(n358), .IN4(n367), .Q(n361) );
  OA22X1 U580 ( .IN1(n698), .IN2(n380), .IN3(n697), .IN4(n378), .Q(n360) );
  OA22X1 U581 ( .IN1(n363), .IN2(n367), .IN3(n362), .IN4(n369), .Q(n365) );
  OA22X1 U582 ( .IN1(n704), .IN2(n380), .IN3(n703), .IN4(n378), .Q(n364) );
  NAND3X0 U583 ( .IN1(input_factor_01[22]), .IN2(n366), .IN3(
        input_factor_02[22]), .QN(n372) );
  OA22X1 U584 ( .IN1(n370), .IN2(n369), .IN3(n368), .IN4(n367), .Q(n371) );
  OR3X1 U585 ( .IN1(n375), .IN2(n374), .IN3(n373), .Q(n376) );
  AO22X1 U586 ( .IN1(input_factor_02[0]), .IN2(n401), .IN3(input_factor_01[0]), 
        .IN4(n399), .Q(N176) );
  AO22X1 U587 ( .IN1(input_factor_02[1]), .IN2(n401), .IN3(input_factor_01[1]), 
        .IN4(n399), .Q(N177) );
  AO22X1 U588 ( .IN1(input_factor_02[2]), .IN2(n401), .IN3(input_factor_01[2]), 
        .IN4(n399), .Q(N178) );
  AO22X1 U589 ( .IN1(input_factor_02[3]), .IN2(n401), .IN3(input_factor_01[3]), 
        .IN4(n399), .Q(N179) );
  AO22X1 U590 ( .IN1(input_factor_02[4]), .IN2(n401), .IN3(input_factor_01[4]), 
        .IN4(n399), .Q(N180) );
  AO22X1 U591 ( .IN1(input_factor_02[5]), .IN2(n401), .IN3(input_factor_01[5]), 
        .IN4(n399), .Q(N181) );
  AO22X1 U592 ( .IN1(input_factor_02[6]), .IN2(n401), .IN3(input_factor_01[6]), 
        .IN4(n399), .Q(N182) );
  AO22X1 U593 ( .IN1(input_factor_02[7]), .IN2(n401), .IN3(input_factor_01[7]), 
        .IN4(n399), .Q(N183) );
  AO22X1 U594 ( .IN1(input_factor_02[8]), .IN2(n401), .IN3(input_factor_01[8]), 
        .IN4(n399), .Q(N184) );
  AO22X1 U595 ( .IN1(input_factor_02[9]), .IN2(n401), .IN3(input_factor_01[9]), 
        .IN4(n399), .Q(N185) );
  AO22X1 U596 ( .IN1(input_factor_02[10]), .IN2(n401), .IN3(
        input_factor_01[10]), .IN4(n399), .Q(N186) );
  AO22X1 U597 ( .IN1(input_factor_02[11]), .IN2(n401), .IN3(
        input_factor_01[11]), .IN4(n399), .Q(N187) );
  AO22X1 U598 ( .IN1(input_factor_02[12]), .IN2(n401), .IN3(
        input_factor_01[12]), .IN4(n399), .Q(N188) );
  AO22X1 U599 ( .IN1(input_factor_02[13]), .IN2(n401), .IN3(
        input_factor_01[13]), .IN4(n399), .Q(N189) );
  AO22X1 U600 ( .IN1(input_factor_02[14]), .IN2(n401), .IN3(
        input_factor_01[14]), .IN4(n399), .Q(N190) );
  AO22X1 U601 ( .IN1(input_factor_02[15]), .IN2(n401), .IN3(
        input_factor_01[15]), .IN4(n399), .Q(N191) );
  AO22X1 U602 ( .IN1(input_factor_02[16]), .IN2(n401), .IN3(
        input_factor_01[16]), .IN4(n399), .Q(N192) );
  AO22X1 U603 ( .IN1(input_factor_02[17]), .IN2(n401), .IN3(
        input_factor_01[17]), .IN4(n399), .Q(N193) );
  AO22X1 U604 ( .IN1(input_factor_02[18]), .IN2(n401), .IN3(
        input_factor_01[18]), .IN4(n399), .Q(N194) );
  AO22X1 U605 ( .IN1(input_factor_02[19]), .IN2(n401), .IN3(
        input_factor_01[19]), .IN4(n399), .Q(N195) );
  AO22X1 U606 ( .IN1(input_factor_02[20]), .IN2(n401), .IN3(
        input_factor_01[20]), .IN4(n399), .Q(N196) );
  AO22X1 U607 ( .IN1(input_factor_02[21]), .IN2(n401), .IN3(
        input_factor_01[21]), .IN4(n399), .Q(N197) );
  AO22X1 U608 ( .IN1(input_factor_02[22]), .IN2(n401), .IN3(
        input_factor_01[22]), .IN4(n399), .Q(N198) );
  MUX21X1 U609 ( .IN1(sub_result[0]), .IN2(add_result[0]), .S(n511), .Q(n823)
         );
  MUX21X1 U610 ( .IN1(sub_result[2]), .IN2(add_result[2]), .S(n511), .Q(n801)
         );
  MUX21X1 U611 ( .IN1(sub_result[3]), .IN2(add_result[3]), .S(n511), .Q(n793)
         );
  MUX21X1 U612 ( .IN1(sub_result[4]), .IN2(add_result[4]), .S(n511), .Q(n802)
         );
  MUX21X1 U613 ( .IN1(sub_result[5]), .IN2(add_result[5]), .S(n511), .Q(n794)
         );
  MUX21X1 U614 ( .IN1(sub_result[6]), .IN2(add_result[6]), .S(n511), .Q(n769)
         );
  MUX21X1 U615 ( .IN1(sub_result[7]), .IN2(add_result[7]), .S(n511), .Q(n761)
         );
  MUX21X1 U616 ( .IN1(sub_result[9]), .IN2(add_result[9]), .S(n511), .Q(n745)
         );
  MUX21X1 U617 ( .IN1(sub_result[10]), .IN2(add_result[10]), .S(n511), .Q(n737) );
  NOR4X0 U618 ( .IN1(add_result[15]), .IN2(add_result[14]), .IN3(
        add_result[13]), .IN4(n14), .QN(n520) );
  NOR4X0 U619 ( .IN1(n511), .IN2(sub_result[14]), .IN3(sub_result[15]), .IN4(
        sub_result[13]), .QN(n518) );
  NOR2X0 U620 ( .IN1(n520), .IN2(n518), .QN(n385) );
  MUX21X1 U621 ( .IN1(sub_result[11]), .IN2(add_result[11]), .S(n511), .Q(n729) );
  MUX21X1 U622 ( .IN1(sub_result[16]), .IN2(add_result[16]), .S(n13), .Q(n404)
         );
  MUX21X1 U623 ( .IN1(sub_result[17]), .IN2(add_result[17]), .S(n13), .Q(n473)
         );
  MUX21X1 U624 ( .IN1(sub_result[20]), .IN2(add_result[20]), .S(n13), .Q(n407)
         );
  INVX0 U625 ( .INP(n407), .ZN(n500) );
  MUX21X1 U626 ( .IN1(sub_result[22]), .IN2(add_result[22]), .S(n13), .Q(n408)
         );
  INVX0 U627 ( .INP(n408), .ZN(n382) );
  MUX21X1 U628 ( .IN1(sub_result[23]), .IN2(add_result[23]), .S(n13), .Q(n403)
         );
  MUX21X1 U629 ( .IN1(sub_result[21]), .IN2(add_result[21]), .S(n13), .Q(n410)
         );
  NOR2X0 U630 ( .IN1(n411), .IN2(n410), .QN(n412) );
  MUX21X1 U631 ( .IN1(sub_result[19]), .IN2(add_result[19]), .S(n13), .Q(n482)
         );
  NOR2X0 U632 ( .IN1(n383), .IN2(n482), .QN(n409) );
  MUX21X1 U633 ( .IN1(sub_result[18]), .IN2(add_result[18]), .S(n13), .Q(n406)
         );
  NOR2X0 U634 ( .IN1(n473), .IN2(n384), .QN(n405) );
  MUX21X1 U635 ( .IN1(sub_result[12]), .IN2(add_result[12]), .S(n13), .Q(n450)
         );
  NOR4X0 U636 ( .IN1(n385), .IN2(n729), .IN3(n564), .IN4(n450), .QN(n724) );
  MUX21X1 U637 ( .IN1(sub_result[8]), .IN2(add_result[8]), .S(n13), .Q(n753)
         );
  NOR3X0 U638 ( .IN1(n745), .IN2(n567), .IN3(n753), .QN(n525) );
  NOR2X0 U639 ( .IN1(n769), .IN2(n386), .QN(n524) );
  NOR2X0 U640 ( .IN1(n802), .IN2(n387), .QN(n532) );
  NOR2X0 U641 ( .IN1(n801), .IN2(n388), .QN(n526) );
  NAND3X0 U642 ( .IN1(n815), .IN2(n807), .IN3(n526), .QN(n562) );
  NOR4X0 U643 ( .IN1(input_factor_02[15]), .IN2(input_factor_02[13]), .IN3(
        input_factor_02[11]), .IN4(input_factor_02[10]), .QN(n398) );
  NOR4X0 U644 ( .IN1(input_factor_02[22]), .IN2(input_factor_02[2]), .IN3(
        input_factor_02[0]), .IN4(input_factor_02[1]), .QN(n397) );
  NOR4X0 U645 ( .IN1(input_factor_02[21]), .IN2(input_factor_02[20]), .IN3(
        input_factor_02[19]), .IN4(input_factor_02[17]), .QN(n396) );
  NOR4X0 U646 ( .IN1(input_factor_02[31]), .IN2(input_factor_02[24]), .IN3(
        input_factor_02[18]), .IN4(input_factor_02[16]), .QN(n391) );
  NAND4X0 U647 ( .IN1(n391), .IN2(n390), .IN3(n389), .IN4(n662), .QN(n394) );
  NOR4X0 U648 ( .IN1(input_factor_02[9]), .IN2(input_factor_02[7]), .IN3(
        input_factor_02[6]), .IN4(input_factor_02[5]), .QN(n392) );
  NAND3X0 U649 ( .IN1(n392), .IN2(n612), .IN3(n608), .QN(n393) );
  NOR4X0 U650 ( .IN1(input_factor_02[12]), .IN2(input_factor_02[8]), .IN3(n394), .IN4(n393), .QN(n395) );
  OR2X1 U651 ( .IN1(n399), .IN2(n8), .Q(n400) );
  AO222X1 U652 ( .IN1(input_factor_02[31]), .IN2(input_factor_01[31]), .IN3(
        input_factor_02[31]), .IN4(n401), .IN5(input_factor_01[31]), .IN6(n400), .Q(n402) );
  AND2X1 U653 ( .IN1(n562), .IN2(n402), .Q(N211) );
  MUX21X1 U654 ( .IN1(n823), .IN2(n821), .S(add_sub_result_24_), .Q(N226) );
  MUX21X1 U655 ( .IN1(n821), .IN2(n801), .S(add_sub_result_24_), .Q(N227) );
  MUX21X1 U656 ( .IN1(n801), .IN2(n793), .S(add_sub_result_24_), .Q(N228) );
  MUX21X1 U657 ( .IN1(n793), .IN2(n802), .S(add_sub_result_24_), .Q(N229) );
  MUX21X1 U658 ( .IN1(n802), .IN2(n794), .S(add_sub_result_24_), .Q(N230) );
  MUX21X1 U659 ( .IN1(n794), .IN2(n769), .S(add_sub_result_24_), .Q(N231) );
  MUX21X1 U660 ( .IN1(n769), .IN2(n761), .S(add_sub_result_24_), .Q(N232) );
  MUX21X1 U661 ( .IN1(n761), .IN2(n753), .S(add_sub_result_24_), .Q(N233) );
  MUX21X1 U662 ( .IN1(n753), .IN2(n745), .S(add_sub_result_24_), .Q(N234) );
  MUX21X1 U663 ( .IN1(n745), .IN2(n737), .S(add_sub_result_24_), .Q(N235) );
  MUX21X1 U664 ( .IN1(n737), .IN2(n729), .S(add_sub_result_24_), .Q(N236) );
  MUX21X1 U665 ( .IN1(n729), .IN2(n450), .S(add_sub_result_24_), .Q(N237) );
  MUX21X1 U666 ( .IN1(sub_result[13]), .IN2(add_result[13]), .S(n13), .Q(n455)
         );
  MUX21X1 U667 ( .IN1(n450), .IN2(n455), .S(add_sub_result_24_), .Q(N238) );
  MUX21X1 U668 ( .IN1(sub_result[14]), .IN2(add_result[14]), .S(n13), .Q(n509)
         );
  MUX21X1 U669 ( .IN1(n455), .IN2(n509), .S(add_sub_result_24_), .Q(N239) );
  MUX21X1 U670 ( .IN1(sub_result[15]), .IN2(add_result[15]), .S(n13), .Q(n464)
         );
  MUX21X1 U671 ( .IN1(n509), .IN2(n464), .S(add_sub_result_24_), .Q(N240) );
  MUX21X1 U672 ( .IN1(n464), .IN2(n404), .S(add_sub_result_24_), .Q(N241) );
  MUX21X1 U673 ( .IN1(n404), .IN2(n473), .S(add_sub_result_24_), .Q(N242) );
  MUX21X1 U674 ( .IN1(n473), .IN2(n406), .S(add_sub_result_24_), .Q(N243) );
  MUX21X1 U675 ( .IN1(n406), .IN2(n482), .S(add_sub_result_24_), .Q(N244) );
  MUX21X1 U676 ( .IN1(n482), .IN2(n407), .S(add_sub_result_24_), .Q(N245) );
  MUX21X1 U677 ( .IN1(n407), .IN2(n410), .S(add_sub_result_24_), .Q(N246) );
  MUX21X1 U678 ( .IN1(n410), .IN2(n408), .S(add_sub_result_24_), .Q(N247) );
  MUX21X1 U679 ( .IN1(n408), .IN2(n403), .S(add_sub_result_24_), .Q(N248) );
  NAND4X0 U680 ( .IN1(n504), .IN2(n493), .IN3(n497), .IN4(n495), .QN(N256) );
  INVX0 U681 ( .INP(n410), .ZN(n496) );
  NOR2X0 U682 ( .IN1(n496), .IN2(n411), .QN(n427) );
  NAND4X0 U683 ( .IN1(n504), .IN2(n491), .IN3(n497), .IN4(n499), .QN(N257) );
  NAND3X0 U684 ( .IN1(n412), .IN2(n500), .IN3(n482), .QN(n501) );
  NAND4X0 U685 ( .IN1(n504), .IN2(n493), .IN3(n501), .IN4(n491), .QN(N258) );
  NOR2X0 U686 ( .IN1(n815), .IN2(n495), .QN(N260) );
  INVX0 U687 ( .INP(n495), .ZN(n429) );
  AO22X1 U688 ( .IN1(n429), .IN2(n821), .IN3(n427), .IN4(n823), .Q(N261) );
  INVX0 U689 ( .INP(n497), .ZN(n428) );
  AO222X1 U690 ( .IN1(n823), .IN2(n428), .IN3(n821), .IN4(n427), .IN5(n801), 
        .IN6(n429), .Q(N262) );
  OA22X1 U691 ( .IN1(n807), .IN2(n497), .IN3(n815), .IN4(n501), .Q(n414) );
  OA22X1 U692 ( .IN1(n813), .IN2(n499), .IN3(n811), .IN4(n495), .Q(n413) );
  OA22X1 U693 ( .IN1(n791), .IN2(n495), .IN3(n811), .IN4(n499), .Q(n417) );
  OA22X1 U694 ( .IN1(n807), .IN2(n501), .IN3(n815), .IN4(n493), .Q(n416) );
  NAND3X0 U695 ( .IN1(n417), .IN2(n416), .IN3(n415), .QN(N264) );
  OA22X1 U696 ( .IN1(n781), .IN2(n495), .IN3(n811), .IN4(n497), .Q(n421) );
  OA22X1 U697 ( .IN1(n813), .IN2(n501), .IN3(n807), .IN4(n493), .Q(n420) );
  INVX0 U698 ( .INP(n491), .ZN(n422) );
  NAND4X0 U699 ( .IN1(n421), .IN2(n420), .IN3(n419), .IN4(n418), .QN(N265) );
  OA22X1 U700 ( .IN1(n791), .IN2(n497), .IN3(n811), .IN4(n501), .Q(n426) );
  OA22X1 U701 ( .IN1(n782), .IN2(n495), .IN3(n781), .IN4(n499), .Q(n425) );
  OA22X1 U702 ( .IN1(n813), .IN2(n493), .IN3(n815), .IN4(n504), .Q(n424) );
  NAND4X0 U703 ( .IN1(n426), .IN2(n425), .IN3(n424), .IN4(n423), .QN(N266) );
  NOR4X0 U704 ( .IN1(n429), .IN2(n428), .IN3(n427), .IN4(N258), .QN(n563) );
  OA22X1 U705 ( .IN1(n813), .IN2(n491), .IN3(n811), .IN4(n493), .Q(n433) );
  OA22X1 U706 ( .IN1(n774), .IN2(n495), .IN3(n781), .IN4(n497), .Q(n432) );
  OA22X1 U707 ( .IN1(n782), .IN2(n499), .IN3(n791), .IN4(n501), .Q(n431) );
  OA22X1 U708 ( .IN1(n807), .IN2(n504), .IN3(n815), .IN4(n839), .Q(n430) );
  NAND4X0 U709 ( .IN1(n433), .IN2(n432), .IN3(n431), .IN4(n430), .QN(N267) );
  OA22X1 U710 ( .IN1(n791), .IN2(n493), .IN3(n811), .IN4(n491), .Q(n437) );
  OA22X1 U711 ( .IN1(n766), .IN2(n495), .IN3(n782), .IN4(n497), .Q(n436) );
  OA22X1 U712 ( .IN1(n774), .IN2(n499), .IN3(n781), .IN4(n501), .Q(n435) );
  OA22X1 U713 ( .IN1(n813), .IN2(n504), .IN3(n807), .IN4(n839), .Q(n434) );
  NAND4X0 U714 ( .IN1(n437), .IN2(n436), .IN3(n435), .IN4(n434), .QN(N268) );
  OA22X1 U715 ( .IN1(n781), .IN2(n493), .IN3(n791), .IN4(n491), .Q(n441) );
  OA22X1 U716 ( .IN1(n758), .IN2(n495), .IN3(n774), .IN4(n497), .Q(n440) );
  OA22X1 U717 ( .IN1(n766), .IN2(n499), .IN3(n782), .IN4(n501), .Q(n439) );
  OA22X1 U718 ( .IN1(n813), .IN2(n839), .IN3(n811), .IN4(n504), .Q(n438) );
  NAND4X0 U719 ( .IN1(n441), .IN2(n440), .IN3(n439), .IN4(n438), .QN(N269) );
  OA22X1 U720 ( .IN1(n782), .IN2(n493), .IN3(n781), .IN4(n491), .Q(n445) );
  OA22X1 U721 ( .IN1(n766), .IN2(n497), .IN3(n750), .IN4(n495), .Q(n444) );
  OA22X1 U722 ( .IN1(n758), .IN2(n499), .IN3(n774), .IN4(n501), .Q(n443) );
  OA22X1 U723 ( .IN1(n791), .IN2(n504), .IN3(n811), .IN4(n839), .Q(n442) );
  NAND4X0 U724 ( .IN1(n445), .IN2(n444), .IN3(n443), .IN4(n442), .QN(N270) );
  OA22X1 U725 ( .IN1(n774), .IN2(n493), .IN3(n782), .IN4(n491), .Q(n449) );
  OA22X1 U726 ( .IN1(n742), .IN2(n495), .IN3(n758), .IN4(n497), .Q(n448) );
  OA22X1 U727 ( .IN1(n766), .IN2(n501), .IN3(n750), .IN4(n499), .Q(n447) );
  OA22X1 U728 ( .IN1(n781), .IN2(n504), .IN3(n791), .IN4(n839), .Q(n446) );
  NAND4X0 U729 ( .IN1(n449), .IN2(n448), .IN3(n447), .IN4(n446), .QN(N271) );
  OA22X1 U730 ( .IN1(n766), .IN2(n493), .IN3(n774), .IN4(n491), .Q(n454) );
  OA22X1 U731 ( .IN1(n734), .IN2(n495), .IN3(n750), .IN4(n497), .Q(n453) );
  OA22X1 U732 ( .IN1(n742), .IN2(n499), .IN3(n758), .IN4(n501), .Q(n452) );
  OA22X1 U733 ( .IN1(n782), .IN2(n504), .IN3(n781), .IN4(n839), .Q(n451) );
  NAND4X0 U734 ( .IN1(n454), .IN2(n453), .IN3(n452), .IN4(n451), .QN(N272) );
  OA22X1 U735 ( .IN1(n766), .IN2(n491), .IN3(n758), .IN4(n493), .Q(n459) );
  OA22X1 U736 ( .IN1(n742), .IN2(n497), .IN3(n723), .IN4(n495), .Q(n458) );
  OA22X1 U737 ( .IN1(n734), .IN2(n499), .IN3(n750), .IN4(n501), .Q(n457) );
  OA22X1 U738 ( .IN1(n774), .IN2(n504), .IN3(n782), .IN4(n839), .Q(n456) );
  NAND4X0 U739 ( .IN1(n459), .IN2(n458), .IN3(n457), .IN4(n456), .QN(N273) );
  OA22X1 U740 ( .IN1(n750), .IN2(n493), .IN3(n758), .IN4(n491), .Q(n463) );
  INVX0 U741 ( .INP(n509), .ZN(n503) );
  OA22X1 U742 ( .IN1(n503), .IN2(n495), .IN3(n734), .IN4(n497), .Q(n462) );
  OA22X1 U743 ( .IN1(n742), .IN2(n501), .IN3(n723), .IN4(n499), .Q(n461) );
  OA22X1 U744 ( .IN1(n766), .IN2(n504), .IN3(n774), .IN4(n839), .Q(n460) );
  NAND4X0 U745 ( .IN1(n463), .IN2(n462), .IN3(n461), .IN4(n460), .QN(N274) );
  OA22X1 U746 ( .IN1(n742), .IN2(n493), .IN3(n750), .IN4(n491), .Q(n468) );
  OA22X1 U747 ( .IN1(n565), .IN2(n495), .IN3(n723), .IN4(n497), .Q(n467) );
  OA22X1 U748 ( .IN1(n503), .IN2(n499), .IN3(n734), .IN4(n501), .Q(n466) );
  OA22X1 U749 ( .IN1(n766), .IN2(n839), .IN3(n758), .IN4(n504), .Q(n465) );
  NAND4X0 U750 ( .IN1(n468), .IN2(n467), .IN3(n466), .IN4(n465), .QN(N275) );
  OA22X1 U751 ( .IN1(n734), .IN2(n493), .IN3(n742), .IN4(n491), .Q(n472) );
  OA22X1 U752 ( .IN1(n503), .IN2(n497), .IN3(n492), .IN4(n495), .Q(n471) );
  OA22X1 U753 ( .IN1(n565), .IN2(n499), .IN3(n723), .IN4(n501), .Q(n470) );
  OA22X1 U754 ( .IN1(n750), .IN2(n504), .IN3(n758), .IN4(n839), .Q(n469) );
  NAND4X0 U755 ( .IN1(n472), .IN2(n471), .IN3(n470), .IN4(n469), .QN(N276) );
  OA22X1 U756 ( .IN1(n734), .IN2(n491), .IN3(n723), .IN4(n493), .Q(n477) );
  INVX0 U757 ( .INP(n473), .ZN(n494) );
  OA22X1 U758 ( .IN1(n565), .IN2(n497), .IN3(n494), .IN4(n495), .Q(n476) );
  OA22X1 U759 ( .IN1(n503), .IN2(n501), .IN3(n492), .IN4(n499), .Q(n475) );
  OA22X1 U760 ( .IN1(n742), .IN2(n504), .IN3(n750), .IN4(n839), .Q(n474) );
  NAND4X0 U761 ( .IN1(n477), .IN2(n476), .IN3(n475), .IN4(n474), .QN(N277) );
  OA22X1 U762 ( .IN1(n503), .IN2(n493), .IN3(n723), .IN4(n491), .Q(n481) );
  OA22X1 U763 ( .IN1(n502), .IN2(n495), .IN3(n492), .IN4(n497), .Q(n480) );
  OA22X1 U764 ( .IN1(n565), .IN2(n501), .IN3(n494), .IN4(n499), .Q(n479) );
  OA22X1 U765 ( .IN1(n734), .IN2(n504), .IN3(n742), .IN4(n839), .Q(n478) );
  NAND4X0 U766 ( .IN1(n481), .IN2(n480), .IN3(n479), .IN4(n478), .QN(N278) );
  OA22X1 U767 ( .IN1(n565), .IN2(n493), .IN3(n503), .IN4(n491), .Q(n486) );
  INVX0 U768 ( .INP(n482), .ZN(n498) );
  OA22X1 U769 ( .IN1(n494), .IN2(n497), .IN3(n498), .IN4(n495), .Q(n485) );
  OA22X1 U770 ( .IN1(n502), .IN2(n499), .IN3(n492), .IN4(n501), .Q(n484) );
  OA22X1 U771 ( .IN1(n734), .IN2(n839), .IN3(n723), .IN4(n504), .Q(n483) );
  NAND4X0 U772 ( .IN1(n486), .IN2(n485), .IN3(n484), .IN4(n483), .QN(N279) );
  OA22X1 U773 ( .IN1(n565), .IN2(n491), .IN3(n492), .IN4(n493), .Q(n490) );
  OA22X1 U774 ( .IN1(n502), .IN2(n497), .IN3(n500), .IN4(n495), .Q(n489) );
  OA22X1 U775 ( .IN1(n494), .IN2(n501), .IN3(n498), .IN4(n499), .Q(n488) );
  OA22X1 U776 ( .IN1(n503), .IN2(n504), .IN3(n723), .IN4(n839), .Q(n487) );
  NAND4X0 U777 ( .IN1(n490), .IN2(n489), .IN3(n488), .IN4(n487), .QN(N280) );
  OA22X1 U778 ( .IN1(n494), .IN2(n493), .IN3(n492), .IN4(n491), .Q(n508) );
  OA22X1 U779 ( .IN1(n498), .IN2(n497), .IN3(n496), .IN4(n495), .Q(n507) );
  OA22X1 U780 ( .IN1(n502), .IN2(n501), .IN3(n500), .IN4(n499), .Q(n506) );
  OA22X1 U781 ( .IN1(n565), .IN2(n504), .IN3(n503), .IN4(n839), .Q(n505) );
  NAND4X0 U782 ( .IN1(n508), .IN2(n507), .IN3(n506), .IN4(n505), .QN(N281) );
  NAND3X0 U783 ( .IN1(n509), .IN2(n522), .IN3(n565), .QN(n722) );
  AO22X1 U784 ( .IN1(n520), .IN2(add_result[12]), .IN3(n518), .IN4(
        sub_result[12]), .Q(n510) );
  INVX0 U785 ( .INP(n722), .ZN(n516) );
  NOR3X0 U786 ( .IN1(add_result[14]), .IN2(add_result[15]), .IN3(n14), .QN(
        n513) );
  NOR3X0 U787 ( .IN1(n511), .IN2(sub_result[14]), .IN3(sub_result[15]), .QN(
        n512) );
  AO22X1 U788 ( .IN1(n513), .IN2(add_result[13]), .IN3(n512), .IN4(
        sub_result[13]), .Q(n514) );
  NOR2X0 U789 ( .IN1(n516), .IN2(n515), .QN(N308) );
  INVX0 U790 ( .INP(add_result[12]), .ZN(n519) );
  INVX0 U791 ( .INP(sub_result[12]), .ZN(n517) );
  AO22X1 U792 ( .IN1(n520), .IN2(n519), .IN3(n518), .IN4(n517), .Q(n521) );
  NAND3X0 U793 ( .IN1(n522), .IN2(n729), .IN3(n521), .QN(n816) );
  NAND4X0 U794 ( .IN1(N308), .IN2(n816), .IN3(n799), .IN4(n790), .QN(n783) );
  NAND4X0 U795 ( .IN1(n799), .IN2(n722), .IN3(n728), .IN4(n783), .QN(N306) );
  NAND4X0 U796 ( .IN1(n790), .IN2(n721), .IN3(n728), .IN4(n783), .QN(N307) );
  AO22X1 U797 ( .IN1(exponent_factor_21[0]), .IN2(n825), .IN3(
        exponent_factor_12[0]), .IN4(n709), .Q(N34) );
  NAND3X0 U798 ( .IN1(n811), .IN2(n532), .IN3(n801), .QN(n545) );
  NAND3X0 U799 ( .IN1(n781), .IN2(n524), .IN3(n802), .QN(n540) );
  NAND3X0 U800 ( .IN1(n774), .IN2(n525), .IN3(n769), .QN(n541) );
  NAND3X0 U801 ( .IN1(n813), .IN2(n807), .IN3(n811), .QN(n523) );
  AND2X1 U802 ( .IN1(n540), .IN2(n542), .Q(n527) );
  NAND4X0 U803 ( .IN1(n529), .IN2(n527), .IN3(n541), .IN4(n543), .QN(n528) );
  NAND4X0 U804 ( .IN1(n545), .IN2(n540), .IN3(n541), .IN4(n528), .QN(N346) );
  NAND3X0 U805 ( .IN1(n527), .IN2(n544), .IN3(n528), .QN(N347) );
  NOR2X0 U806 ( .IN1(n815), .IN2(n543), .QN(N349) );
  AO22X1 U807 ( .IN1(exponent_factor_21[1]), .IN2(n825), .IN3(
        exponent_factor_12[1]), .IN4(n709), .Q(N35) );
  OAI22X1 U808 ( .IN1(n807), .IN2(n543), .IN3(n815), .IN4(n541), .QN(N350) );
  OAI222X1 U809 ( .IN1(n542), .IN2(n815), .IN3(n541), .IN4(n807), .IN5(n543), 
        .IN6(n813), .QN(N351) );
  OA22X1 U810 ( .IN1(n813), .IN2(n541), .IN3(n811), .IN4(n543), .Q(n531) );
  OA22X1 U811 ( .IN1(n807), .IN2(n542), .IN3(n815), .IN4(n540), .Q(n530) );
  OA22X1 U812 ( .IN1(n791), .IN2(n543), .IN3(n811), .IN4(n541), .Q(n535) );
  OA22X1 U813 ( .IN1(n813), .IN2(n542), .IN3(n807), .IN4(n540), .Q(n534) );
  AND2X1 U814 ( .IN1(n532), .IN2(n793), .Q(n546) );
  NAND3X0 U815 ( .IN1(n535), .IN2(n534), .IN3(n533), .QN(N353) );
  OA22X1 U816 ( .IN1(n781), .IN2(n543), .IN3(n791), .IN4(n541), .Q(n539) );
  OA22X1 U817 ( .IN1(n813), .IN2(n540), .IN3(n815), .IN4(n545), .Q(n538) );
  OR2X1 U818 ( .IN1(n542), .IN2(n811), .Q(n536) );
  NAND4X0 U819 ( .IN1(n539), .IN2(n538), .IN3(n537), .IN4(n536), .QN(N354) );
  OA22X1 U820 ( .IN1(n781), .IN2(n541), .IN3(n811), .IN4(n540), .Q(n550) );
  OA22X1 U821 ( .IN1(n782), .IN2(n543), .IN3(n791), .IN4(n542), .Q(n549) );
  OA22X1 U822 ( .IN1(n807), .IN2(n545), .IN3(n815), .IN4(n544), .Q(n548) );
  NAND4X0 U823 ( .IN1(n550), .IN2(n549), .IN3(n548), .IN4(n547), .QN(N355) );
  AO22X1 U824 ( .IN1(exponent_factor_21[2]), .IN2(n825), .IN3(
        exponent_factor_12[2]), .IN4(n709), .Q(N36) );
  AO22X1 U825 ( .IN1(exponent_factor_21[3]), .IN2(n825), .IN3(
        exponent_factor_12[3]), .IN4(n709), .Q(N37) );
  AO22X1 U826 ( .IN1(exponent_factor_21[4]), .IN2(n825), .IN3(
        exponent_factor_12[4]), .IN4(n709), .Q(N38) );
  OR4X1 U827 ( .IN1(input_factor_01[27]), .IN2(input_factor_01[30]), .IN3(
        input_factor_01[29]), .IN4(input_factor_01[23]), .Q(n551) );
  NOR4X0 U828 ( .IN1(input_factor_01[25]), .IN2(input_factor_01[24]), .IN3(
        n552), .IN4(n551), .QN(n561) );
  NOR4X0 U829 ( .IN1(input_factor_01[22]), .IN2(input_factor_01[21]), .IN3(
        input_factor_01[20]), .IN4(input_factor_01[19]), .QN(n560) );
  NOR4X0 U830 ( .IN1(input_factor_01[31]), .IN2(input_factor_01[18]), .IN3(
        input_factor_01[17]), .IN4(input_factor_01[16]), .QN(n559) );
  NAND4X0 U831 ( .IN1(n623), .IN2(n619), .IN3(n615), .IN4(n611), .QN(n557) );
  NAND4X0 U832 ( .IN1(n607), .IN2(n603), .IN3(n553), .IN4(n599), .QN(n556) );
  NAND4X0 U833 ( .IN1(n667), .IN2(n661), .IN3(n655), .IN4(n649), .QN(n555) );
  NAND4X0 U834 ( .IN1(n643), .IN2(n637), .IN3(n631), .IN4(n627), .QN(n554) );
  NOR4X0 U835 ( .IN1(n557), .IN2(n556), .IN3(n555), .IN4(n554), .QN(n558) );
  NAND3X0 U836 ( .IN1(n562), .IN2(n15), .IN3(n711), .QN(n571) );
  AOI22X1 U837 ( .IN1(input_factor_01[23]), .IN2(n8), .IN3(n716), .IN4(
        add_output_exponent_w1[0]), .QN(n575) );
  OA21X1 U838 ( .IN1(n565), .IN2(n564), .IN3(n563), .Q(n568) );
  INVX0 U839 ( .INP(n571), .ZN(n569) );
  INVX0 U840 ( .INP(n783), .ZN(n566) );
  OA21X1 U841 ( .IN1(n766), .IN2(n567), .IN3(n566), .Q(n572) );
  AOI22X1 U842 ( .IN1(n713), .IN2(add_output_exponent_w2[0]), .IN3(n715), 
        .IN4(add_output_exponent_w4[0]), .QN(n574) );
  NAND2X0 U843 ( .IN1(input_factor_02[23]), .IN2(n16), .QN(n581) );
  NAND4X0 U844 ( .IN1(n575), .IN2(n574), .IN3(n573), .IN4(n581), .QN(N380) );
  AOI22X1 U845 ( .IN1(input_factor_01[24]), .IN2(n8), .IN3(input_factor_02[24]), .IN4(n16), .QN(n579) );
  AOI22X1 U846 ( .IN1(n714), .IN2(add_output_exponent_w3[1]), .IN3(n713), 
        .IN4(add_output_exponent_w2[1]), .QN(n578) );
  NAND4X0 U847 ( .IN1(n579), .IN2(n578), .IN3(n577), .IN4(n576), .QN(N381) );
  AOI22X1 U848 ( .IN1(input_factor_01[25]), .IN2(n8), .IN3(n716), .IN4(
        add_output_exponent_w1[2]), .QN(n583) );
  AOI22X1 U849 ( .IN1(n714), .IN2(add_output_exponent_w3[2]), .IN3(n713), 
        .IN4(add_output_exponent_w2[2]), .QN(n582) );
  NAND4X0 U850 ( .IN1(n583), .IN2(n582), .IN3(n581), .IN4(n580), .QN(N382) );
  AOI22X1 U851 ( .IN1(input_factor_01[26]), .IN2(n8), .IN3(n716), .IN4(
        add_output_exponent_w1[3]), .QN(n586) );
  AOI22X1 U852 ( .IN1(n713), .IN2(add_output_exponent_w2[3]), .IN3(n715), 
        .IN4(add_output_exponent_w4[3]), .QN(n585) );
  NAND4X0 U853 ( .IN1(n586), .IN2(n585), .IN3(n584), .IN4(n594), .QN(N383) );
  AOI22X1 U854 ( .IN1(input_factor_01[27]), .IN2(n8), .IN3(n716), .IN4(
        add_output_exponent_w1[4]), .QN(n589) );
  AOI22X1 U855 ( .IN1(n713), .IN2(add_output_exponent_w2[4]), .IN3(n715), 
        .IN4(add_output_exponent_w4[4]), .QN(n588) );
  NAND4X0 U856 ( .IN1(n589), .IN2(n588), .IN3(n594), .IN4(n587), .QN(N384) );
  AOI22X1 U857 ( .IN1(input_factor_01[28]), .IN2(n8), .IN3(n716), .IN4(
        add_output_exponent_w1[5]), .QN(n592) );
  AOI22X1 U858 ( .IN1(n713), .IN2(add_output_exponent_w2[5]), .IN3(n715), 
        .IN4(add_output_exponent_w4[5]), .QN(n591) );
  NAND4X0 U859 ( .IN1(n592), .IN2(n591), .IN3(n594), .IN4(n590), .QN(N385) );
  AOI22X1 U860 ( .IN1(input_factor_01[29]), .IN2(n8), .IN3(n716), .IN4(
        add_output_exponent_w1[6]), .QN(n596) );
  AOI22X1 U861 ( .IN1(n714), .IN2(add_output_exponent_w3[6]), .IN3(n713), 
        .IN4(add_output_exponent_w2[6]), .QN(n595) );
  NAND4X0 U862 ( .IN1(n596), .IN2(n595), .IN3(n594), .IN4(n593), .QN(N386) );
  AO22X1 U864 ( .IN1(input_factor_01[30]), .IN2(n8), .IN3(n716), .IN4(
        add_output_exponent_w1[7]), .Q(n598) );
  AO22X1 U865 ( .IN1(n714), .IN2(add_output_exponent_w3[7]), .IN3(n713), .IN4(
        add_output_exponent_w2[7]), .Q(n597) );
  AO222X1 U866 ( .IN1(input_factor_02[0]), .IN2(n16), .IN3(n8), .IN4(
        input_factor_01[0]), .IN5(n716), .IN6(pre_sig_res_01[0]), .Q(N388) );
  AOI22X1 U867 ( .IN1(n713), .IN2(pre_sig_res_02[1]), .IN3(n716), .IN4(
        pre_sig_res_01[1]), .QN(n602) );
  OA22X1 U868 ( .IN1(n600), .IN2(n711), .IN3(n599), .IN4(n15), .Q(n601) );
  AO22X1 U869 ( .IN1(exponent_factor_21[5]), .IN2(n825), .IN3(
        exponent_factor_12[5]), .IN4(n709), .Q(N39) );
  AOI22X1 U870 ( .IN1(n713), .IN2(pre_sig_res_02[2]), .IN3(n716), .IN4(
        pre_sig_res_01[2]), .QN(n606) );
  OA22X1 U871 ( .IN1(n604), .IN2(n711), .IN3(n603), .IN4(n15), .Q(n605) );
  AOI22X1 U872 ( .IN1(n713), .IN2(pre_sig_res_02[3]), .IN3(n716), .IN4(
        pre_sig_res_01[3]), .QN(n610) );
  OA22X1 U873 ( .IN1(n608), .IN2(n711), .IN3(n607), .IN4(n15), .Q(n609) );
  AOI22X1 U874 ( .IN1(n713), .IN2(pre_sig_res_02[4]), .IN3(n716), .IN4(
        pre_sig_res_01[4]), .QN(n614) );
  OA22X1 U875 ( .IN1(n612), .IN2(n711), .IN3(n611), .IN4(n15), .Q(n613) );
  AOI22X1 U876 ( .IN1(n713), .IN2(pre_sig_res_02[5]), .IN3(n716), .IN4(
        pre_sig_res_01[5]), .QN(n618) );
  OA22X1 U877 ( .IN1(n616), .IN2(n711), .IN3(n615), .IN4(n15), .Q(n617) );
  AOI22X1 U878 ( .IN1(n713), .IN2(pre_sig_res_02[6]), .IN3(n716), .IN4(
        pre_sig_res_01[6]), .QN(n622) );
  OA22X1 U879 ( .IN1(n620), .IN2(n711), .IN3(n619), .IN4(n15), .Q(n621) );
  AOI22X1 U880 ( .IN1(n713), .IN2(pre_sig_res_02[7]), .IN3(n716), .IN4(
        pre_sig_res_01[7]), .QN(n626) );
  OA22X1 U881 ( .IN1(n624), .IN2(n711), .IN3(n623), .IN4(n15), .Q(n625) );
  AOI22X1 U882 ( .IN1(n713), .IN2(pre_sig_res_02[8]), .IN3(n716), .IN4(
        pre_sig_res_01[8]), .QN(n630) );
  OA22X1 U883 ( .IN1(n628), .IN2(n711), .IN3(n627), .IN4(n15), .Q(n629) );
  OA22X1 U884 ( .IN1(n632), .IN2(n711), .IN3(n631), .IN4(n15), .Q(n636) );
  NAND4X0 U885 ( .IN1(n636), .IN2(n635), .IN3(n634), .IN4(n633), .QN(N397) );
  OA22X1 U886 ( .IN1(n638), .IN2(n711), .IN3(n637), .IN4(n15), .Q(n642) );
  NAND4X0 U887 ( .IN1(n642), .IN2(n641), .IN3(n640), .IN4(n639), .QN(N398) );
  OA22X1 U888 ( .IN1(n644), .IN2(n711), .IN3(n643), .IN4(n15), .Q(n648) );
  NAND4X0 U889 ( .IN1(n648), .IN2(n647), .IN3(n646), .IN4(n645), .QN(N399) );
  AO22X1 U890 ( .IN1(exponent_factor_21[6]), .IN2(n825), .IN3(
        exponent_factor_12[6]), .IN4(n709), .Q(N40) );
  OA22X1 U891 ( .IN1(n650), .IN2(n711), .IN3(n649), .IN4(n15), .Q(n654) );
  NAND4X0 U892 ( .IN1(n654), .IN2(n653), .IN3(n652), .IN4(n651), .QN(N400) );
  OA22X1 U893 ( .IN1(n656), .IN2(n711), .IN3(n655), .IN4(n15), .Q(n660) );
  NAND4X0 U894 ( .IN1(n660), .IN2(n659), .IN3(n658), .IN4(n657), .QN(N401) );
  OA22X1 U895 ( .IN1(n662), .IN2(n711), .IN3(n661), .IN4(n15), .Q(n666) );
  NAND4X0 U896 ( .IN1(n666), .IN2(n665), .IN3(n664), .IN4(n663), .QN(N402) );
  OA22X1 U897 ( .IN1(n668), .IN2(n711), .IN3(n667), .IN4(n15), .Q(n672) );
  NAND4X0 U898 ( .IN1(n672), .IN2(n671), .IN3(n670), .IN4(n669), .QN(N403) );
  OA22X1 U899 ( .IN1(n674), .IN2(n711), .IN3(n673), .IN4(n15), .Q(n678) );
  AOI22X1 U900 ( .IN1(n714), .IN2(pre_sig_res_03[16]), .IN3(n713), .IN4(
        pre_sig_res_02[16]), .QN(n677) );
  NAND4X0 U901 ( .IN1(n678), .IN2(n677), .IN3(n676), .IN4(n675), .QN(N404) );
  OA22X1 U902 ( .IN1(n680), .IN2(n711), .IN3(n679), .IN4(n15), .Q(n684) );
  AOI22X1 U903 ( .IN1(n714), .IN2(pre_sig_res_03[17]), .IN3(n713), .IN4(
        pre_sig_res_02[17]), .QN(n683) );
  NAND4X0 U904 ( .IN1(n684), .IN2(n683), .IN3(n682), .IN4(n681), .QN(N405) );
  OA22X1 U905 ( .IN1(n686), .IN2(n711), .IN3(n685), .IN4(n15), .Q(n690) );
  AOI22X1 U906 ( .IN1(n714), .IN2(pre_sig_res_03[18]), .IN3(n713), .IN4(
        pre_sig_res_02[18]), .QN(n689) );
  NAND4X0 U907 ( .IN1(n690), .IN2(n689), .IN3(n688), .IN4(n687), .QN(N406) );
  OA22X1 U908 ( .IN1(n692), .IN2(n711), .IN3(n691), .IN4(n15), .Q(n696) );
  AOI22X1 U909 ( .IN1(n714), .IN2(pre_sig_res_03[19]), .IN3(n713), .IN4(
        pre_sig_res_02[19]), .QN(n695) );
  NAND4X0 U910 ( .IN1(n696), .IN2(n695), .IN3(n694), .IN4(n693), .QN(N407) );
  OA22X1 U911 ( .IN1(n698), .IN2(n711), .IN3(n697), .IN4(n15), .Q(n702) );
  AOI22X1 U912 ( .IN1(n714), .IN2(pre_sig_res_03[20]), .IN3(n713), .IN4(
        pre_sig_res_02[20]), .QN(n701) );
  NAND4X0 U913 ( .IN1(n702), .IN2(n701), .IN3(n700), .IN4(n699), .QN(N408) );
  OA22X1 U914 ( .IN1(n704), .IN2(n711), .IN3(n703), .IN4(n15), .Q(n708) );
  AOI22X1 U915 ( .IN1(n714), .IN2(pre_sig_res_03[21]), .IN3(n713), .IN4(
        pre_sig_res_02[21]), .QN(n707) );
  NAND4X0 U916 ( .IN1(n708), .IN2(n707), .IN3(n706), .IN4(n705), .QN(N409) );
  AO22X1 U917 ( .IN1(exponent_factor_21[7]), .IN2(n825), .IN3(
        exponent_factor_12[7]), .IN4(n709), .Q(N41) );
  OA22X1 U918 ( .IN1(n712), .IN2(n711), .IN3(n710), .IN4(n15), .Q(n720) );
  AOI22X1 U919 ( .IN1(n714), .IN2(pre_sig_res_03[22]), .IN3(n713), .IN4(
        pre_sig_res_02[22]), .QN(n719) );
  NAND4X0 U920 ( .IN1(n720), .IN2(n719), .IN3(n718), .IN4(n717), .QN(N410) );
  NOR2X0 U921 ( .IN1(n862), .IN2(n721), .QN(n822) );
  NOR2X0 U922 ( .IN1(n722), .IN2(n862), .QN(n824) );
  OA22X1 U923 ( .IN1(n734), .IN2(n812), .IN3(n723), .IN4(n810), .Q(n733) );
  OA22X1 U924 ( .IN1(n750), .IN2(n816), .IN3(n774), .IN4(n783), .Q(n727) );
  INVX0 U925 ( .INP(rst_n), .ZN(n826) );
  NAND3X0 U926 ( .IN1(n725), .IN2(n745), .IN3(n724), .QN(n726) );
  OA22X1 U927 ( .IN1(n862), .IN2(n727), .IN3(n826), .IN4(n726), .Q(n732) );
  NAND4X0 U928 ( .IN1(n733), .IN2(n732), .IN3(n731), .IN4(n730), .QN(n861) );
  OA22X1 U929 ( .IN1(n734), .IN2(n810), .IN3(n742), .IN4(n812), .Q(n741) );
  OA22X1 U930 ( .IN1(n774), .IN2(n790), .IN3(n782), .IN4(n783), .Q(n736) );
  OA22X1 U931 ( .IN1(n766), .IN2(n799), .IN3(n758), .IN4(n816), .Q(n735) );
  AO21X1 U932 ( .IN1(n736), .IN2(n735), .IN3(n862), .Q(n740) );
  NAND4X0 U933 ( .IN1(n741), .IN2(n740), .IN3(n739), .IN4(n738), .QN(n860) );
  OA22X1 U934 ( .IN1(n742), .IN2(n810), .IN3(n750), .IN4(n812), .Q(n749) );
  OA22X1 U935 ( .IN1(n782), .IN2(n790), .IN3(n781), .IN4(n783), .Q(n744) );
  OA22X1 U936 ( .IN1(n766), .IN2(n816), .IN3(n774), .IN4(n799), .Q(n743) );
  AO21X1 U937 ( .IN1(n744), .IN2(n743), .IN3(n862), .Q(n748) );
  NAND4X0 U938 ( .IN1(n749), .IN2(n748), .IN3(n747), .IN4(n746), .QN(n859) );
  OA22X1 U939 ( .IN1(n750), .IN2(n810), .IN3(n758), .IN4(n812), .Q(n757) );
  OA22X1 U940 ( .IN1(n781), .IN2(n790), .IN3(n791), .IN4(n783), .Q(n752) );
  OA22X1 U941 ( .IN1(n774), .IN2(n816), .IN3(n782), .IN4(n799), .Q(n751) );
  AO21X1 U942 ( .IN1(n752), .IN2(n751), .IN3(n862), .Q(n756) );
  NAND4X0 U943 ( .IN1(n757), .IN2(n756), .IN3(n755), .IN4(n754), .QN(n858) );
  OA22X1 U944 ( .IN1(n766), .IN2(n812), .IN3(n758), .IN4(n810), .Q(n765) );
  OA22X1 U945 ( .IN1(n791), .IN2(n790), .IN3(n811), .IN4(n783), .Q(n760) );
  OA22X1 U946 ( .IN1(n782), .IN2(n816), .IN3(n781), .IN4(n799), .Q(n759) );
  AO21X1 U947 ( .IN1(n760), .IN2(n759), .IN3(n862), .Q(n764) );
  NAND4X0 U948 ( .IN1(n765), .IN2(n764), .IN3(n763), .IN4(n762), .QN(n857) );
  OA22X1 U949 ( .IN1(n766), .IN2(n810), .IN3(n774), .IN4(n812), .Q(n773) );
  OA22X1 U950 ( .IN1(n813), .IN2(n783), .IN3(n811), .IN4(n790), .Q(n768) );
  OA22X1 U951 ( .IN1(n781), .IN2(n816), .IN3(n791), .IN4(n799), .Q(n767) );
  AO21X1 U952 ( .IN1(n768), .IN2(n767), .IN3(n862), .Q(n772) );
  NAND4X0 U953 ( .IN1(n773), .IN2(n772), .IN3(n771), .IN4(n770), .QN(n856) );
  OA22X1 U954 ( .IN1(n774), .IN2(n810), .IN3(n782), .IN4(n812), .Q(n780) );
  OA22X1 U955 ( .IN1(n813), .IN2(n790), .IN3(n807), .IN4(n783), .Q(n776) );
  OA22X1 U956 ( .IN1(n791), .IN2(n816), .IN3(n811), .IN4(n799), .Q(n775) );
  AO21X1 U957 ( .IN1(n776), .IN2(n775), .IN3(n862), .Q(n779) );
  NAND4X0 U958 ( .IN1(n780), .IN2(n779), .IN3(n778), .IN4(n777), .QN(n855) );
  OA22X1 U959 ( .IN1(n782), .IN2(n810), .IN3(n781), .IN4(n812), .Q(n789) );
  OA22X1 U960 ( .IN1(n807), .IN2(n790), .IN3(n815), .IN4(n783), .Q(n785) );
  OA22X1 U961 ( .IN1(n813), .IN2(n799), .IN3(n811), .IN4(n816), .Q(n784) );
  AO21X1 U962 ( .IN1(n785), .IN2(n784), .IN3(n862), .Q(n788) );
  NAND4X0 U963 ( .IN1(n789), .IN2(n788), .IN3(n787), .IN4(n786), .QN(n854) );
  OA222X1 U964 ( .IN1(n816), .IN2(n813), .IN3(n790), .IN4(n815), .IN5(n799), 
        .IN6(n807), .Q(n792) );
  OA22X1 U965 ( .IN1(n862), .IN2(n792), .IN3(n791), .IN4(n812), .Q(n798) );
  NAND4X0 U966 ( .IN1(n798), .IN2(n797), .IN3(n796), .IN4(n795), .QN(n853) );
  OA22X1 U967 ( .IN1(n807), .IN2(n816), .IN3(n815), .IN4(n799), .Q(n800) );
  OA22X1 U968 ( .IN1(n811), .IN2(n812), .IN3(n800), .IN4(n826), .Q(n806) );
  NAND4X0 U969 ( .IN1(n806), .IN2(n805), .IN3(n804), .IN4(n803), .QN(n852) );
  AOI22X1 U970 ( .IN1(pre_sig_res_03[11]), .IN2(n826), .IN3(n814), .IN4(n823), 
        .QN(n809) );
  OA22X1 U971 ( .IN1(n813), .IN2(n810), .IN3(n807), .IN4(n812), .Q(n808) );
  OA22X1 U972 ( .IN1(n813), .IN2(n812), .IN3(n811), .IN4(n810), .Q(n820) );
  OR3X1 U973 ( .IN1(n816), .IN2(n826), .IN3(n815), .Q(n818) );
  NAND4X0 U974 ( .IN1(n820), .IN2(n819), .IN3(n818), .IN4(n817), .QN(n850) );
  AO222X1 U975 ( .IN1(n823), .IN2(n822), .IN3(n821), .IN4(n824), .IN5(n826), 
        .IN6(pre_sig_res_03[10]), .Q(n849) );
  AO22X1 U976 ( .IN1(pre_sig_res_03[9]), .IN2(n826), .IN3(n824), .IN4(n823), 
        .Q(n848) );
  NOR2X0 U977 ( .IN1(n825), .IN2(n862), .QN(n835) );
  AOI22X1 U978 ( .IN1(input_factor_01[23]), .IN2(n835), .IN3(n862), .IN4(
        larger_exponent[0]), .QN(n828) );
  NOR2X0 U979 ( .IN1(n827), .IN2(n826), .QN(n831) );
  NAND2X0 U980 ( .IN1(input_factor_02[23]), .IN2(n831), .QN(n829) );
  AO222X1 U981 ( .IN1(input_factor_01[24]), .IN2(n835), .IN3(n862), .IN4(
        larger_exponent[1]), .IN5(input_factor_02[24]), .IN6(n831), .Q(n846)
         );
  AOI22X1 U982 ( .IN1(input_factor_01[25]), .IN2(n835), .IN3(n862), .IN4(
        larger_exponent[2]), .QN(n830) );
  AOI22X1 U983 ( .IN1(input_factor_01[26]), .IN2(n835), .IN3(n862), .IN4(
        larger_exponent[3]), .QN(n832) );
  AOI22X1 U984 ( .IN1(input_factor_01[27]), .IN2(n835), .IN3(n862), .IN4(
        larger_exponent[4]), .QN(n833) );
  AOI22X1 U985 ( .IN1(input_factor_01[28]), .IN2(n835), .IN3(n862), .IN4(
        larger_exponent[5]), .QN(n834) );
  AOI22X1 U986 ( .IN1(input_factor_01[29]), .IN2(n835), .IN3(n862), .IN4(
        larger_exponent[6]), .QN(n837) );
endmodule


module add_145 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_146 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_147 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_148 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_149 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_150 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_151 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_152 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_153 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_154 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_155 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_156 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_157 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_158 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_159 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_160 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_161 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_162 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_163 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_164 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_165 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_166 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_167 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_168 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(b), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(b), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module adder24_3 ( clk, rst_n, a, b, cin, out );
  input [23:0] a;
  input [23:0] b;
  output [24:0] out;
  input clk, rst_n, cin;
  wire   c_tmp;
  wire   [24:0] s;
  wire   [22:0] c;

  add_168 add_01 ( .s(s[0]), .a(a[0]), .b(b[0]), .ci(1'b0), .co(c[0]) );
  add_167 add_02 ( .s(s[1]), .a(a[1]), .b(b[1]), .ci(c[0]), .co(c[1]) );
  add_166 add_03 ( .s(s[2]), .a(a[2]), .b(b[2]), .ci(c[1]), .co(c[2]) );
  add_165 add_04 ( .s(s[3]), .a(a[3]), .b(b[3]), .ci(c[2]), .co(c[3]) );
  add_164 add_05 ( .s(s[4]), .a(a[4]), .b(b[4]), .ci(c[3]), .co(c[4]) );
  add_163 add_06 ( .s(s[5]), .a(a[5]), .b(b[5]), .ci(c[4]), .co(c[5]) );
  add_162 add_07 ( .s(s[6]), .a(a[6]), .b(b[6]), .ci(c[5]), .co(c[6]) );
  add_161 add_08 ( .s(s[7]), .a(a[7]), .b(b[7]), .ci(c[6]), .co(c[7]) );
  add_160 add_09 ( .s(s[8]), .a(a[8]), .b(b[8]), .ci(c[7]), .co(c[8]) );
  add_159 add_10 ( .s(s[9]), .a(a[9]), .b(b[9]), .ci(c[8]), .co(c[9]) );
  add_158 add_11 ( .s(s[10]), .a(a[10]), .b(b[10]), .ci(c[9]), .co(c[10]) );
  add_157 add_12 ( .s(s[11]), .a(a[11]), .b(b[11]), .ci(c_tmp), .co(c[11]) );
  add_156 add_13 ( .s(s[12]), .a(a[12]), .b(b[12]), .ci(c[11]), .co(c[12]) );
  add_155 add_14 ( .s(s[13]), .a(a[13]), .b(b[13]), .ci(c[12]), .co(c[13]) );
  add_154 add_15 ( .s(s[14]), .a(a[14]), .b(b[14]), .ci(c[13]), .co(c[14]) );
  add_153 add_16 ( .s(s[15]), .a(a[15]), .b(b[15]), .ci(c[14]), .co(c[15]) );
  add_152 add_17 ( .s(s[16]), .a(a[16]), .b(b[16]), .ci(c[15]), .co(c[16]) );
  add_151 add_18 ( .s(s[17]), .a(a[17]), .b(b[17]), .ci(c[16]), .co(c[17]) );
  add_150 add_19 ( .s(s[18]), .a(a[18]), .b(b[18]), .ci(c[17]), .co(c[18]) );
  add_149 add_20 ( .s(s[19]), .a(a[19]), .b(b[19]), .ci(c[18]), .co(c[19]) );
  add_148 add_21 ( .s(s[20]), .a(a[20]), .b(b[20]), .ci(c[19]), .co(c[20]) );
  add_147 add_22 ( .s(s[21]), .a(a[21]), .b(b[21]), .ci(c[20]), .co(c[21]) );
  add_146 add_23 ( .s(s[22]), .a(a[22]), .b(b[22]), .ci(c[21]), .co(c[22]) );
  add_145 add_24 ( .s(s[23]), .a(a[23]), .b(b[23]), .ci(c[22]), .co(s[24]) );
  DFFARX1 out_reg_10_ ( .D(s[10]), .CLK(clk), .RSTB(rst_n), .Q(out[10]) );
  DFFARX1 out_reg_9_ ( .D(s[9]), .CLK(clk), .RSTB(rst_n), .Q(out[9]) );
  DFFARX1 out_reg_8_ ( .D(s[8]), .CLK(clk), .RSTB(rst_n), .Q(out[8]) );
  DFFARX1 out_reg_7_ ( .D(s[7]), .CLK(clk), .RSTB(rst_n), .Q(out[7]) );
  DFFARX1 out_reg_6_ ( .D(s[6]), .CLK(clk), .RSTB(rst_n), .Q(out[6]) );
  DFFARX1 out_reg_5_ ( .D(s[5]), .CLK(clk), .RSTB(rst_n), .Q(out[5]) );
  DFFARX1 out_reg_4_ ( .D(s[4]), .CLK(clk), .RSTB(rst_n), .Q(out[4]) );
  DFFARX1 out_reg_3_ ( .D(s[3]), .CLK(clk), .RSTB(rst_n), .Q(out[3]) );
  DFFARX1 out_reg_2_ ( .D(s[2]), .CLK(clk), .RSTB(rst_n), .Q(out[2]) );
  DFFARX1 out_reg_1_ ( .D(s[1]), .CLK(clk), .RSTB(rst_n), .Q(out[1]) );
  DFFARX1 out_reg_0_ ( .D(s[0]), .CLK(clk), .RSTB(rst_n), .Q(out[0]) );
  DFFARX1 c_tmp_reg ( .D(c[10]), .CLK(clk), .RSTB(rst_n), .Q(c_tmp) );
  DFFARX1 out_reg_24_ ( .D(s[24]), .CLK(clk), .RSTB(rst_n), .Q(out[24]) );
  DFFARX1 out_reg_23_ ( .D(s[23]), .CLK(clk), .RSTB(rst_n), .Q(out[23]) );
  DFFARX1 out_reg_22_ ( .D(s[22]), .CLK(clk), .RSTB(rst_n), .Q(out[22]) );
  DFFARX1 out_reg_21_ ( .D(s[21]), .CLK(clk), .RSTB(rst_n), .Q(out[21]) );
  DFFARX1 out_reg_20_ ( .D(s[20]), .CLK(clk), .RSTB(rst_n), .Q(out[20]) );
  DFFARX1 out_reg_19_ ( .D(s[19]), .CLK(clk), .RSTB(rst_n), .Q(out[19]) );
  DFFARX1 out_reg_18_ ( .D(s[18]), .CLK(clk), .RSTB(rst_n), .Q(out[18]) );
  DFFARX1 out_reg_17_ ( .D(s[17]), .CLK(clk), .RSTB(rst_n), .Q(out[17]) );
  DFFARX1 out_reg_16_ ( .D(s[16]), .CLK(clk), .RSTB(rst_n), .Q(out[16]) );
  DFFARX1 out_reg_15_ ( .D(s[15]), .CLK(clk), .RSTB(rst_n), .Q(out[15]) );
  DFFARX1 out_reg_14_ ( .D(s[14]), .CLK(clk), .RSTB(rst_n), .Q(out[14]) );
  DFFARX1 out_reg_13_ ( .D(s[13]), .CLK(clk), .RSTB(rst_n), .Q(out[13]) );
  DFFARX1 out_reg_12_ ( .D(s[12]), .CLK(clk), .RSTB(rst_n), .Q(out[12]) );
  DFFARX1 out_reg_11_ ( .D(s[11]), .CLK(clk), .RSTB(rst_n), .Q(out[11]) );
endmodule


module add_169 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_170 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_171 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_172 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_173 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_174 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_175 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_176 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_177 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_178 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_179 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_180 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_181 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_182 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_183 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_184 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_185 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_186 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_187 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_188 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_189 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_190 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_191 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_192 ( s, a, ci, co, b_BAR );
  input a, ci, b_BAR;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(b_BAR), .IN2(n1), .QN(co) );
  INVX0 U2 ( .INP(a), .ZN(n1) );
  MUX21X1 U3 ( .IN1(a), .IN2(n1), .S(b_BAR), .Q(s) );
endmodule


module adder24_4 ( clk, rst_n, a, b, cin, out );
  input [23:0] a;
  input [23:0] b;
  output [24:0] out;
  input clk, rst_n, cin;
  wire   c_tmp, n_1_net_, n_2_net_, n_3_net_, n_4_net_, n_5_net_, n_6_net_,
         n_7_net_, n_8_net_, n_9_net_, n_10_net_, n_11_net_, n_12_net_,
         n_13_net_, n_14_net_, n_15_net_, n_16_net_, n_17_net_, n_18_net_,
         n_19_net_, n_20_net_, n_21_net_, n_22_net_, n_23_net_;
  wire   [24:0] s;
  wire   [23:0] c;

  add_192 add_01 ( .s(s[0]), .a(a[0]), .ci(1'b1), .co(c[0]), .b_BAR(b[0]) );
  add_191 add_02 ( .s(s[1]), .a(a[1]), .b(n_1_net_), .ci(c[0]), .co(c[1]) );
  add_190 add_03 ( .s(s[2]), .a(a[2]), .b(n_2_net_), .ci(c[1]), .co(c[2]) );
  add_189 add_04 ( .s(s[3]), .a(a[3]), .b(n_3_net_), .ci(c[2]), .co(c[3]) );
  add_188 add_05 ( .s(s[4]), .a(a[4]), .b(n_4_net_), .ci(c[3]), .co(c[4]) );
  add_187 add_06 ( .s(s[5]), .a(a[5]), .b(n_5_net_), .ci(c[4]), .co(c[5]) );
  add_186 add_07 ( .s(s[6]), .a(a[6]), .b(n_6_net_), .ci(c[5]), .co(c[6]) );
  add_185 add_08 ( .s(s[7]), .a(a[7]), .b(n_7_net_), .ci(c[6]), .co(c[7]) );
  add_184 add_09 ( .s(s[8]), .a(a[8]), .b(n_8_net_), .ci(c[7]), .co(c[8]) );
  add_183 add_10 ( .s(s[9]), .a(a[9]), .b(n_9_net_), .ci(c[8]), .co(c[9]) );
  add_182 add_11 ( .s(s[10]), .a(a[10]), .b(n_10_net_), .ci(c[9]), .co(c[10])
         );
  add_181 add_12 ( .s(s[11]), .a(a[11]), .b(n_11_net_), .ci(c_tmp), .co(c[11])
         );
  add_180 add_13 ( .s(s[12]), .a(a[12]), .b(n_12_net_), .ci(c[11]), .co(c[12])
         );
  add_179 add_14 ( .s(s[13]), .a(a[13]), .b(n_13_net_), .ci(c[12]), .co(c[13])
         );
  add_178 add_15 ( .s(s[14]), .a(a[14]), .b(n_14_net_), .ci(c[13]), .co(c[14])
         );
  add_177 add_16 ( .s(s[15]), .a(a[15]), .b(n_15_net_), .ci(c[14]), .co(c[15])
         );
  add_176 add_17 ( .s(s[16]), .a(a[16]), .b(n_16_net_), .ci(c[15]), .co(c[16])
         );
  add_175 add_18 ( .s(s[17]), .a(a[17]), .b(n_17_net_), .ci(c[16]), .co(c[17])
         );
  add_174 add_19 ( .s(s[18]), .a(a[18]), .b(n_18_net_), .ci(c[17]), .co(c[18])
         );
  add_173 add_20 ( .s(s[19]), .a(a[19]), .b(n_19_net_), .ci(c[18]), .co(c[19])
         );
  add_172 add_21 ( .s(s[20]), .a(a[20]), .b(n_20_net_), .ci(c[19]), .co(c[20])
         );
  add_171 add_22 ( .s(s[21]), .a(a[21]), .b(n_21_net_), .ci(c[20]), .co(c[21])
         );
  add_170 add_23 ( .s(s[22]), .a(a[22]), .b(n_22_net_), .ci(c[21]), .co(c[22])
         );
  add_169 add_24 ( .s(s[23]), .a(a[23]), .b(n_23_net_), .ci(c[22]), .co(c[23])
         );
  DFFARX1 out_reg_10_ ( .D(s[10]), .CLK(clk), .RSTB(rst_n), .Q(out[10]) );
  DFFARX1 out_reg_9_ ( .D(s[9]), .CLK(clk), .RSTB(rst_n), .Q(out[9]) );
  DFFARX1 out_reg_8_ ( .D(s[8]), .CLK(clk), .RSTB(rst_n), .Q(out[8]) );
  DFFARX1 out_reg_7_ ( .D(s[7]), .CLK(clk), .RSTB(rst_n), .Q(out[7]) );
  DFFARX1 out_reg_6_ ( .D(s[6]), .CLK(clk), .RSTB(rst_n), .Q(out[6]) );
  DFFARX1 out_reg_5_ ( .D(s[5]), .CLK(clk), .RSTB(rst_n), .Q(out[5]) );
  DFFARX1 out_reg_4_ ( .D(s[4]), .CLK(clk), .RSTB(rst_n), .Q(out[4]) );
  DFFARX1 out_reg_3_ ( .D(s[3]), .CLK(clk), .RSTB(rst_n), .Q(out[3]) );
  DFFARX1 out_reg_2_ ( .D(s[2]), .CLK(clk), .RSTB(rst_n), .Q(out[2]) );
  DFFARX1 out_reg_1_ ( .D(s[1]), .CLK(clk), .RSTB(rst_n), .Q(out[1]) );
  DFFARX1 out_reg_0_ ( .D(s[0]), .CLK(clk), .RSTB(rst_n), .Q(out[0]) );
  DFFARX1 c_tmp_reg ( .D(c[10]), .CLK(clk), .RSTB(rst_n), .Q(c_tmp) );
  DFFARX1 out_reg_24_ ( .D(s[24]), .CLK(clk), .RSTB(rst_n), .Q(out[24]) );
  DFFARX1 out_reg_23_ ( .D(s[23]), .CLK(clk), .RSTB(rst_n), .Q(out[23]) );
  DFFARX1 out_reg_22_ ( .D(s[22]), .CLK(clk), .RSTB(rst_n), .Q(out[22]) );
  DFFARX1 out_reg_21_ ( .D(s[21]), .CLK(clk), .RSTB(rst_n), .Q(out[21]) );
  DFFARX1 out_reg_20_ ( .D(s[20]), .CLK(clk), .RSTB(rst_n), .Q(out[20]) );
  DFFARX1 out_reg_19_ ( .D(s[19]), .CLK(clk), .RSTB(rst_n), .Q(out[19]) );
  DFFARX1 out_reg_18_ ( .D(s[18]), .CLK(clk), .RSTB(rst_n), .Q(out[18]) );
  DFFARX1 out_reg_17_ ( .D(s[17]), .CLK(clk), .RSTB(rst_n), .Q(out[17]) );
  DFFARX1 out_reg_16_ ( .D(s[16]), .CLK(clk), .RSTB(rst_n), .Q(out[16]) );
  DFFARX1 out_reg_15_ ( .D(s[15]), .CLK(clk), .RSTB(rst_n), .Q(out[15]) );
  DFFARX1 out_reg_14_ ( .D(s[14]), .CLK(clk), .RSTB(rst_n), .Q(out[14]) );
  DFFARX1 out_reg_13_ ( .D(s[13]), .CLK(clk), .RSTB(rst_n), .Q(out[13]) );
  DFFARX1 out_reg_12_ ( .D(s[12]), .CLK(clk), .RSTB(rst_n), .Q(out[12]) );
  DFFARX1 out_reg_11_ ( .D(s[11]), .CLK(clk), .RSTB(rst_n), .Q(out[11]) );
  INVX0 U3 ( .INP(b[1]), .ZN(n_1_net_) );
  INVX0 U4 ( .INP(b[2]), .ZN(n_2_net_) );
  INVX0 U5 ( .INP(b[3]), .ZN(n_3_net_) );
  INVX0 U6 ( .INP(b[4]), .ZN(n_4_net_) );
  INVX0 U7 ( .INP(b[5]), .ZN(n_5_net_) );
  INVX0 U8 ( .INP(b[6]), .ZN(n_6_net_) );
  INVX0 U9 ( .INP(b[7]), .ZN(n_7_net_) );
  INVX0 U10 ( .INP(b[8]), .ZN(n_8_net_) );
  INVX0 U11 ( .INP(b[9]), .ZN(n_9_net_) );
  INVX0 U12 ( .INP(b[10]), .ZN(n_10_net_) );
  INVX0 U13 ( .INP(c[23]), .ZN(s[24]) );
  INVX0 U14 ( .INP(b[11]), .ZN(n_11_net_) );
  INVX0 U15 ( .INP(b[12]), .ZN(n_12_net_) );
  INVX0 U16 ( .INP(b[13]), .ZN(n_13_net_) );
  INVX0 U17 ( .INP(b[14]), .ZN(n_14_net_) );
  INVX0 U18 ( .INP(b[15]), .ZN(n_15_net_) );
  INVX0 U19 ( .INP(b[16]), .ZN(n_16_net_) );
  INVX0 U20 ( .INP(b[17]), .ZN(n_17_net_) );
  INVX0 U21 ( .INP(b[18]), .ZN(n_18_net_) );
  INVX0 U22 ( .INP(b[19]), .ZN(n_19_net_) );
  INVX0 U23 ( .INP(b[20]), .ZN(n_20_net_) );
  INVX0 U24 ( .INP(b[21]), .ZN(n_21_net_) );
  INVX0 U25 ( .INP(b[22]), .ZN(n_22_net_) );
  INVX0 U26 ( .INP(b[23]), .ZN(n_23_net_) );
endmodule


module add_113 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  XNOR2X1 U1 ( .IN1(ci), .IN2(a), .Q(s) );
endmodule


module add_114 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_115 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_116 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_117 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_118 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_119 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_120 ( s, a, ci, co, b_BAR );
  input a, ci, b_BAR;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(b_BAR), .IN2(n1), .QN(co) );
  INVX0 U2 ( .INP(a), .ZN(n1) );
  MUX21X1 U3 ( .IN1(a), .IN2(n1), .S(b_BAR), .Q(s) );
endmodule


module adder8_9 ( out, a, b, cin );
  output [7:0] out;
  input [7:0] a;
  input [7:0] b;
  input cin;
  wire   n_1_net_, n_2_net_, n_4_net_;
  wire   [6:0] c;

  add_120 add_01 ( .s(out[0]), .a(a[0]), .ci(1'b1), .co(c[0]), .b_BAR(b[0]) );
  add_119 add_02 ( .s(out[1]), .a(a[1]), .b(n_1_net_), .ci(c[0]), .co(c[1]) );
  add_118 add_03 ( .s(out[2]), .a(a[2]), .b(n_2_net_), .ci(c[1]), .co(c[2]) );
  add_117 add_04 ( .s(out[3]), .a(a[3]), .b(1'b1), .ci(c[2]), .co(c[3]) );
  add_116 add_05 ( .s(out[4]), .a(a[4]), .b(n_4_net_), .ci(c[3]), .co(c[4]) );
  add_115 add_06 ( .s(out[5]), .a(a[5]), .b(1'b1), .ci(c[4]), .co(c[5]) );
  add_114 add_07 ( .s(out[6]), .a(a[6]), .b(1'b1), .ci(c[5]), .co(c[6]) );
  add_113 add_08 ( .s(out[7]), .a(a[7]), .b(1'b1), .ci(c[6]) );
  INVX0 U1 ( .INP(b[1]), .ZN(n_1_net_) );
  INVX0 U2 ( .INP(b[2]), .ZN(n_2_net_) );
  INVX0 U3 ( .INP(b[4]), .ZN(n_4_net_) );
endmodule


module add_121 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  XNOR2X1 U1 ( .IN1(ci), .IN2(a), .Q(s) );
endmodule


module add_122 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_123 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_124 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_125 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_126 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_127 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_128 ( s, a, ci, co, b_BAR );
  input a, ci, b_BAR;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(b_BAR), .IN2(n1), .QN(co) );
  INVX0 U2 ( .INP(a), .ZN(n1) );
  MUX21X1 U3 ( .IN1(a), .IN2(n1), .S(b_BAR), .Q(s) );
endmodule


module adder8_10 ( out, a, b, cin );
  output [7:0] out;
  input [7:0] a;
  input [7:0] b;
  input cin;
  wire   n_1_net_, n_2_net_, n_3_net_;
  wire   [6:0] c;

  add_128 add_01 ( .s(out[0]), .a(a[0]), .ci(1'b1), .co(c[0]), .b_BAR(b[0]) );
  add_127 add_02 ( .s(out[1]), .a(a[1]), .b(n_1_net_), .ci(c[0]), .co(c[1]) );
  add_126 add_03 ( .s(out[2]), .a(a[2]), .b(n_2_net_), .ci(c[1]), .co(c[2]) );
  add_125 add_04 ( .s(out[3]), .a(a[3]), .b(n_3_net_), .ci(c[2]), .co(c[3]) );
  add_124 add_05 ( .s(out[4]), .a(a[4]), .b(1'b1), .ci(c[3]), .co(c[4]) );
  add_123 add_06 ( .s(out[5]), .a(a[5]), .b(1'b1), .ci(c[4]), .co(c[5]) );
  add_122 add_07 ( .s(out[6]), .a(a[6]), .b(1'b1), .ci(c[5]), .co(c[6]) );
  add_121 add_08 ( .s(out[7]), .a(a[7]), .b(1'b1), .ci(c[6]) );
  INVX0 U1 ( .INP(b[1]), .ZN(n_1_net_) );
  INVX0 U2 ( .INP(b[2]), .ZN(n_2_net_) );
  INVX0 U3 ( .INP(b[3]), .ZN(n_3_net_) );
endmodule


module add_129 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  XNOR2X1 U1 ( .IN1(ci), .IN2(a), .Q(s) );
endmodule


module add_130 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_131 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_132 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_133 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_134 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_135 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_136 ( s, a, ci, co, b_BAR );
  input a, ci, b_BAR;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(b_BAR), .IN2(n1), .QN(co) );
  INVX0 U2 ( .INP(a), .ZN(n1) );
  MUX21X1 U3 ( .IN1(a), .IN2(n1), .S(b_BAR), .Q(s) );
endmodule


module adder8_11 ( out, a, b, cin );
  output [7:0] out;
  input [7:0] a;
  input [7:0] b;
  input cin;
  wire   n_1_net_, n_2_net_, n_3_net_;
  wire   [6:0] c;

  add_136 add_01 ( .s(out[0]), .a(a[0]), .ci(1'b1), .co(c[0]), .b_BAR(b[0]) );
  add_135 add_02 ( .s(out[1]), .a(a[1]), .b(n_1_net_), .ci(c[0]), .co(c[1]) );
  add_134 add_03 ( .s(out[2]), .a(a[2]), .b(n_2_net_), .ci(c[1]), .co(c[2]) );
  add_133 add_04 ( .s(out[3]), .a(a[3]), .b(n_3_net_), .ci(c[2]), .co(c[3]) );
  add_132 add_05 ( .s(out[4]), .a(a[4]), .b(1'b1), .ci(c[3]), .co(c[4]) );
  add_131 add_06 ( .s(out[5]), .a(a[5]), .b(1'b1), .ci(c[4]), .co(c[5]) );
  add_130 add_07 ( .s(out[6]), .a(a[6]), .b(1'b1), .ci(c[5]), .co(c[6]) );
  add_129 add_08 ( .s(out[7]), .a(a[7]), .b(1'b1), .ci(c[6]) );
  INVX0 U1 ( .INP(b[1]), .ZN(n_1_net_) );
  INVX0 U2 ( .INP(b[2]), .ZN(n_2_net_) );
  INVX0 U3 ( .INP(b[3]), .ZN(n_3_net_) );
endmodule


module add_137 ( s, a, b, co, ci_BAR );
  input a, b, ci_BAR;
  output s, co;


  XNOR2X1 U1 ( .IN1(a), .IN2(ci_BAR), .Q(s) );
endmodule


module add_138 ( s, a, b, ci, co_BAR );
  input a, b, ci;
  output s, co_BAR;


  NAND2X0 U1 ( .IN1(ci), .IN2(a), .QN(co_BAR) );
  OA21X1 U2 ( .IN1(ci), .IN2(a), .IN3(co_BAR), .Q(s) );
endmodule


module add_139 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_140 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_141 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_142 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_143 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_144 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(b), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(b), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module adder8_12 ( out, a, b, cin );
  output [7:0] out;
  input [7:0] a;
  input [7:0] b;
  input cin;

  wire   [6:0] c;

  add_144 add_01 ( .s(out[0]), .a(a[0]), .b(b[0]), .ci(1'b0), .co(c[0]) );
  add_143 add_02 ( .s(out[1]), .a(a[1]), .b(1'b0), .ci(c[0]), .co(c[1]) );
  add_142 add_03 ( .s(out[2]), .a(a[2]), .b(1'b0), .ci(c[1]), .co(c[2]) );
  add_141 add_04 ( .s(out[3]), .a(a[3]), .b(1'b0), .ci(c[2]), .co(c[3]) );
  add_140 add_05 ( .s(out[4]), .a(a[4]), .b(1'b0), .ci(c[3]), .co(c[4]) );
  add_139 add_06 ( .s(out[5]), .a(a[5]), .b(1'b0), .ci(c[4]), .co(c[5]) );
  add_138 add_07 ( .s(out[6]), .a(a[6]), .b(1'b0), .ci(c[5]), .co_BAR(c[6]) );
  add_137 add_08 ( .s(out[7]), .a(a[7]), .b(1'b0), .ci_BAR(c[6]) );
endmodule


module add_193 ( s, a, ci, co, b_BAR );
  input a, ci, b_BAR;
  output s, co;


  XNOR2X1 U1 ( .IN1(ci), .IN2(a), .Q(s) );
endmodule


module add_194 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_195 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_196 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_197 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_198 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_199 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_200 ( s, a, ci, co, b_BAR );
  input a, ci, b_BAR;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(b_BAR), .IN2(n1), .QN(co) );
  INVX0 U2 ( .INP(a), .ZN(n1) );
  MUX21X1 U3 ( .IN1(a), .IN2(n1), .S(b_BAR), .Q(s) );
endmodule


module adder8_13 ( out, a, b, cin );
  output [7:0] out;
  input [7:0] a;
  input [7:0] b;
  input cin;
  wire   n_1_net_, n_2_net_, n_3_net_, n_4_net_, n_5_net_, n_6_net_;
  wire   [6:0] c;

  add_200 add_01 ( .s(out[0]), .a(a[0]), .ci(1'b1), .co(c[0]), .b_BAR(b[0]) );
  add_199 add_02 ( .s(out[1]), .a(a[1]), .b(n_1_net_), .ci(c[0]), .co(c[1]) );
  add_198 add_03 ( .s(out[2]), .a(a[2]), .b(n_2_net_), .ci(c[1]), .co(c[2]) );
  add_197 add_04 ( .s(out[3]), .a(a[3]), .b(n_3_net_), .ci(c[2]), .co(c[3]) );
  add_196 add_05 ( .s(out[4]), .a(a[4]), .b(n_4_net_), .ci(c[3]), .co(c[4]) );
  add_195 add_06 ( .s(out[5]), .a(a[5]), .b(n_5_net_), .ci(c[4]), .co(c[5]) );
  add_194 add_07 ( .s(out[6]), .a(a[6]), .b(n_6_net_), .ci(c[5]), .co(c[6]) );
  add_193 add_08 ( .s(out[7]), .a(a[7]), .ci(c[6]), .b_BAR(1'b0) );
  INVX0 U1 ( .INP(b[1]), .ZN(n_1_net_) );
  INVX0 U2 ( .INP(b[2]), .ZN(n_2_net_) );
  INVX0 U3 ( .INP(b[3]), .ZN(n_3_net_) );
  INVX0 U4 ( .INP(b[4]), .ZN(n_4_net_) );
  INVX0 U5 ( .INP(b[5]), .ZN(n_5_net_) );
  INVX0 U6 ( .INP(b[6]), .ZN(n_6_net_) );
endmodule


module add_201 ( s, a, ci, co, b_BAR );
  input a, ci, b_BAR;
  output s, co;


  XNOR2X1 U1 ( .IN1(b_BAR), .IN2(ci), .Q(s) );
endmodule


module add_202 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_203 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_204 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_205 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_206 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_207 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_208 ( s, a, ci, co, b_BAR );
  input a, ci, b_BAR;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(b_BAR), .IN2(n1), .QN(co) );
  INVX0 U2 ( .INP(a), .ZN(n1) );
  MUX21X1 U3 ( .IN1(a), .IN2(n1), .S(b_BAR), .Q(s) );
endmodule


module adder8_14 ( out, a, b, cin );
  output [7:0] out;
  input [7:0] a;
  input [7:0] b;
  input cin;
  wire   n_1_net_, n_2_net_, n_3_net_, n_4_net_, n_5_net_, n_6_net_;
  wire   [6:0] c;

  add_208 add_01 ( .s(out[0]), .a(a[0]), .ci(1'b1), .co(c[0]), .b_BAR(b[0]) );
  add_207 add_02 ( .s(out[1]), .a(a[1]), .b(n_1_net_), .ci(c[0]), .co(c[1]) );
  add_206 add_03 ( .s(out[2]), .a(a[2]), .b(n_2_net_), .ci(c[1]), .co(c[2]) );
  add_205 add_04 ( .s(out[3]), .a(a[3]), .b(n_3_net_), .ci(c[2]), .co(c[3]) );
  add_204 add_05 ( .s(out[4]), .a(a[4]), .b(n_4_net_), .ci(c[3]), .co(c[4]) );
  add_203 add_06 ( .s(out[5]), .a(a[5]), .b(n_5_net_), .ci(c[4]), .co(c[5]) );
  add_202 add_07 ( .s(out[6]), .a(a[6]), .b(n_6_net_), .ci(c[5]), .co(c[6]) );
  add_201 add_08 ( .s(out[7]), .a(1'b0), .ci(c[6]), .b_BAR(b[7]) );
  INVX0 U1 ( .INP(b[1]), .ZN(n_1_net_) );
  INVX0 U2 ( .INP(b[2]), .ZN(n_2_net_) );
  INVX0 U3 ( .INP(b[3]), .ZN(n_3_net_) );
  INVX0 U4 ( .INP(b[4]), .ZN(n_4_net_) );
  INVX0 U5 ( .INP(b[5]), .ZN(n_5_net_) );
  INVX0 U6 ( .INP(b[6]), .ZN(n_6_net_) );
endmodule


module floating_point_adder_2 ( clk, rst_n, input_factor_01, input_factor_02, 
        output_adder );
  input [31:0] input_factor_01;
  input [31:0] input_factor_02;
  output [31:0] output_adder;
  input clk, rst_n;
  wire   N34, N35, N36, N37, N38, N39, N40, N41, N152, N153, N154, N155, N156,
         N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, N167,
         N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178,
         N179, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189,
         N190, N191, N192, N193, N194, N195, N196, N197, N198,
         add_sub_result_24_, N211, shift_temp_01_0_, N226, N227, N228, N229,
         N230, N231, N232, N233, N234, N235, N236, N237, N238, N239, N240,
         N241, N242, N243, N244, N245, N246, N247, N248, N256, N257, N258,
         N260, N261, N262, N263, N264, N265, N266, N267, N268, N269, N270,
         N271, N272, N273, N274, N275, N276, N277, N278, N279, N280, N281,
         N306, N307, N308, N346, N347, N348, N349, N350, N351, N352, N353,
         N354, N355, N380, N381, N382, N383, N384, N385, N386, N387, N388,
         N389, N390, N391, N392, N393, N394, N395, N396, N397, N398, N399,
         N400, N401, N402, N403, N404, N405, N406, N407, N408, N409, N410, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844;
  wire   [7:0] exp_diff_value;
  wire   [7:0] exponent_factor_21;
  wire   [7:0] exponent_factor_12;
  wire   [23:0] shift_smaller_factor;
  wire   [22:0] larger_factor;
  wire   [7:0] larger_exponent;
  wire   [24:0] add_result;
  wire   [24:0] sub_result;
  wire   [22:0] pre_sig_res_01;
  wire   [3:0] shift_temp_02;
  wire   [22:1] pre_sig_res_02;
  wire   [2:0] shift_temp_03;
  wire   [22:9] pre_sig_res_03;
  wire   [4:0] shift_temp_04;
  wire   [22:16] pre_sig_res_04;
  wire   [7:0] add_output_exponent_w1;
  wire   [7:0] add_output_exponent_w2;
  wire   [7:0] add_output_exponent_w3;
  wire   [7:0] add_output_exponent_w4;

  adder8_14 adder8_01 ( .out(exponent_factor_21), .a({1'b0, 
        input_factor_02[29:23]}), .b(input_factor_01[30:23]), .cin(1'b1) );
  adder8_13 adder8_02 ( .out(exponent_factor_12), .a(input_factor_01[30:23]), 
        .b({1'b0, input_factor_02[29:23]}), .cin(1'b1) );
  adder24_4 adder24_01 ( .clk(clk), .rst_n(rst_n), .a({shift_temp_04[4], 
        larger_factor}), .b(shift_smaller_factor), .cin(1'b1), .out(sub_result) );
  adder24_3 adder24_02 ( .clk(clk), .rst_n(rst_n), .a({shift_temp_04[4], 
        larger_factor}), .b(shift_smaller_factor), .cin(1'b0), .out(add_result) );
  adder8_12 adder8_03 ( .out(add_output_exponent_w1), .a(larger_exponent), .b(
        {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, shift_temp_01_0_}), .cin(
        1'b0) );
  adder8_11 adder8_04 ( .out(add_output_exponent_w2), .a(larger_exponent), .b(
        {1'b0, 1'b0, 1'b0, 1'b0, shift_temp_02}), .cin(1'b1) );
  adder8_10 adder8_05 ( .out(add_output_exponent_w3), .a(larger_exponent), .b(
        {1'b0, 1'b0, 1'b0, 1'b0, shift_temp_04[4], shift_temp_03}), .cin(1'b1)
         );
  adder8_9 adder8_06 ( .out(add_output_exponent_w4), .a(larger_exponent), .b({
        1'b0, 1'b0, 1'b0, shift_temp_04[4], 1'b0, shift_temp_04[2:0]}), .cin(
        1'b1) );
  DFFARX1 exp_diff_value_reg_7_ ( .D(N41), .CLK(clk), .RSTB(rst_n), .Q(
        exp_diff_value[7]) );
  DFFARX1 exp_diff_value_reg_6_ ( .D(N40), .CLK(clk), .RSTB(rst_n), .Q(
        exp_diff_value[6]) );
  DFFARX1 exp_diff_value_reg_5_ ( .D(N39), .CLK(clk), .RSTB(rst_n), .Q(
        exp_diff_value[5]) );
  DFFARX1 exp_diff_value_reg_4_ ( .D(N38), .CLK(clk), .RSTB(rst_n), .Q(
        exp_diff_value[4]) );
  DFFARX1 exp_diff_value_reg_3_ ( .D(N37), .CLK(clk), .RSTB(rst_n), .Q(
        exp_diff_value[3]), .QN(n4) );
  DFFARX1 exp_diff_value_reg_2_ ( .D(N36), .CLK(clk), .RSTB(rst_n), .Q(
        exp_diff_value[2]), .QN(n1) );
  DFFARX1 exp_diff_value_reg_1_ ( .D(N35), .CLK(clk), .RSTB(rst_n), .Q(
        exp_diff_value[1]), .QN(n2) );
  DFFARX1 exp_diff_value_reg_0_ ( .D(N34), .CLK(clk), .RSTB(rst_n), .Q(
        exp_diff_value[0]), .QN(n3) );
  DFFARX1 larger_factor_reg_22_ ( .D(N198), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[22]) );
  DFFARX1 larger_factor_reg_21_ ( .D(N197), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[21]) );
  DFFARX1 larger_factor_reg_20_ ( .D(N196), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[20]) );
  DFFARX1 larger_factor_reg_19_ ( .D(N195), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[19]) );
  DFFARX1 larger_factor_reg_18_ ( .D(N194), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[18]) );
  DFFARX1 larger_factor_reg_17_ ( .D(N193), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[17]) );
  DFFARX1 larger_factor_reg_16_ ( .D(N192), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[16]) );
  DFFARX1 larger_factor_reg_15_ ( .D(N191), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[15]) );
  DFFARX1 larger_factor_reg_14_ ( .D(N190), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[14]) );
  DFFARX1 larger_factor_reg_13_ ( .D(N189), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[13]) );
  DFFARX1 larger_factor_reg_12_ ( .D(N188), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[12]) );
  DFFARX1 larger_factor_reg_11_ ( .D(N187), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[11]) );
  DFFARX1 larger_factor_reg_10_ ( .D(N186), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[10]) );
  DFFARX1 larger_factor_reg_9_ ( .D(N185), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[9]) );
  DFFARX1 larger_factor_reg_8_ ( .D(N184), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[8]) );
  DFFARX1 larger_factor_reg_7_ ( .D(N183), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[7]) );
  DFFARX1 larger_factor_reg_6_ ( .D(N182), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[6]) );
  DFFARX1 larger_factor_reg_5_ ( .D(N181), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[5]) );
  DFFARX1 larger_factor_reg_4_ ( .D(N180), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[4]) );
  DFFARX1 larger_factor_reg_3_ ( .D(N179), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[3]) );
  DFFARX1 larger_factor_reg_2_ ( .D(N178), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[2]) );
  DFFARX1 larger_factor_reg_1_ ( .D(N177), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[1]) );
  DFFARX1 larger_factor_reg_0_ ( .D(N176), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[0]) );
  DFFARX1 shift_smaller_factor_reg_23_ ( .D(N175), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[23]) );
  DFFARX1 shift_smaller_factor_reg_22_ ( .D(N174), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[22]) );
  DFFARX1 shift_smaller_factor_reg_21_ ( .D(N173), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[21]) );
  DFFARX1 shift_smaller_factor_reg_20_ ( .D(N172), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[20]) );
  DFFARX1 shift_smaller_factor_reg_19_ ( .D(N171), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[19]) );
  DFFARX1 shift_smaller_factor_reg_18_ ( .D(N170), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[18]) );
  DFFARX1 shift_smaller_factor_reg_17_ ( .D(N169), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[17]) );
  DFFARX1 shift_smaller_factor_reg_16_ ( .D(N168), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[16]) );
  DFFARX1 shift_smaller_factor_reg_15_ ( .D(N167), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[15]) );
  DFFARX1 shift_smaller_factor_reg_14_ ( .D(N166), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[14]) );
  DFFARX1 shift_smaller_factor_reg_13_ ( .D(N165), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[13]) );
  DFFARX1 shift_smaller_factor_reg_12_ ( .D(N164), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[12]) );
  DFFARX1 shift_smaller_factor_reg_11_ ( .D(N163), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[11]) );
  DFFARX1 shift_smaller_factor_reg_10_ ( .D(N162), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[10]) );
  DFFARX1 shift_smaller_factor_reg_9_ ( .D(N161), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[9]) );
  DFFARX1 shift_smaller_factor_reg_8_ ( .D(N160), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[8]) );
  DFFARX1 shift_smaller_factor_reg_7_ ( .D(N159), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[7]) );
  DFFARX1 shift_smaller_factor_reg_6_ ( .D(N158), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[6]) );
  DFFARX1 shift_smaller_factor_reg_5_ ( .D(N157), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[5]) );
  DFFARX1 shift_smaller_factor_reg_4_ ( .D(N156), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[4]) );
  DFFARX1 shift_smaller_factor_reg_3_ ( .D(N155), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[3]) );
  DFFARX1 shift_smaller_factor_reg_2_ ( .D(N154), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[2]) );
  DFFARX1 shift_smaller_factor_reg_1_ ( .D(N153), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[1]) );
  DFFARX1 shift_smaller_factor_reg_0_ ( .D(N152), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[0]) );
  DFFX1 larger_exponent_reg_7_ ( .D(n822), .CLK(clk), .Q(larger_exponent[7])
         );
  DFFX1 larger_exponent_reg_6_ ( .D(n823), .CLK(clk), .Q(larger_exponent[6])
         );
  DFFX1 larger_exponent_reg_5_ ( .D(n824), .CLK(clk), .Q(larger_exponent[5])
         );
  DFFX1 larger_exponent_reg_4_ ( .D(n825), .CLK(clk), .Q(larger_exponent[4])
         );
  DFFX1 larger_exponent_reg_3_ ( .D(n826), .CLK(clk), .Q(larger_exponent[3])
         );
  DFFX1 larger_exponent_reg_2_ ( .D(n827), .CLK(clk), .Q(larger_exponent[2])
         );
  DFFX1 larger_exponent_reg_1_ ( .D(n828), .CLK(clk), .Q(larger_exponent[1])
         );
  DFFX1 larger_exponent_reg_0_ ( .D(n829), .CLK(clk), .Q(larger_exponent[0])
         );
  DFFARX1 shift_temp_04_reg_4_ ( .D(1'b1), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_04[4]) );
  DFFARX1 shift_temp_01_reg_0_ ( .D(add_sub_result_24_), .CLK(clk), .RSTB(
        rst_n), .Q(shift_temp_01_0_) );
  DFFARX1 pre_sig_res_02_reg_1_ ( .D(N260), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[1]) );
  DFFARX1 pre_sig_res_02_reg_2_ ( .D(N261), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[2]) );
  DFFARX1 pre_sig_res_02_reg_3_ ( .D(N262), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[3]) );
  DFFARX1 pre_sig_res_02_reg_4_ ( .D(N263), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[4]) );
  DFFARX1 pre_sig_res_02_reg_5_ ( .D(N264), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[5]) );
  DFFARX1 pre_sig_res_02_reg_6_ ( .D(N265), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[6]) );
  DFFARX1 pre_sig_res_02_reg_7_ ( .D(N266), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[7]) );
  DFFARX1 shift_temp_02_reg_2_ ( .D(N258), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_02[2]) );
  DFFASX1 shift_temp_02_reg_3_ ( .D(n821), .CLK(clk), .SETB(rst_n), .QN(
        shift_temp_02[3]) );
  DFFARX1 pre_sig_res_02_reg_8_ ( .D(N267), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[8]) );
  DFFARX1 pre_sig_res_02_reg_9_ ( .D(N268), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[9]) );
  DFFARX1 pre_sig_res_02_reg_10_ ( .D(N269), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[10]) );
  DFFARX1 pre_sig_res_02_reg_11_ ( .D(N270), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[11]) );
  DFFARX1 pre_sig_res_02_reg_12_ ( .D(N271), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[12]) );
  DFFARX1 pre_sig_res_02_reg_13_ ( .D(N272), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[13]) );
  DFFARX1 pre_sig_res_02_reg_14_ ( .D(N273), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[14]) );
  DFFARX1 pre_sig_res_02_reg_15_ ( .D(N274), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[15]) );
  DFFARX1 pre_sig_res_02_reg_16_ ( .D(N275), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[16]) );
  DFFARX1 pre_sig_res_02_reg_17_ ( .D(N276), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[17]) );
  DFFARX1 pre_sig_res_02_reg_18_ ( .D(N277), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[18]) );
  DFFARX1 pre_sig_res_02_reg_19_ ( .D(N278), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[19]) );
  DFFARX1 pre_sig_res_02_reg_20_ ( .D(N279), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[20]) );
  DFFARX1 pre_sig_res_02_reg_21_ ( .D(N280), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[21]) );
  DFFARX1 pre_sig_res_02_reg_22_ ( .D(N281), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[22]) );
  DFFARX1 shift_temp_02_reg_1_ ( .D(N257), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_02[1]) );
  DFFARX1 shift_temp_02_reg_0_ ( .D(N256), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_02[0]) );
  DFFX1 pre_sig_res_03_reg_9_ ( .D(n830), .CLK(clk), .Q(pre_sig_res_03[9]) );
  DFFX1 pre_sig_res_03_reg_10_ ( .D(n831), .CLK(clk), .Q(pre_sig_res_03[10])
         );
  DFFX1 pre_sig_res_03_reg_12_ ( .D(n832), .CLK(clk), .Q(pre_sig_res_03[12])
         );
  DFFX1 pre_sig_res_03_reg_11_ ( .D(n833), .CLK(clk), .Q(pre_sig_res_03[11])
         );
  DFFX1 pre_sig_res_03_reg_13_ ( .D(n834), .CLK(clk), .Q(pre_sig_res_03[13])
         );
  DFFX1 pre_sig_res_03_reg_14_ ( .D(n835), .CLK(clk), .Q(pre_sig_res_03[14])
         );
  DFFARX1 shift_temp_03_reg_2_ ( .D(N308), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_03[2]) );
  DFFARX1 shift_temp_03_reg_0_ ( .D(N306), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_03[0]) );
  DFFARX1 shift_temp_03_reg_1_ ( .D(N307), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_03[1]) );
  DFFX1 pre_sig_res_03_reg_15_ ( .D(n836), .CLK(clk), .Q(pre_sig_res_03[15])
         );
  DFFX1 pre_sig_res_03_reg_16_ ( .D(n837), .CLK(clk), .Q(pre_sig_res_03[16])
         );
  DFFX1 pre_sig_res_03_reg_17_ ( .D(n838), .CLK(clk), .Q(pre_sig_res_03[17])
         );
  DFFX1 pre_sig_res_03_reg_18_ ( .D(n839), .CLK(clk), .Q(pre_sig_res_03[18])
         );
  DFFX1 pre_sig_res_03_reg_19_ ( .D(n840), .CLK(clk), .Q(pre_sig_res_03[19])
         );
  DFFX1 pre_sig_res_03_reg_20_ ( .D(n841), .CLK(clk), .Q(pre_sig_res_03[20])
         );
  DFFX1 pre_sig_res_03_reg_21_ ( .D(n842), .CLK(clk), .Q(pre_sig_res_03[21])
         );
  DFFX1 pre_sig_res_03_reg_22_ ( .D(n843), .CLK(clk), .Q(pre_sig_res_03[22])
         );
  DFFARX1 pre_sig_res_04_reg_16_ ( .D(N349), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_04[16]) );
  DFFARX1 pre_sig_res_04_reg_17_ ( .D(N350), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_04[17]) );
  DFFARX1 pre_sig_res_04_reg_18_ ( .D(N351), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_04[18]) );
  DFFARX1 pre_sig_res_04_reg_19_ ( .D(N352), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_04[19]) );
  DFFARX1 pre_sig_res_04_reg_20_ ( .D(N353), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_04[20]) );
  DFFARX1 pre_sig_res_04_reg_21_ ( .D(N354), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_04[21]) );
  DFFARX1 pre_sig_res_04_reg_22_ ( .D(N355), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_04[22]) );
  DFFARX1 add_output_sign_reg ( .D(N211), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[31]) );
  DFFARX1 pre_sig_res_01_reg_0_ ( .D(N226), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[0]) );
  DFFARX1 pre_sig_res_01_reg_1_ ( .D(N227), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[1]) );
  DFFARX1 pre_sig_res_01_reg_2_ ( .D(N228), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[2]) );
  DFFARX1 pre_sig_res_01_reg_3_ ( .D(N229), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[3]) );
  DFFARX1 pre_sig_res_01_reg_4_ ( .D(N230), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[4]) );
  DFFARX1 pre_sig_res_01_reg_5_ ( .D(N231), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[5]) );
  DFFARX1 pre_sig_res_01_reg_6_ ( .D(N232), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[6]) );
  DFFARX1 pre_sig_res_01_reg_7_ ( .D(N233), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[7]) );
  DFFARX1 pre_sig_res_01_reg_8_ ( .D(N234), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[8]) );
  DFFARX1 pre_sig_res_01_reg_9_ ( .D(N235), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[9]) );
  DFFARX1 pre_sig_res_01_reg_10_ ( .D(N236), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[10]) );
  DFFARX1 pre_sig_res_01_reg_11_ ( .D(N237), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[11]) );
  DFFARX1 pre_sig_res_01_reg_12_ ( .D(N238), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[12]) );
  DFFARX1 pre_sig_res_01_reg_13_ ( .D(N239), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[13]) );
  DFFARX1 pre_sig_res_01_reg_14_ ( .D(N240), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[14]) );
  DFFARX1 pre_sig_res_01_reg_15_ ( .D(N241), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[15]) );
  DFFARX1 pre_sig_res_01_reg_16_ ( .D(N242), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[16]) );
  DFFARX1 pre_sig_res_01_reg_17_ ( .D(N243), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[17]) );
  DFFARX1 pre_sig_res_01_reg_18_ ( .D(N244), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[18]) );
  DFFARX1 pre_sig_res_01_reg_19_ ( .D(N245), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[19]) );
  DFFARX1 pre_sig_res_01_reg_20_ ( .D(N246), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[20]) );
  DFFARX1 pre_sig_res_01_reg_21_ ( .D(N247), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[21]) );
  DFFARX1 pre_sig_res_01_reg_22_ ( .D(N248), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[22]) );
  DFFARX1 shift_temp_04_reg_2_ ( .D(N348), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_04[2]) );
  DFFARX1 shift_temp_04_reg_1_ ( .D(N347), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_04[1]) );
  DFFARX1 shift_temp_04_reg_0_ ( .D(N346), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_04[0]) );
  DFFARX1 add_output_exponent_reg_7_ ( .D(N387), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[30]) );
  DFFARX1 add_output_exponent_reg_6_ ( .D(N386), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[29]) );
  DFFARX1 add_output_exponent_reg_5_ ( .D(N385), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[28]) );
  DFFARX1 add_output_exponent_reg_4_ ( .D(N384), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[27]) );
  DFFARX1 add_output_exponent_reg_3_ ( .D(N383), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[26]) );
  DFFARX1 add_output_exponent_reg_2_ ( .D(N382), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[25]) );
  DFFARX1 add_output_exponent_reg_1_ ( .D(N381), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[24]) );
  DFFARX1 add_output_exponent_reg_0_ ( .D(N380), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[23]) );
  DFFARX1 add_output_significands_reg_22_ ( .D(N410), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[22]) );
  DFFARX1 add_output_significands_reg_21_ ( .D(N409), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[21]) );
  DFFARX1 add_output_significands_reg_20_ ( .D(N408), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[20]) );
  DFFARX1 add_output_significands_reg_19_ ( .D(N407), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[19]) );
  DFFARX1 add_output_significands_reg_18_ ( .D(N406), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[18]) );
  DFFARX1 add_output_significands_reg_17_ ( .D(N405), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[17]) );
  DFFARX1 add_output_significands_reg_16_ ( .D(N404), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[16]) );
  DFFARX1 add_output_significands_reg_15_ ( .D(N403), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[15]) );
  DFFARX1 add_output_significands_reg_14_ ( .D(N402), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[14]) );
  DFFARX1 add_output_significands_reg_13_ ( .D(N401), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[13]) );
  DFFARX1 add_output_significands_reg_12_ ( .D(N400), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[12]) );
  DFFARX1 add_output_significands_reg_11_ ( .D(N399), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[11]) );
  DFFARX1 add_output_significands_reg_10_ ( .D(N398), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[10]) );
  DFFARX1 add_output_significands_reg_9_ ( .D(N397), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[9]) );
  DFFARX1 add_output_significands_reg_8_ ( .D(N396), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[8]) );
  DFFARX1 add_output_significands_reg_7_ ( .D(N395), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[7]) );
  DFFARX1 add_output_significands_reg_6_ ( .D(N394), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[6]) );
  DFFARX1 add_output_significands_reg_5_ ( .D(N393), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[5]) );
  DFFARX1 add_output_significands_reg_4_ ( .D(N392), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[4]) );
  DFFARX1 add_output_significands_reg_3_ ( .D(N391), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[3]) );
  DFFARX1 add_output_significands_reg_2_ ( .D(N390), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[2]) );
  DFFARX1 add_output_significands_reg_1_ ( .D(N389), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[1]) );
  DFFARX1 add_output_significands_reg_0_ ( .D(N388), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[0]) );
  INVX1 U5 ( .INP(rst_n), .ZN(n844) );
  NAND2X0 U3 ( .IN1(input_factor_02[11]), .IN2(n638), .QN(n57) );
  NAND2X0 U4 ( .IN1(n482), .IN2(n395), .QN(n562) );
  NAND2X0 U6 ( .IN1(input_factor_02[16]), .IN2(n370), .QN(n70) );
  NAND2X0 U7 ( .IN1(input_factor_02[24]), .IN2(n541), .QN(n34) );
  NAND2X0 U8 ( .IN1(input_factor_01[27]), .IN2(n588), .QN(n30) );
  NAND2X0 U9 ( .IN1(input_factor_01[26]), .IN2(n582), .QN(n31) );
  NAND2X0 U10 ( .IN1(input_factor_01[28]), .IN2(n594), .QN(n41) );
  NAND2X0 U11 ( .IN1(input_factor_02[28]), .IN2(n593), .QN(n45) );
  NAND2X0 U12 ( .IN1(n801), .IN2(n522), .QN(n381) );
  NAND2X0 U13 ( .IN1(n771), .IN2(n514), .QN(n380) );
  NAND2X0 U14 ( .IN1(n764), .IN2(n515), .QN(n379) );
  NAND2X0 U15 ( .IN1(n740), .IN2(n714), .QN(n559) );
  NAND2X0 U16 ( .IN1(n399), .IN2(n492), .QN(n377) );
  NAND2X0 U17 ( .IN1(n490), .IN2(n402), .QN(n376) );
  NAND2X0 U18 ( .IN1(n375), .IN2(n568), .QN(n401) );
  NAND2X0 U19 ( .IN1(n91), .IN2(n90), .QN(n217) );
  NAND2X0 U20 ( .IN1(n166), .IN2(n165), .QN(n250) );
  NAND2X0 U21 ( .IN1(n200), .IN2(n199), .QN(n269) );
  NAND2X0 U22 ( .IN1(exp_diff_value[1]), .IN2(exp_diff_value[0]), .QN(n198) );
  NAND2X0 U23 ( .IN1(exp_diff_value[1]), .IN2(n3), .QN(n196) );
  NAND2X0 U24 ( .IN1(exp_diff_value[0]), .IN2(n2), .QN(n197) );
  NAND2X0 U25 ( .IN1(n353), .IN2(n217), .QN(n218) );
  NAND2X0 U26 ( .IN1(n698), .IN2(n268), .QN(n248) );
  NAND2X0 U27 ( .IN1(n164), .IN2(n163), .QN(n246) );
  NAND2X0 U28 ( .IN1(n353), .IN2(n250), .QN(n251) );
  NAND2X0 U29 ( .IN1(n268), .IN2(n817), .QN(n252) );
  NAND2X0 U30 ( .IN1(n195), .IN2(n194), .QN(n265) );
  NAND2X0 U31 ( .IN1(n353), .IN2(n269), .QN(n270) );
  NAND2X0 U32 ( .IN1(n126), .IN2(n125), .QN(n230) );
  NAND2X0 U33 ( .IN1(n70), .IN2(n71), .QN(n18) );
  NAND2X0 U34 ( .IN1(n693), .IN2(n2), .QN(n120) );
  NAND2X0 U35 ( .IN1(input_factor_02[19]), .IN2(n683), .QN(n65) );
  NAND2X0 U36 ( .IN1(n702), .IN2(n3), .QN(n147) );
  NAND2X0 U37 ( .IN1(input_factor_01[23]), .IN2(n557), .QN(n32) );
  NAND2X0 U38 ( .IN1(n542), .IN2(input_factor_02[25]), .QN(n33) );
  NAND2X0 U39 ( .IN1(input_factor_02[27]), .IN2(n587), .QN(n24) );
  NAND2X0 U40 ( .IN1(input_factor_02[26]), .IN2(n581), .QN(n22) );
  NAND2X0 U41 ( .IN1(n373), .IN2(n74), .QN(n176) );
  NAND2X0 U42 ( .IN1(n706), .IN2(pre_sig_res_01[9]), .QN(n630) );
  NAND2X0 U43 ( .IN1(n706), .IN2(pre_sig_res_01[10]), .QN(n636) );
  NAND2X0 U44 ( .IN1(n706), .IN2(pre_sig_res_01[11]), .QN(n642) );
  NAND2X0 U45 ( .IN1(n706), .IN2(pre_sig_res_01[13]), .QN(n651) );
  NAND2X0 U46 ( .IN1(n706), .IN2(pre_sig_res_01[14]), .QN(n657) );
  NAND2X0 U47 ( .IN1(n706), .IN2(pre_sig_res_01[15]), .QN(n663) );
  NAND2X0 U48 ( .IN1(n706), .IN2(pre_sig_res_01[16]), .QN(n667) );
  NAND2X0 U49 ( .IN1(n706), .IN2(pre_sig_res_01[17]), .QN(n673) );
  NAND2X0 U50 ( .IN1(n706), .IN2(pre_sig_res_01[18]), .QN(n679) );
  NAND2X0 U51 ( .IN1(n706), .IN2(pre_sig_res_01[19]), .QN(n685) );
  NAND2X0 U52 ( .IN1(n706), .IN2(pre_sig_res_01[21]), .QN(n694) );
  NAND2X0 U53 ( .IN1(n706), .IN2(pre_sig_res_01[22]), .QN(n707) );
  NAND2X0 U54 ( .IN1(n706), .IN2(add_output_exponent_w1[0]), .QN(n569) );
  NAND2X0 U55 ( .IN1(n706), .IN2(add_output_exponent_w1[1]), .QN(n573) );
  NAND2X0 U56 ( .IN1(n706), .IN2(add_output_exponent_w1[2]), .QN(n577) );
  NAND2X0 U57 ( .IN1(n706), .IN2(add_output_exponent_w1[3]), .QN(n583) );
  NAND2X0 U58 ( .IN1(n706), .IN2(add_output_exponent_w1[4]), .QN(n589) );
  NAND2X0 U59 ( .IN1(n706), .IN2(add_output_exponent_w1[5]), .QN(n595) );
  NAND2X0 U60 ( .IN1(n706), .IN2(add_output_exponent_w1[6]), .QN(n601) );
  NAND2X0 U61 ( .IN1(n516), .IN2(n811), .QN(n534) );
  NAND2X0 U62 ( .IN1(n513), .IN2(n522), .QN(n519) );
  NAND2X0 U63 ( .IN1(n176), .IN2(n360), .QN(n391) );
  NAND2X0 U64 ( .IN1(n514), .IN2(n784), .QN(n532) );
  NAND2X0 U65 ( .IN1(n515), .IN2(n751), .QN(n533) );
  NAND2X0 U66 ( .IN1(n756), .IN2(n740), .QN(n715) );
  NAND2X0 U67 ( .IN1(n714), .IN2(n727), .QN(n789) );
  NAND2X0 U68 ( .IN1(n512), .IN2(n500), .QN(n718) );
  NAND2X0 U69 ( .IN1(n512), .IN2(n504), .QN(n711) );
  NAND2X0 U70 ( .IN1(n395), .IN2(n394), .QN(n494) );
  NAND2X0 U71 ( .IN1(n412), .IN2(n813), .QN(n409) );
  NAND2X0 U72 ( .IN1(n399), .IN2(n396), .QN(n483) );
  NAND2X0 U73 ( .IN1(n402), .IN2(n397), .QN(n487) );
  NAND2X0 U74 ( .IN1(n398), .IN2(n568), .QN(n485) );
  NAND2X0 U75 ( .IN1(n162), .IN2(n161), .QN(n167) );
  NAND2X0 U76 ( .IN1(n268), .IN2(n4), .QN(n177) );
  NAND2X0 U77 ( .IN1(n817), .IN2(n372), .QN(n271) );
  NAND2X0 U78 ( .IN1(n698), .IN2(n372), .QN(n232) );
  NAND2X0 U79 ( .IN1(n191), .IN2(n190), .QN(n201) );
  NAND2X0 U80 ( .IN1(n89), .IN2(n88), .QN(n215) );
  NAND2X0 U81 ( .IN1(n218), .IN2(n219), .QN(n16) );
  NAND2X0 U82 ( .IN1(n4), .IN2(n1), .QN(n275) );
  NAND2X0 U83 ( .IN1(n251), .IN2(n253), .QN(n14) );
  NAND2X0 U84 ( .IN1(n354), .IN2(n207), .QN(n262) );
  NAND2X0 U85 ( .IN1(n270), .IN2(n273), .QN(n12) );
  NAND2X0 U86 ( .IN1(exp_diff_value[3]), .IN2(n354), .QN(n330) );
  NAND2X0 U87 ( .IN1(n307), .IN2(n1), .QN(n322) );
  NAND2X0 U88 ( .IN1(n330), .IN2(n329), .QN(n331) );
  NAND2X0 U89 ( .IN1(n353), .IN2(n4), .QN(n347) );
  NAND2X0 U90 ( .IN1(n354), .IN2(n4), .QN(n349) );
  NAND2X0 U91 ( .IN1(n363), .IN2(n69), .QN(n360) );
  NAND2X0 U92 ( .IN1(n2), .IN2(n147), .QN(n367) );
  NAND2X0 U93 ( .IN1(n371), .IN2(n353), .QN(n366) );
  NAND2X0 U94 ( .IN1(n354), .IN2(n371), .QN(n364) );
  NAND2X0 U95 ( .IN1(n608), .IN2(n607), .QN(N390) );
  NAND2X0 U96 ( .IN1(n610), .IN2(n609), .QN(N391) );
  NAND2X0 U97 ( .IN1(n612), .IN2(n611), .QN(N392) );
  NAND2X0 U98 ( .IN1(n616), .IN2(n615), .QN(N393) );
  NAND2X0 U99 ( .IN1(n618), .IN2(n617), .QN(N394) );
  NAND2X0 U100 ( .IN1(n621), .IN2(n620), .QN(N395) );
  NAND2X0 U101 ( .IN1(n625), .IN2(n624), .QN(N396) );
  NAND2X0 U102 ( .IN1(n704), .IN2(pre_sig_res_03[9]), .QN(n628) );
  NAND2X0 U103 ( .IN1(n703), .IN2(pre_sig_res_02[9]), .QN(n629) );
  NAND2X0 U104 ( .IN1(n704), .IN2(pre_sig_res_03[10]), .QN(n634) );
  NAND2X0 U105 ( .IN1(n703), .IN2(pre_sig_res_02[10]), .QN(n635) );
  NAND2X0 U106 ( .IN1(n704), .IN2(pre_sig_res_03[11]), .QN(n640) );
  NAND2X0 U107 ( .IN1(n703), .IN2(pre_sig_res_02[11]), .QN(n641) );
  NAND2X0 U108 ( .IN1(n7), .IN2(n8), .QN(N400) );
  NAND2X0 U109 ( .IN1(pre_sig_res_01[12]), .IN2(n706), .QN(n8) );
  NAND2X0 U110 ( .IN1(n704), .IN2(pre_sig_res_03[13]), .QN(n649) );
  NAND2X0 U111 ( .IN1(n703), .IN2(pre_sig_res_02[13]), .QN(n650) );
  NAND2X0 U112 ( .IN1(n704), .IN2(pre_sig_res_03[14]), .QN(n655) );
  NAND2X0 U113 ( .IN1(n703), .IN2(pre_sig_res_02[14]), .QN(n656) );
  NAND2X0 U114 ( .IN1(n704), .IN2(pre_sig_res_03[15]), .QN(n661) );
  NAND2X0 U115 ( .IN1(n703), .IN2(pre_sig_res_02[15]), .QN(n662) );
  NAND2X0 U116 ( .IN1(n705), .IN2(pre_sig_res_04[16]), .QN(n668) );
  NAND2X0 U117 ( .IN1(n705), .IN2(pre_sig_res_04[17]), .QN(n674) );
  NAND2X0 U118 ( .IN1(n705), .IN2(pre_sig_res_04[18]), .QN(n680) );
  NAND2X0 U119 ( .IN1(n705), .IN2(pre_sig_res_04[19]), .QN(n686) );
  NAND2X0 U120 ( .IN1(n5), .IN2(n6), .QN(N408) );
  NAND2X0 U121 ( .IN1(n705), .IN2(pre_sig_res_04[20]), .QN(n6) );
  NAND2X0 U122 ( .IN1(n705), .IN2(pre_sig_res_04[21]), .QN(n695) );
  NAND2X0 U123 ( .IN1(n705), .IN2(pre_sig_res_04[22]), .QN(n708) );
  NAND2X0 U124 ( .IN1(n705), .IN2(add_output_exponent_w4[0]), .QN(n570) );
  NAND2X0 U125 ( .IN1(n705), .IN2(add_output_exponent_w4[1]), .QN(n574) );
  NAND2X0 U126 ( .IN1(n705), .IN2(add_output_exponent_w4[2]), .QN(n578) );
  NAND2X0 U127 ( .IN1(n705), .IN2(add_output_exponent_w4[3]), .QN(n584) );
  NAND2X0 U128 ( .IN1(n705), .IN2(add_output_exponent_w4[4]), .QN(n590) );
  NAND2X0 U129 ( .IN1(n705), .IN2(add_output_exponent_w4[5]), .QN(n596) );
  NAND2X0 U130 ( .IN1(n705), .IN2(add_output_exponent_w4[6]), .QN(n602) );
  NAND2X0 U131 ( .IN1(n9), .IN2(n10), .QN(N387) );
  NAND2X0 U132 ( .IN1(n705), .IN2(add_output_exponent_w4[7]), .QN(n10) );
  NAND2X0 U133 ( .IN1(n519), .IN2(n518), .QN(N348) );
  NAND2X0 U134 ( .IN1(n536), .IN2(n791), .QN(n537) );
  NAND2X0 U135 ( .IN1(n536), .IN2(n811), .QN(n527) );
  NAND2X0 U136 ( .IN1(n536), .IN2(n813), .QN(n523) );
  NAND2X0 U137 ( .IN1(n521), .IN2(n520), .QN(N352) );
  NAND2X0 U138 ( .IN1(pre_sig_res_03[22]), .IN2(n815), .QN(n720) );
  NAND2X0 U139 ( .IN1(n804), .IN2(n719), .QN(n721) );
  NAND2X0 U140 ( .IN1(pre_sig_res_03[21]), .IN2(n815), .QN(n728) );
  NAND2X0 U141 ( .IN1(n804), .IN2(n727), .QN(n729) );
  NAND2X0 U142 ( .IN1(pre_sig_res_03[20]), .IN2(n815), .QN(n736) );
  NAND2X0 U143 ( .IN1(n804), .IN2(n735), .QN(n737) );
  NAND2X0 U144 ( .IN1(pre_sig_res_03[19]), .IN2(n815), .QN(n744) );
  NAND2X0 U145 ( .IN1(n804), .IN2(n743), .QN(n745) );
  NAND2X0 U146 ( .IN1(pre_sig_res_03[18]), .IN2(n815), .QN(n752) );
  NAND2X0 U147 ( .IN1(n804), .IN2(n751), .QN(n753) );
  NAND2X0 U148 ( .IN1(pre_sig_res_03[17]), .IN2(n815), .QN(n760) );
  NAND2X0 U149 ( .IN1(n804), .IN2(n759), .QN(n761) );
  NAND2X0 U150 ( .IN1(pre_sig_res_03[16]), .IN2(n815), .QN(n767) );
  NAND2X0 U151 ( .IN1(n804), .IN2(n784), .QN(n768) );
  NAND2X0 U152 ( .IN1(pre_sig_res_03[15]), .IN2(n815), .QN(n776) );
  NAND2X0 U153 ( .IN1(n804), .IN2(n792), .QN(n777) );
  NAND2X0 U154 ( .IN1(n711), .IN2(n718), .QN(n505) );
  NAND2X0 U155 ( .IN1(pre_sig_res_03[14]), .IN2(n844), .QN(n786) );
  NAND2X0 U156 ( .IN1(n814), .IN2(n784), .QN(n785) );
  NAND2X0 U157 ( .IN1(n804), .IN2(n783), .QN(n787) );
  NAND2X0 U158 ( .IN1(pre_sig_res_03[13]), .IN2(n815), .QN(n794) );
  NAND2X0 U159 ( .IN1(n814), .IN2(n792), .QN(n793) );
  NAND2X0 U160 ( .IN1(n804), .IN2(n791), .QN(n795) );
  NAND2X0 U161 ( .IN1(n799), .IN2(n798), .QN(n833) );
  NAND2X0 U162 ( .IN1(pre_sig_res_03[12]), .IN2(n815), .QN(n807) );
  NAND2X0 U163 ( .IN1(n804), .IN2(n811), .QN(n809) );
  NAND2X0 U164 ( .IN1(n412), .IN2(n811), .QN(n413) );
  NAND2X0 U165 ( .IN1(n417), .IN2(n792), .QN(n408) );
  NAND2X0 U166 ( .IN1(n418), .IN2(n791), .QN(n405) );
  NAND2X0 U167 ( .IN1(n404), .IN2(n403), .QN(N263) );
  NAND2X0 U168 ( .IN1(n308), .IN2(input_factor_01[0]), .QN(n119) );
  NAND2X0 U169 ( .IN1(n146), .IN2(n145), .QN(N153) );
  NAND2X0 U170 ( .IN1(n308), .IN2(input_factor_01[2]), .QN(n172) );
  NAND2X0 U171 ( .IN1(n308), .IN2(input_factor_01[3]), .QN(n206) );
  NAND2X0 U172 ( .IN1(input_factor_01[4]), .IN2(n308), .QN(n222) );
  NAND2X0 U173 ( .IN1(input_factor_01[6]), .IN2(n308), .QN(n256) );
  NAND2X0 U174 ( .IN1(input_factor_01[7]), .IN2(n308), .QN(n277) );
  NAND2X0 U175 ( .IN1(input_factor_01[12]), .IN2(n308), .QN(n309) );
  NAND2X0 U176 ( .IN1(n338), .IN2(n337), .QN(N168) );
  NAND2X0 U177 ( .IN1(n342), .IN2(n341), .QN(N169) );
  NAND2X0 U178 ( .IN1(n346), .IN2(n345), .QN(N170) );
  NAND2X0 U179 ( .IN1(n352), .IN2(n351), .QN(N171) );
  NAND2X0 U180 ( .IN1(n362), .IN2(n361), .QN(N173) );
  NAND2X0 U181 ( .IN1(n369), .IN2(n368), .QN(N174) );
  NAND2X0 U182 ( .IN1(n374), .IN2(n373), .QN(N175) );
  INVX0 U183 ( .INP(n391), .ZN(n390) );
  NOR2X0 U184 ( .IN1(n817), .IN2(n844), .QN(n818) );
  NOR2X0 U185 ( .IN1(n816), .IN2(n815), .QN(n819) );
  INVX0 U186 ( .INP(n561), .ZN(n821) );
  INVX0 U187 ( .INP(n417), .ZN(n489) );
  NOR2X0 U188 ( .IN1(n718), .IN2(n815), .QN(n804) );
  INVX0 U189 ( .INP(n812), .ZN(n802) );
  INVX0 U190 ( .INP(n791), .ZN(n803) );
  INVX0 U191 ( .INP(n792), .ZN(n781) );
  INVX0 U192 ( .INP(n759), .ZN(n772) );
  NOR2X0 U193 ( .IN1(n564), .IN2(n567), .QN(n703) );
  NOR2X0 U194 ( .IN1(n565), .IN2(n567), .QN(n704) );
  INVX0 U195 ( .INP(n735), .ZN(n748) );
  INVX0 U196 ( .INP(n454), .ZN(n563) );
  INVX0 U197 ( .INP(n562), .ZN(n512) );
  INVX0 U198 ( .INP(n743), .ZN(n756) );
  NOR2X0 U199 ( .IN1(n568), .IN2(n567), .QN(n706) );
  INVX0 U200 ( .INP(n689), .ZN(n700) );
  NAND2X0 U201 ( .IN1(exp_diff_value[2]), .IN2(n4), .QN(n214) );
  INVX0 U202 ( .INP(n197), .ZN(n185) );
  INVX0 U203 ( .INP(n196), .ZN(n193) );
  NOR2X0 U204 ( .IN1(n363), .IN2(n74), .QN(n817) );
  INVX0 U205 ( .INP(n308), .ZN(n359) );
  NOR2X0 U206 ( .IN1(exp_diff_value[1]), .IN2(exp_diff_value[0]), .QN(n370) );
  INVX0 U207 ( .INP(n176), .ZN(n698) );
  INVX0 U208 ( .INP(n396), .ZN(n492) );
  NOR2X0 U209 ( .IN1(add_sub_result_24_), .IN2(n393), .QN(n568) );
  MUX21X1 U210 ( .IN1(add_result[24]), .IN2(sub_result[24]), .S(n20), .Q(
        add_sub_result_24_) );
  INVX0 U211 ( .INP(n394), .ZN(n482) );
  INVX0 U212 ( .INP(n21), .ZN(n20) );
  INVX0 U213 ( .INP(n501), .ZN(n21) );
  INVX0 U214 ( .INP(n727), .ZN(n740) );
  INVX0 U215 ( .INP(n751), .ZN(n764) );
  INVX0 U216 ( .INP(n784), .ZN(n771) );
  INVX0 U217 ( .INP(n783), .ZN(n801) );
  INVX0 U218 ( .INP(n811), .ZN(n797) );
  INVX0 U219 ( .INP(n813), .ZN(n805) );
  MUX21X1 U220 ( .IN1(input_factor_01[31]), .IN2(n547), .S(input_factor_02[31]), .Q(n501) );
  INVX0 U221 ( .INP(input_factor_01[31]), .ZN(n547) );
  INVX0 U222 ( .INP(n373), .ZN(n363) );
  NAND2X0 U223 ( .IN1(input_factor_02[29]), .IN2(n599), .QN(n46) );
  INVX0 U224 ( .INP(input_factor_02[23]), .ZN(n557) );
  INVX0 U225 ( .INP(input_factor_02[29]), .ZN(n600) );
  NAND4X0 U226 ( .IN1(n29), .IN2(n28), .IN3(n543), .IN4(n32), .QN(n373) );
  INVX0 U227 ( .INP(n445), .ZN(n713) );
  INVX0 U228 ( .INP(n719), .ZN(n732) );
  INVX0 U229 ( .INP(n814), .ZN(n800) );
  INVX0 U230 ( .INP(n440), .ZN(n724) );
  NOR2X0 U231 ( .IN1(n15), .IN2(n16), .QN(n221) );
  NOR2X0 U232 ( .IN1(n355), .IN2(n252), .QN(n15) );
  NOR2X0 U233 ( .IN1(n646), .IN2(n645), .QN(n7) );
  NOR2X0 U234 ( .IN1(n13), .IN2(n14), .QN(n255) );
  NOR2X0 U235 ( .IN1(n365), .IN2(n252), .QN(n13) );
  NOR2X0 U236 ( .IN1(n11), .IN2(n12), .QN(n276) );
  NOR2X0 U237 ( .IN1(n271), .IN2(n272), .QN(n11) );
  NOR2X0 U238 ( .IN1(n691), .IN2(n690), .QN(n5) );
  NOR2X0 U239 ( .IN1(n606), .IN2(n605), .QN(n9) );
  NAND3X0 U240 ( .IN1(n492), .IN2(n399), .IN3(n463), .QN(n481) );
  OR2X1 U241 ( .IN1(n559), .IN2(n748), .Q(n780) );
  NOR2X0 U242 ( .IN1(n17), .IN2(n18), .QN(n211) );
  NOR2X0 U243 ( .IN1(n684), .IN2(n198), .QN(n17) );
  INVX0 U244 ( .INP(n370), .ZN(n19) );
  NOR4X0 U245 ( .IN1(n389), .IN2(n388), .IN3(n387), .IN4(n386), .QN(n689) );
  MUX21X1 U246 ( .IN1(add_result[1]), .IN2(sub_result[1]), .S(n501), .Q(n811)
         );
  INVX0 U247 ( .INP(input_factor_01[29]), .ZN(n599) );
  OA222X1 U248 ( .IN1(input_factor_02[29]), .IN2(n599), .IN3(n600), .IN4(
        input_factor_01[29]), .IN5(input_factor_01[23]), .IN6(n557), .Q(n29)
         );
  INVX0 U249 ( .INP(input_factor_01[25]), .ZN(n542) );
  INVX0 U250 ( .INP(n33), .ZN(n27) );
  NOR2X0 U251 ( .IN1(input_factor_02[25]), .IN2(n542), .QN(n38) );
  INVX0 U252 ( .INP(input_factor_02[28]), .ZN(n594) );
  INVX0 U253 ( .INP(input_factor_02[26]), .ZN(n582) );
  INVX0 U254 ( .INP(input_factor_01[28]), .ZN(n593) );
  INVX0 U255 ( .INP(input_factor_01[26]), .ZN(n581) );
  NAND4X0 U256 ( .IN1(n41), .IN2(n31), .IN3(n45), .IN4(n22), .QN(n26) );
  INVX0 U257 ( .INP(input_factor_01[27]), .ZN(n587) );
  INVX0 U258 ( .INP(input_factor_02[27]), .ZN(n588) );
  INVX0 U259 ( .INP(input_factor_01[24]), .ZN(n541) );
  NOR2X0 U260 ( .IN1(n541), .IN2(input_factor_02[24]), .QN(n36) );
  INVX0 U261 ( .INP(n36), .ZN(n23) );
  NAND4X0 U262 ( .IN1(n24), .IN2(n30), .IN3(n34), .IN4(n23), .QN(n25) );
  NOR4X0 U263 ( .IN1(n27), .IN2(n38), .IN3(n26), .IN4(n25), .QN(n28) );
  INVX0 U264 ( .INP(input_factor_01[30]), .ZN(n543) );
  INVX0 U265 ( .INP(n30), .ZN(n44) );
  INVX0 U266 ( .INP(n31), .ZN(n40) );
  INVX0 U267 ( .INP(n32), .ZN(n35) );
  OA221X1 U268 ( .IN1(n36), .IN2(n35), .IN3(n36), .IN4(n34), .IN5(n33), .Q(n37) );
  OA22X1 U269 ( .IN1(n38), .IN2(n37), .IN3(input_factor_01[26]), .IN4(n582), 
        .Q(n39) );
  OA22X1 U270 ( .IN1(n40), .IN2(n39), .IN3(input_factor_01[27]), .IN4(n588), 
        .Q(n43) );
  INVX0 U271 ( .INP(n41), .ZN(n42) );
  AO221X1 U272 ( .IN1(n45), .IN2(n44), .IN3(n45), .IN4(n43), .IN5(n42), .Q(n47) );
  AO221X1 U273 ( .IN1(n47), .IN2(n46), .IN3(n600), .IN4(input_factor_01[29]), 
        .IN5(input_factor_01[30]), .Q(n74) );
  INVX0 U274 ( .INP(input_factor_02[22]), .ZN(n702) );
  INVX0 U275 ( .INP(input_factor_02[21]), .ZN(n693) );
  INVX0 U276 ( .INP(input_factor_02[18]), .ZN(n678) );
  INVX0 U277 ( .INP(input_factor_02[17]), .ZN(n672) );
  INVX0 U278 ( .INP(input_factor_02[16]), .ZN(n666) );
  INVX0 U279 ( .INP(input_factor_02[15]), .ZN(n660) );
  INVX0 U280 ( .INP(input_factor_02[14]), .ZN(n654) );
  INVX0 U281 ( .INP(input_factor_02[13]), .ZN(n648) );
  INVX0 U282 ( .INP(input_factor_02[10]), .ZN(n633) );
  INVX0 U283 ( .INP(input_factor_02[9]), .ZN(n627) );
  INVX0 U284 ( .INP(input_factor_02[8]), .ZN(n623) );
  INVX0 U285 ( .INP(input_factor_02[7]), .ZN(n274) );
  INVX0 U286 ( .INP(input_factor_02[6]), .ZN(n254) );
  INVX0 U287 ( .INP(input_factor_02[5]), .ZN(n614) );
  INVX0 U288 ( .INP(input_factor_02[4]), .ZN(n220) );
  INVX0 U289 ( .INP(input_factor_02[3]), .ZN(n189) );
  INVX0 U290 ( .INP(input_factor_02[2]), .ZN(n160) );
  INVX0 U291 ( .INP(input_factor_02[0]), .ZN(n76) );
  AO21X1 U292 ( .IN1(input_factor_01[0]), .IN2(n76), .IN3(input_factor_01[1]), 
        .Q(n48) );
  AO222X1 U293 ( .IN1(input_factor_01[2]), .IN2(n160), .IN3(input_factor_01[2]), .IN4(n48), .IN5(n160), .IN6(n48), .Q(n49) );
  AO222X1 U294 ( .IN1(input_factor_01[3]), .IN2(n189), .IN3(input_factor_01[3]), .IN4(n49), .IN5(n189), .IN6(n49), .Q(n50) );
  AO222X1 U295 ( .IN1(input_factor_01[4]), .IN2(n220), .IN3(input_factor_01[4]), .IN4(n50), .IN5(n220), .IN6(n50), .Q(n51) );
  AO222X1 U296 ( .IN1(input_factor_01[5]), .IN2(n614), .IN3(input_factor_01[5]), .IN4(n51), .IN5(n614), .IN6(n51), .Q(n52) );
  AO222X1 U297 ( .IN1(input_factor_01[6]), .IN2(n254), .IN3(input_factor_01[6]), .IN4(n52), .IN5(n254), .IN6(n52), .Q(n53) );
  AO222X1 U298 ( .IN1(input_factor_01[7]), .IN2(n274), .IN3(input_factor_01[7]), .IN4(n53), .IN5(n274), .IN6(n53), .Q(n54) );
  AO222X1 U299 ( .IN1(input_factor_01[8]), .IN2(n623), .IN3(input_factor_01[8]), .IN4(n54), .IN5(n623), .IN6(n54), .Q(n55) );
  AO222X1 U300 ( .IN1(input_factor_01[9]), .IN2(n627), .IN3(input_factor_01[9]), .IN4(n55), .IN5(n627), .IN6(n55), .Q(n56) );
  AO222X1 U301 ( .IN1(input_factor_01[10]), .IN2(n633), .IN3(
        input_factor_01[10]), .IN4(n56), .IN5(n633), .IN6(n56), .Q(n58) );
  INVX0 U302 ( .INP(input_factor_01[11]), .ZN(n638) );
  INVX0 U303 ( .INP(input_factor_02[11]), .ZN(n639) );
  AO221X1 U304 ( .IN1(n58), .IN2(n57), .IN3(n639), .IN4(input_factor_01[11]), 
        .IN5(input_factor_01[12]), .Q(n59) );
  AO222X1 U305 ( .IN1(input_factor_01[13]), .IN2(n648), .IN3(
        input_factor_01[13]), .IN4(n59), .IN5(n648), .IN6(n59), .Q(n60) );
  AO222X1 U306 ( .IN1(input_factor_01[14]), .IN2(n654), .IN3(
        input_factor_01[14]), .IN4(n60), .IN5(n654), .IN6(n60), .Q(n61) );
  AO222X1 U307 ( .IN1(input_factor_01[15]), .IN2(n660), .IN3(
        input_factor_01[15]), .IN4(n61), .IN5(n660), .IN6(n61), .Q(n62) );
  AO222X1 U308 ( .IN1(input_factor_01[16]), .IN2(n666), .IN3(
        input_factor_01[16]), .IN4(n62), .IN5(n666), .IN6(n62), .Q(n63) );
  AO222X1 U309 ( .IN1(input_factor_01[17]), .IN2(n672), .IN3(
        input_factor_01[17]), .IN4(n63), .IN5(n672), .IN6(n63), .Q(n64) );
  AO222X1 U310 ( .IN1(input_factor_01[18]), .IN2(n678), .IN3(
        input_factor_01[18]), .IN4(n64), .IN5(n678), .IN6(n64), .Q(n66) );
  INVX0 U311 ( .INP(input_factor_01[19]), .ZN(n683) );
  INVX0 U312 ( .INP(input_factor_02[19]), .ZN(n684) );
  AO221X1 U313 ( .IN1(n66), .IN2(n65), .IN3(n684), .IN4(input_factor_01[19]), 
        .IN5(input_factor_01[20]), .Q(n67) );
  AO222X1 U314 ( .IN1(input_factor_01[21]), .IN2(n693), .IN3(
        input_factor_01[21]), .IN4(n67), .IN5(n693), .IN6(n67), .Q(n68) );
  AO222X1 U315 ( .IN1(input_factor_01[22]), .IN2(n702), .IN3(
        input_factor_01[22]), .IN4(n68), .IN5(n702), .IN6(n68), .Q(n69) );
  INVX0 U316 ( .INP(input_factor_01[1]), .ZN(n143) );
  NOR2X0 U317 ( .IN1(n390), .IN2(n143), .QN(N177) );
  INVX0 U318 ( .INP(input_factor_01[12]), .ZN(n644) );
  NOR2X0 U319 ( .IN1(n390), .IN2(n644), .QN(N188) );
  INVX0 U320 ( .INP(input_factor_01[20]), .ZN(n546) );
  NOR2X0 U321 ( .IN1(n390), .IN2(n546), .QN(N196) );
  AO22X1 U322 ( .IN1(input_factor_01[30]), .IN2(rst_n), .IN3(n844), .IN4(
        larger_exponent[7]), .Q(n822) );
  NOR2X0 U324 ( .IN1(n373), .IN2(n69), .QN(n308) );
  OA22X1 U325 ( .IN1(n678), .IN2(n196), .IN3(n672), .IN4(n197), .Q(n71) );
  NAND3X0 U326 ( .IN1(n19), .IN2(n147), .IN3(n120), .QN(n356) );
  MUX21X1 U327 ( .IN1(n211), .IN2(n356), .S(exp_diff_value[2]), .Q(n335) );
  AO22X1 U328 ( .IN1(input_factor_01[18]), .IN2(n193), .IN3(
        input_factor_01[16]), .IN4(n370), .Q(n73) );
  INVX0 U329 ( .INP(n198), .ZN(n192) );
  AO22X1 U330 ( .IN1(input_factor_01[19]), .IN2(n192), .IN3(
        input_factor_01[17]), .IN4(n185), .Q(n72) );
  NOR2X0 U331 ( .IN1(n73), .IN2(n72), .QN(n208) );
  INVX0 U332 ( .INP(input_factor_01[22]), .ZN(n699) );
  INVX0 U333 ( .INP(input_factor_01[21]), .ZN(n692) );
  AO222X1 U334 ( .IN1(n193), .IN2(n699), .IN3(n185), .IN4(n692), .IN5(n370), 
        .IN6(n546), .Q(n355) );
  MUX21X1 U335 ( .IN1(n208), .IN2(n355), .S(exp_diff_value[2]), .Q(n336) );
  INVX0 U336 ( .INP(n817), .ZN(n816) );
  OA22X1 U337 ( .IN1(n335), .IN2(n176), .IN3(n336), .IN4(n816), .Q(n77) );
  NOR3X0 U338 ( .IN1(exp_diff_value[5]), .IN2(exp_diff_value[6]), .IN3(
        exp_diff_value[7]), .QN(n75) );
  AND2X1 U339 ( .IN1(exp_diff_value[4]), .IN2(n75), .Q(n268) );
  OA22X1 U340 ( .IN1(n77), .IN2(n177), .IN3(n76), .IN4(n360), .Q(n118) );
  AO22X1 U341 ( .IN1(input_factor_01[10]), .IN2(n193), .IN3(input_factor_01[8]), .IN4(n370), .Q(n80) );
  AO22X1 U342 ( .IN1(input_factor_01[11]), .IN2(n192), .IN3(input_factor_01[9]), .IN4(n185), .Q(n79) );
  NOR2X0 U343 ( .IN1(n80), .IN2(n79), .QN(n210) );
  AO22X1 U344 ( .IN1(input_factor_01[14]), .IN2(n193), .IN3(
        input_factor_01[12]), .IN4(n370), .Q(n82) );
  AO22X1 U345 ( .IN1(input_factor_01[15]), .IN2(n192), .IN3(
        input_factor_01[13]), .IN4(n185), .Q(n81) );
  NOR2X0 U346 ( .IN1(n82), .IN2(n81), .QN(n209) );
  MUX21X1 U347 ( .IN1(n210), .IN2(n209), .S(exp_diff_value[2]), .Q(n283) );
  AO22X1 U348 ( .IN1(input_factor_01[2]), .IN2(n193), .IN3(input_factor_01[0]), 
        .IN4(n370), .Q(n84) );
  AO22X1 U349 ( .IN1(input_factor_01[3]), .IN2(n192), .IN3(input_factor_01[1]), 
        .IN4(n185), .Q(n83) );
  NOR2X0 U350 ( .IN1(n84), .IN2(n83), .QN(n87) );
  AO22X1 U351 ( .IN1(input_factor_01[6]), .IN2(n193), .IN3(input_factor_01[4]), 
        .IN4(n370), .Q(n86) );
  AO22X1 U352 ( .IN1(input_factor_01[7]), .IN2(n192), .IN3(input_factor_01[5]), 
        .IN4(n185), .Q(n85) );
  NOR2X0 U353 ( .IN1(n86), .IN2(n85), .QN(n216) );
  OA222X1 U354 ( .IN1(n4), .IN2(n283), .IN3(n275), .IN4(n87), .IN5(n214), 
        .IN6(n216), .Q(n116) );
  NOR4X0 U355 ( .IN1(exp_diff_value[4]), .IN2(exp_diff_value[5]), .IN3(
        exp_diff_value[6]), .IN4(exp_diff_value[7]), .QN(n372) );
  AO222X1 U356 ( .IN1(input_factor_02[0]), .IN2(n370), .IN3(input_factor_02[3]), .IN4(n192), .IN5(input_factor_02[2]), .IN6(n193), .Q(n92) );
  INVX0 U357 ( .INP(n275), .ZN(n371) );
  OA22X1 U358 ( .IN1(n633), .IN2(n196), .IN3(n623), .IN4(n19), .Q(n89) );
  OA22X1 U359 ( .IN1(n639), .IN2(n198), .IN3(n627), .IN4(n197), .Q(n88) );
  AO222X1 U360 ( .IN1(input_factor_02[15]), .IN2(n192), .IN3(
        input_factor_02[13]), .IN4(n185), .IN5(input_factor_02[14]), .IN6(n193), .Q(n213) );
  MUX21X1 U361 ( .IN1(n215), .IN2(n213), .S(exp_diff_value[2]), .Q(n281) );
  OA22X1 U362 ( .IN1(n254), .IN2(n196), .IN3(n220), .IN4(n19), .Q(n91) );
  OA22X1 U363 ( .IN1(n614), .IN2(n197), .IN3(n274), .IN4(n198), .Q(n90) );
  INVX0 U364 ( .INP(n214), .ZN(n207) );
  AOI222X1 U365 ( .IN1(n92), .IN2(n371), .IN3(exp_diff_value[3]), .IN4(n281), 
        .IN5(n217), .IN6(n207), .QN(n93) );
  OA22X1 U366 ( .IN1(n116), .IN2(n271), .IN3(n93), .IN4(n232), .Q(n117) );
  NAND3X0 U367 ( .IN1(n119), .IN2(n118), .IN3(n117), .QN(N152) );
  AO222X1 U368 ( .IN1(input_factor_02[18]), .IN2(n185), .IN3(
        input_factor_02[19]), .IN4(n193), .IN5(input_factor_02[17]), .IN6(n370), .Q(n229) );
  INVX0 U369 ( .INP(n229), .ZN(n121) );
  AOI22X1 U370 ( .IN1(input_factor_02[22]), .IN2(n185), .IN3(n3), .IN4(n120), 
        .QN(n358) );
  MUX21X1 U371 ( .IN1(n121), .IN2(n358), .S(exp_diff_value[2]), .Q(n339) );
  AO22X1 U372 ( .IN1(input_factor_01[19]), .IN2(n193), .IN3(
        input_factor_01[17]), .IN4(n370), .Q(n123) );
  AO22X1 U373 ( .IN1(input_factor_01[20]), .IN2(n192), .IN3(
        input_factor_01[18]), .IN4(n185), .Q(n122) );
  NOR2X0 U374 ( .IN1(n123), .IN2(n122), .QN(n226) );
  AO22X1 U375 ( .IN1(input_factor_01[22]), .IN2(n185), .IN3(
        input_factor_01[21]), .IN4(n3), .Q(n124) );
  NOR2X0 U376 ( .IN1(n193), .IN2(n124), .QN(n357) );
  MUX21X1 U377 ( .IN1(n226), .IN2(n357), .S(exp_diff_value[2]), .Q(n340) );
  OA22X1 U378 ( .IN1(n176), .IN2(n339), .IN3(n816), .IN4(n340), .Q(n132) );
  AO222X1 U379 ( .IN1(input_factor_02[10]), .IN2(n185), .IN3(
        input_factor_02[9]), .IN4(n370), .IN5(input_factor_02[11]), .IN6(n193), 
        .Q(n231) );
  OA22X1 U380 ( .IN1(n660), .IN2(n196), .IN3(n648), .IN4(n19), .Q(n126) );
  OA22X1 U381 ( .IN1(n654), .IN2(n197), .IN3(n666), .IN4(n198), .Q(n125) );
  MUX21X1 U382 ( .IN1(n231), .IN2(n230), .S(exp_diff_value[2]), .Q(n127) );
  INVX0 U383 ( .INP(n127), .ZN(n287) );
  OA222X1 U384 ( .IN1(n160), .IN2(n197), .IN3(n189), .IN4(n196), .IN5(n220), 
        .IN6(n198), .Q(n130) );
  AO22X1 U385 ( .IN1(input_factor_02[5]), .IN2(n370), .IN3(input_factor_02[7]), 
        .IN4(n193), .Q(n129) );
  AO22X1 U386 ( .IN1(input_factor_02[6]), .IN2(n185), .IN3(input_factor_02[8]), 
        .IN4(n192), .Q(n128) );
  NOR2X0 U387 ( .IN1(n129), .IN2(n128), .QN(n233) );
  OA222X1 U388 ( .IN1(n4), .IN2(n287), .IN3(n275), .IN4(n130), .IN5(n214), 
        .IN6(n233), .Q(n131) );
  OA22X1 U389 ( .IN1(n132), .IN2(n177), .IN3(n131), .IN4(n232), .Q(n146) );
  AO22X1 U390 ( .IN1(input_factor_01[11]), .IN2(n193), .IN3(input_factor_01[9]), .IN4(n370), .Q(n134) );
  AO22X1 U391 ( .IN1(input_factor_01[12]), .IN2(n192), .IN3(
        input_factor_01[10]), .IN4(n185), .Q(n133) );
  NOR2X0 U392 ( .IN1(n134), .IN2(n133), .QN(n228) );
  AO22X1 U393 ( .IN1(input_factor_01[15]), .IN2(n193), .IN3(
        input_factor_01[13]), .IN4(n370), .Q(n136) );
  AO22X1 U394 ( .IN1(input_factor_01[16]), .IN2(n192), .IN3(
        input_factor_01[14]), .IN4(n185), .Q(n135) );
  NOR2X0 U395 ( .IN1(n136), .IN2(n135), .QN(n227) );
  MUX21X1 U396 ( .IN1(n228), .IN2(n227), .S(exp_diff_value[2]), .Q(n288) );
  AO22X1 U397 ( .IN1(input_factor_01[3]), .IN2(n193), .IN3(input_factor_01[1]), 
        .IN4(n370), .Q(n139) );
  AO22X1 U398 ( .IN1(input_factor_01[4]), .IN2(n192), .IN3(input_factor_01[2]), 
        .IN4(n185), .Q(n137) );
  NOR2X0 U399 ( .IN1(n139), .IN2(n137), .QN(n142) );
  AO22X1 U400 ( .IN1(input_factor_01[7]), .IN2(n193), .IN3(input_factor_01[5]), 
        .IN4(n370), .Q(n141) );
  AO22X1 U401 ( .IN1(input_factor_01[8]), .IN2(n192), .IN3(input_factor_01[6]), 
        .IN4(n185), .Q(n140) );
  NOR2X0 U402 ( .IN1(n141), .IN2(n140), .QN(n234) );
  OA222X1 U403 ( .IN1(n4), .IN2(n288), .IN3(n275), .IN4(n142), .IN5(n214), 
        .IN6(n234), .Q(n144) );
  OA22X1 U404 ( .IN1(n144), .IN2(n271), .IN3(n143), .IN4(n359), .Q(n145) );
  OA222X1 U405 ( .IN1(n693), .IN2(n198), .IN3(n678), .IN4(n19), .IN5(n684), 
        .IN6(n197), .Q(n244) );
  MUX21X1 U406 ( .IN1(n244), .IN2(n367), .S(exp_diff_value[2]), .Q(n343) );
  AO22X1 U407 ( .IN1(input_factor_01[20]), .IN2(n193), .IN3(
        input_factor_01[18]), .IN4(n370), .Q(n149) );
  AO22X1 U408 ( .IN1(input_factor_01[21]), .IN2(n192), .IN3(
        input_factor_01[19]), .IN4(n185), .Q(n148) );
  NOR2X0 U409 ( .IN1(n149), .IN2(n148), .QN(n241) );
  AO21X1 U410 ( .IN1(n699), .IN2(n3), .IN3(exp_diff_value[1]), .Q(n365) );
  MUX21X1 U411 ( .IN1(n241), .IN2(n365), .S(exp_diff_value[2]), .Q(n344) );
  OA22X1 U412 ( .IN1(n343), .IN2(n176), .IN3(n344), .IN4(n816), .Q(n150) );
  OA22X1 U413 ( .IN1(n150), .IN2(n177), .IN3(n160), .IN4(n360), .Q(n171) );
  AO22X1 U414 ( .IN1(input_factor_01[12]), .IN2(n193), .IN3(
        input_factor_01[10]), .IN4(n370), .Q(n152) );
  AO22X1 U415 ( .IN1(input_factor_01[13]), .IN2(n192), .IN3(
        input_factor_01[11]), .IN4(n185), .Q(n151) );
  NOR2X0 U416 ( .IN1(n152), .IN2(n151), .QN(n243) );
  AO22X1 U417 ( .IN1(input_factor_01[16]), .IN2(n193), .IN3(
        input_factor_01[14]), .IN4(n370), .Q(n154) );
  AO22X1 U418 ( .IN1(input_factor_01[17]), .IN2(n192), .IN3(
        input_factor_01[15]), .IN4(n185), .Q(n153) );
  NOR2X0 U419 ( .IN1(n154), .IN2(n153), .QN(n242) );
  MUX21X1 U420 ( .IN1(n243), .IN2(n242), .S(exp_diff_value[2]), .Q(n294) );
  AO22X1 U421 ( .IN1(input_factor_01[4]), .IN2(n193), .IN3(input_factor_01[2]), 
        .IN4(n370), .Q(n156) );
  AO22X1 U422 ( .IN1(input_factor_01[5]), .IN2(n192), .IN3(input_factor_01[3]), 
        .IN4(n185), .Q(n155) );
  NOR2X0 U423 ( .IN1(n156), .IN2(n155), .QN(n159) );
  AO22X1 U424 ( .IN1(input_factor_01[8]), .IN2(n193), .IN3(input_factor_01[6]), 
        .IN4(n370), .Q(n158) );
  AO22X1 U425 ( .IN1(input_factor_01[9]), .IN2(n192), .IN3(input_factor_01[7]), 
        .IN4(n185), .Q(n157) );
  NOR2X0 U426 ( .IN1(n158), .IN2(n157), .QN(n249) );
  OA222X1 U427 ( .IN1(n4), .IN2(n294), .IN3(n275), .IN4(n159), .IN5(n214), 
        .IN6(n249), .Q(n169) );
  OA22X1 U428 ( .IN1(n160), .IN2(n19), .IN3(n220), .IN4(n196), .Q(n162) );
  OA22X1 U429 ( .IN1(n189), .IN2(n197), .IN3(n614), .IN4(n198), .Q(n161) );
  AO222X1 U430 ( .IN1(input_factor_02[10]), .IN2(n370), .IN3(
        input_factor_02[13]), .IN4(n192), .IN5(input_factor_02[11]), .IN6(n185), .Q(n247) );
  OA22X1 U431 ( .IN1(n654), .IN2(n19), .IN3(n666), .IN4(n196), .Q(n164) );
  OA22X1 U432 ( .IN1(n660), .IN2(n197), .IN3(n672), .IN4(n198), .Q(n163) );
  MUX21X1 U433 ( .IN1(n247), .IN2(n246), .S(exp_diff_value[2]), .Q(n292) );
  OA22X1 U434 ( .IN1(n254), .IN2(n19), .IN3(n623), .IN4(n196), .Q(n166) );
  OA22X1 U435 ( .IN1(n274), .IN2(n197), .IN3(n627), .IN4(n198), .Q(n165) );
  AOI222X1 U436 ( .IN1(n167), .IN2(n371), .IN3(exp_diff_value[3]), .IN4(n292), 
        .IN5(n250), .IN6(n207), .QN(n168) );
  OA22X1 U437 ( .IN1(n169), .IN2(n271), .IN3(n168), .IN4(n232), .Q(n170) );
  NAND3X0 U438 ( .IN1(n172), .IN2(n171), .IN3(n170), .QN(N154) );
  AO222X1 U439 ( .IN1(input_factor_02[21]), .IN2(n193), .IN3(
        input_factor_02[19]), .IN4(n370), .IN5(input_factor_02[22]), .IN6(n192), .Q(n264) );
  MUX21X1 U440 ( .IN1(n264), .IN2(n370), .S(exp_diff_value[2]), .Q(n173) );
  INVX0 U441 ( .INP(n173), .ZN(n348) );
  AO22X1 U442 ( .IN1(input_factor_01[21]), .IN2(n193), .IN3(
        input_factor_01[19]), .IN4(n370), .Q(n175) );
  AO22X1 U443 ( .IN1(input_factor_01[22]), .IN2(n192), .IN3(
        input_factor_01[20]), .IN4(n185), .Q(n174) );
  NOR2X0 U444 ( .IN1(n175), .IN2(n174), .QN(n260) );
  MUX21X1 U445 ( .IN1(n260), .IN2(n19), .S(exp_diff_value[2]), .Q(n350) );
  OA22X1 U446 ( .IN1(n348), .IN2(n176), .IN3(n350), .IN4(n816), .Q(n178) );
  OA22X1 U447 ( .IN1(n178), .IN2(n177), .IN3(n189), .IN4(n360), .Q(n205) );
  AO22X1 U448 ( .IN1(input_factor_01[13]), .IN2(n193), .IN3(
        input_factor_01[11]), .IN4(n370), .Q(n180) );
  AO22X1 U449 ( .IN1(input_factor_01[14]), .IN2(n192), .IN3(
        input_factor_01[12]), .IN4(n185), .Q(n179) );
  NOR2X0 U450 ( .IN1(n180), .IN2(n179), .QN(n263) );
  AO22X1 U451 ( .IN1(input_factor_01[17]), .IN2(n193), .IN3(
        input_factor_01[15]), .IN4(n370), .Q(n182) );
  AO22X1 U452 ( .IN1(input_factor_01[18]), .IN2(n192), .IN3(
        input_factor_01[16]), .IN4(n185), .Q(n181) );
  NOR2X0 U453 ( .IN1(n182), .IN2(n181), .QN(n261) );
  MUX21X1 U454 ( .IN1(n263), .IN2(n261), .S(exp_diff_value[2]), .Q(n300) );
  AO22X1 U455 ( .IN1(input_factor_01[5]), .IN2(n193), .IN3(input_factor_01[3]), 
        .IN4(n370), .Q(n184) );
  AO22X1 U456 ( .IN1(input_factor_01[6]), .IN2(n192), .IN3(input_factor_01[4]), 
        .IN4(n185), .Q(n183) );
  NOR2X0 U457 ( .IN1(n184), .IN2(n183), .QN(n188) );
  AO22X1 U458 ( .IN1(input_factor_01[9]), .IN2(n193), .IN3(input_factor_01[7]), 
        .IN4(n370), .Q(n187) );
  AO22X1 U459 ( .IN1(input_factor_01[10]), .IN2(n192), .IN3(input_factor_01[8]), .IN4(n185), .Q(n186) );
  NOR2X0 U460 ( .IN1(n187), .IN2(n186), .QN(n272) );
  OA222X1 U461 ( .IN1(n4), .IN2(n300), .IN3(n275), .IN4(n188), .IN5(n214), 
        .IN6(n272), .Q(n203) );
  OA22X1 U462 ( .IN1(n189), .IN2(n19), .IN3(n614), .IN4(n196), .Q(n191) );
  OA22X1 U463 ( .IN1(n254), .IN2(n198), .IN3(n220), .IN4(n197), .Q(n190) );
  AO222X1 U464 ( .IN1(input_factor_02[11]), .IN2(n370), .IN3(
        input_factor_02[13]), .IN4(n193), .IN5(n192), .IN6(input_factor_02[14]), .Q(n266) );
  OA22X1 U465 ( .IN1(n660), .IN2(n19), .IN3(n672), .IN4(n196), .Q(n195) );
  OA22X1 U466 ( .IN1(n678), .IN2(n198), .IN3(n666), .IN4(n197), .Q(n194) );
  MUX21X1 U467 ( .IN1(n266), .IN2(n265), .S(exp_diff_value[2]), .Q(n298) );
  OA22X1 U468 ( .IN1(n274), .IN2(n19), .IN3(n627), .IN4(n196), .Q(n200) );
  OA22X1 U469 ( .IN1(n633), .IN2(n198), .IN3(n623), .IN4(n197), .Q(n199) );
  AOI222X1 U470 ( .IN1(n201), .IN2(n371), .IN3(exp_diff_value[3]), .IN4(n298), 
        .IN5(n269), .IN6(n207), .QN(n202) );
  OA22X1 U471 ( .IN1(n203), .IN2(n271), .IN3(n202), .IN4(n232), .Q(n204) );
  NAND3X0 U472 ( .IN1(n206), .IN2(n205), .IN3(n204), .QN(N155) );
  INVX0 U473 ( .INP(n271), .ZN(n354) );
  MUX21X1 U474 ( .IN1(n209), .IN2(n208), .S(exp_diff_value[2]), .Q(n305) );
  OA22X1 U475 ( .IN1(n210), .IN2(n262), .IN3(n305), .IN4(n330), .Q(n225) );
  INVX0 U476 ( .INP(n211), .ZN(n212) );
  MUX21X1 U477 ( .IN1(n213), .IN2(n212), .S(exp_diff_value[2]), .Q(n304) );
  NOR2X0 U478 ( .IN1(n4), .IN2(n232), .QN(n307) );
  NOR2X0 U479 ( .IN1(n214), .IN2(n232), .QN(n267) );
  AOI22X1 U480 ( .IN1(n304), .IN2(n307), .IN3(n267), .IN4(n215), .QN(n224) );
  OA22X1 U481 ( .IN1(n216), .IN2(n271), .IN3(n356), .IN4(n248), .Q(n219) );
  INVX0 U482 ( .INP(n232), .ZN(n353) );
  OA22X1 U483 ( .IN1(n221), .IN2(n275), .IN3(n220), .IN4(n360), .Q(n223) );
  NAND4X0 U484 ( .IN1(n225), .IN2(n224), .IN3(n223), .IN4(n222), .QN(N156) );
  MUX21X1 U485 ( .IN1(n227), .IN2(n226), .S(exp_diff_value[2]), .Q(n313) );
  OA22X1 U486 ( .IN1(n228), .IN2(n262), .IN3(n330), .IN4(n313), .Q(n240) );
  MUX21X1 U487 ( .IN1(n230), .IN2(n229), .S(exp_diff_value[2]), .Q(n312) );
  AOI22X1 U488 ( .IN1(n307), .IN2(n312), .IN3(n267), .IN4(n231), .QN(n239) );
  INVX0 U489 ( .INP(input_factor_01[5]), .ZN(n613) );
  OA22X1 U490 ( .IN1(n614), .IN2(n360), .IN3(n613), .IN4(n359), .Q(n238) );
  OA22X1 U491 ( .IN1(n234), .IN2(n271), .IN3(n233), .IN4(n232), .Q(n236) );
  OA22X1 U492 ( .IN1(n357), .IN2(n252), .IN3(n358), .IN4(n248), .Q(n235) );
  AO21X1 U493 ( .IN1(n236), .IN2(n235), .IN3(n275), .Q(n237) );
  NAND4X0 U494 ( .IN1(n240), .IN2(n239), .IN3(n238), .IN4(n237), .QN(N157) );
  MUX21X1 U495 ( .IN1(n242), .IN2(n241), .S(exp_diff_value[2]), .Q(n319) );
  OA22X1 U496 ( .IN1(n243), .IN2(n262), .IN3(n319), .IN4(n330), .Q(n259) );
  INVX0 U497 ( .INP(n244), .ZN(n245) );
  MUX21X1 U498 ( .IN1(n246), .IN2(n245), .S(exp_diff_value[2]), .Q(n318) );
  AOI22X1 U499 ( .IN1(n318), .IN2(n307), .IN3(n267), .IN4(n247), .QN(n258) );
  OA22X1 U500 ( .IN1(n249), .IN2(n271), .IN3(n367), .IN4(n248), .Q(n253) );
  OA22X1 U501 ( .IN1(n255), .IN2(n275), .IN3(n254), .IN4(n360), .Q(n257) );
  NAND4X0 U502 ( .IN1(n259), .IN2(n258), .IN3(n257), .IN4(n256), .QN(N158) );
  MUX21X1 U503 ( .IN1(n261), .IN2(n260), .S(exp_diff_value[2]), .Q(n327) );
  OA22X1 U504 ( .IN1(n263), .IN2(n262), .IN3(n327), .IN4(n330), .Q(n280) );
  MUX21X1 U505 ( .IN1(n265), .IN2(n264), .S(exp_diff_value[2]), .Q(n326) );
  AOI22X1 U506 ( .IN1(n326), .IN2(n307), .IN3(n267), .IN4(n266), .QN(n279) );
  NAND3X0 U507 ( .IN1(n268), .IN2(n370), .IN3(n373), .QN(n273) );
  OA22X1 U508 ( .IN1(n276), .IN2(n275), .IN3(n274), .IN4(n360), .Q(n278) );
  NAND4X0 U509 ( .IN1(n280), .IN2(n279), .IN3(n278), .IN4(n277), .QN(N159) );
  INVX0 U510 ( .INP(n307), .ZN(n329) );
  OA22X1 U511 ( .IN1(n336), .IN2(n330), .IN3(n335), .IN4(n329), .Q(n286) );
  INVX0 U512 ( .INP(n281), .ZN(n282) );
  OA22X1 U513 ( .IN1(n283), .IN2(n349), .IN3(n282), .IN4(n347), .Q(n285) );
  INVX0 U514 ( .INP(input_factor_01[8]), .ZN(n622) );
  OA22X1 U515 ( .IN1(n623), .IN2(n360), .IN3(n622), .IN4(n359), .Q(n284) );
  NAND3X0 U516 ( .IN1(n286), .IN2(n285), .IN3(n284), .QN(N160) );
  OA22X1 U517 ( .IN1(n329), .IN2(n339), .IN3(n330), .IN4(n340), .Q(n291) );
  OA22X1 U518 ( .IN1(n349), .IN2(n288), .IN3(n347), .IN4(n287), .Q(n290) );
  INVX0 U519 ( .INP(input_factor_01[9]), .ZN(n626) );
  OA22X1 U520 ( .IN1(n627), .IN2(n360), .IN3(n626), .IN4(n359), .Q(n289) );
  NAND3X0 U521 ( .IN1(n291), .IN2(n290), .IN3(n289), .QN(N161) );
  OA22X1 U522 ( .IN1(n344), .IN2(n330), .IN3(n343), .IN4(n329), .Q(n297) );
  INVX0 U523 ( .INP(n292), .ZN(n293) );
  OA22X1 U524 ( .IN1(n294), .IN2(n349), .IN3(n293), .IN4(n347), .Q(n296) );
  INVX0 U525 ( .INP(input_factor_01[10]), .ZN(n632) );
  OA22X1 U526 ( .IN1(n633), .IN2(n360), .IN3(n632), .IN4(n359), .Q(n295) );
  NAND3X0 U527 ( .IN1(n297), .IN2(n296), .IN3(n295), .QN(N162) );
  OA22X1 U528 ( .IN1(n350), .IN2(n330), .IN3(n348), .IN4(n329), .Q(n303) );
  INVX0 U529 ( .INP(n298), .ZN(n299) );
  OA22X1 U530 ( .IN1(n300), .IN2(n349), .IN3(n299), .IN4(n347), .Q(n302) );
  OA22X1 U531 ( .IN1(n639), .IN2(n360), .IN3(n638), .IN4(n359), .Q(n301) );
  NAND3X0 U532 ( .IN1(n303), .IN2(n302), .IN3(n301), .QN(N163) );
  INVX0 U533 ( .INP(n304), .ZN(n306) );
  OA22X1 U534 ( .IN1(n306), .IN2(n347), .IN3(n305), .IN4(n349), .Q(n311) );
  OR2X1 U535 ( .IN1(n330), .IN2(exp_diff_value[2]), .Q(n321) );
  OA22X1 U536 ( .IN1(n356), .IN2(n322), .IN3(n355), .IN4(n321), .Q(n310) );
  NAND3X0 U537 ( .IN1(n311), .IN2(n310), .IN3(n309), .QN(N164) );
  INVX0 U538 ( .INP(n312), .ZN(n314) );
  OA22X1 U539 ( .IN1(n314), .IN2(n347), .IN3(n313), .IN4(n349), .Q(n317) );
  OA22X1 U540 ( .IN1(n358), .IN2(n322), .IN3(n357), .IN4(n321), .Q(n316) );
  INVX0 U541 ( .INP(input_factor_01[13]), .ZN(n647) );
  OA22X1 U542 ( .IN1(n648), .IN2(n360), .IN3(n647), .IN4(n359), .Q(n315) );
  NAND3X0 U543 ( .IN1(n317), .IN2(n316), .IN3(n315), .QN(N165) );
  INVX0 U544 ( .INP(n318), .ZN(n320) );
  OA22X1 U545 ( .IN1(n320), .IN2(n347), .IN3(n319), .IN4(n349), .Q(n325) );
  OA22X1 U546 ( .IN1(n367), .IN2(n322), .IN3(n365), .IN4(n321), .Q(n324) );
  INVX0 U547 ( .INP(input_factor_01[14]), .ZN(n653) );
  OA22X1 U548 ( .IN1(n654), .IN2(n360), .IN3(n653), .IN4(n359), .Q(n323) );
  NAND3X0 U549 ( .IN1(n325), .IN2(n324), .IN3(n323), .QN(N166) );
  INVX0 U550 ( .INP(n326), .ZN(n328) );
  OA22X1 U551 ( .IN1(n328), .IN2(n347), .IN3(n327), .IN4(n349), .Q(n334) );
  INVX0 U552 ( .INP(input_factor_01[15]), .ZN(n659) );
  OA22X1 U553 ( .IN1(n660), .IN2(n360), .IN3(n659), .IN4(n359), .Q(n333) );
  NAND3X0 U554 ( .IN1(n331), .IN2(n1), .IN3(n370), .QN(n332) );
  NAND3X0 U555 ( .IN1(n334), .IN2(n333), .IN3(n332), .QN(N167) );
  OA22X1 U556 ( .IN1(n336), .IN2(n349), .IN3(n335), .IN4(n347), .Q(n338) );
  INVX0 U557 ( .INP(input_factor_01[16]), .ZN(n665) );
  OA22X1 U558 ( .IN1(n666), .IN2(n360), .IN3(n665), .IN4(n359), .Q(n337) );
  OA22X1 U559 ( .IN1(n349), .IN2(n340), .IN3(n347), .IN4(n339), .Q(n342) );
  INVX0 U560 ( .INP(input_factor_01[17]), .ZN(n671) );
  OA22X1 U561 ( .IN1(n672), .IN2(n360), .IN3(n671), .IN4(n359), .Q(n341) );
  OA22X1 U562 ( .IN1(n344), .IN2(n349), .IN3(n343), .IN4(n347), .Q(n346) );
  INVX0 U563 ( .INP(input_factor_01[18]), .ZN(n677) );
  OA22X1 U564 ( .IN1(n678), .IN2(n360), .IN3(n677), .IN4(n359), .Q(n345) );
  OA22X1 U565 ( .IN1(n350), .IN2(n349), .IN3(n348), .IN4(n347), .Q(n352) );
  OA22X1 U566 ( .IN1(n684), .IN2(n360), .IN3(n683), .IN4(n359), .Q(n351) );
  OAI222X1 U567 ( .IN1(n366), .IN2(n356), .IN3(n359), .IN4(n546), .IN5(n364), 
        .IN6(n355), .QN(N172) );
  OA22X1 U568 ( .IN1(n358), .IN2(n366), .IN3(n357), .IN4(n364), .Q(n362) );
  OA22X1 U569 ( .IN1(n693), .IN2(n360), .IN3(n692), .IN4(n359), .Q(n361) );
  NAND3X0 U570 ( .IN1(input_factor_01[22]), .IN2(input_factor_02[22]), .IN3(
        n363), .QN(n369) );
  OA22X1 U571 ( .IN1(n367), .IN2(n366), .IN3(n365), .IN4(n364), .Q(n368) );
  NAND3X0 U572 ( .IN1(n372), .IN2(n371), .IN3(n370), .QN(n374) );
  MUX21X1 U573 ( .IN1(input_factor_01[0]), .IN2(input_factor_02[0]), .S(n390), 
        .Q(N176) );
  MUX21X1 U574 ( .IN1(input_factor_01[2]), .IN2(input_factor_02[2]), .S(n390), 
        .Q(N178) );
  MUX21X1 U575 ( .IN1(input_factor_01[3]), .IN2(input_factor_02[3]), .S(n390), 
        .Q(N179) );
  MUX21X1 U576 ( .IN1(input_factor_01[4]), .IN2(input_factor_02[4]), .S(n390), 
        .Q(N180) );
  MUX21X1 U577 ( .IN1(input_factor_01[5]), .IN2(input_factor_02[5]), .S(n390), 
        .Q(N181) );
  MUX21X1 U578 ( .IN1(input_factor_01[6]), .IN2(input_factor_02[6]), .S(n390), 
        .Q(N182) );
  MUX21X1 U579 ( .IN1(input_factor_01[7]), .IN2(input_factor_02[7]), .S(n390), 
        .Q(N183) );
  MUX21X1 U580 ( .IN1(input_factor_01[8]), .IN2(input_factor_02[8]), .S(n390), 
        .Q(N184) );
  MUX21X1 U581 ( .IN1(input_factor_01[9]), .IN2(input_factor_02[9]), .S(n390), 
        .Q(N185) );
  MUX21X1 U582 ( .IN1(input_factor_01[10]), .IN2(input_factor_02[10]), .S(n390), .Q(N186) );
  MUX21X1 U583 ( .IN1(input_factor_01[11]), .IN2(input_factor_02[11]), .S(n390), .Q(N187) );
  MUX21X1 U584 ( .IN1(input_factor_01[13]), .IN2(input_factor_02[13]), .S(n390), .Q(N189) );
  MUX21X1 U585 ( .IN1(input_factor_01[14]), .IN2(input_factor_02[14]), .S(n390), .Q(N190) );
  MUX21X1 U586 ( .IN1(input_factor_01[15]), .IN2(input_factor_02[15]), .S(n390), .Q(N191) );
  MUX21X1 U587 ( .IN1(input_factor_01[16]), .IN2(input_factor_02[16]), .S(n390), .Q(N192) );
  MUX21X1 U588 ( .IN1(input_factor_01[17]), .IN2(input_factor_02[17]), .S(n390), .Q(N193) );
  MUX21X1 U589 ( .IN1(input_factor_01[18]), .IN2(input_factor_02[18]), .S(n390), .Q(N194) );
  MUX21X1 U590 ( .IN1(input_factor_01[19]), .IN2(input_factor_02[19]), .S(n390), .Q(N195) );
  MUX21X1 U591 ( .IN1(input_factor_01[21]), .IN2(input_factor_02[21]), .S(n390), .Q(N197) );
  MUX21X1 U592 ( .IN1(input_factor_01[22]), .IN2(input_factor_02[22]), .S(n390), .Q(N198) );
  MUX21X1 U593 ( .IN1(add_result[0]), .IN2(sub_result[0]), .S(n501), .Q(n813)
         );
  MUX21X1 U594 ( .IN1(add_result[2]), .IN2(sub_result[2]), .S(n501), .Q(n791)
         );
  MUX21X1 U595 ( .IN1(add_result[3]), .IN2(sub_result[3]), .S(n501), .Q(n783)
         );
  MUX21X1 U596 ( .IN1(add_result[4]), .IN2(sub_result[4]), .S(n501), .Q(n792)
         );
  MUX21X1 U597 ( .IN1(add_result[5]), .IN2(sub_result[5]), .S(n501), .Q(n784)
         );
  MUX21X1 U598 ( .IN1(add_result[6]), .IN2(sub_result[6]), .S(n501), .Q(n759)
         );
  MUX21X1 U599 ( .IN1(add_result[7]), .IN2(sub_result[7]), .S(n501), .Q(n751)
         );
  MUX21X1 U600 ( .IN1(add_result[9]), .IN2(sub_result[9]), .S(n501), .Q(n735)
         );
  MUX21X1 U601 ( .IN1(add_result[10]), .IN2(sub_result[10]), .S(n501), .Q(n727) );
  NOR4X0 U602 ( .IN1(n501), .IN2(add_result[14]), .IN3(add_result[15]), .IN4(
        add_result[13]), .QN(n510) );
  NOR4X0 U603 ( .IN1(sub_result[15]), .IN2(sub_result[14]), .IN3(
        sub_result[13]), .IN4(n21), .QN(n508) );
  NOR2X0 U604 ( .IN1(n510), .IN2(n508), .QN(n378) );
  MUX21X1 U605 ( .IN1(add_result[11]), .IN2(sub_result[11]), .S(n501), .Q(n719) );
  MUX21X1 U606 ( .IN1(add_result[16]), .IN2(sub_result[16]), .S(n20), .Q(n394)
         );
  MUX21X1 U607 ( .IN1(add_result[17]), .IN2(sub_result[17]), .S(n20), .Q(n463)
         );
  MUX21X1 U608 ( .IN1(add_result[20]), .IN2(sub_result[20]), .S(n20), .Q(n397)
         );
  INVX0 U609 ( .INP(n397), .ZN(n490) );
  MUX21X1 U610 ( .IN1(add_result[22]), .IN2(sub_result[22]), .S(n20), .Q(n398)
         );
  INVX0 U611 ( .INP(n398), .ZN(n375) );
  MUX21X1 U612 ( .IN1(add_result[23]), .IN2(sub_result[23]), .S(n20), .Q(n393)
         );
  MUX21X1 U613 ( .IN1(add_result[21]), .IN2(sub_result[21]), .S(n20), .Q(n400)
         );
  NOR2X0 U614 ( .IN1(n401), .IN2(n400), .QN(n402) );
  MUX21X1 U615 ( .IN1(add_result[19]), .IN2(sub_result[19]), .S(n20), .Q(n472)
         );
  NOR2X0 U616 ( .IN1(n376), .IN2(n472), .QN(n399) );
  MUX21X1 U617 ( .IN1(add_result[18]), .IN2(sub_result[18]), .S(n20), .Q(n396)
         );
  NOR2X0 U618 ( .IN1(n463), .IN2(n377), .QN(n395) );
  MUX21X1 U619 ( .IN1(add_result[12]), .IN2(sub_result[12]), .S(n20), .Q(n440)
         );
  NOR4X0 U620 ( .IN1(n378), .IN2(n719), .IN3(n562), .IN4(n440), .QN(n714) );
  MUX21X1 U621 ( .IN1(add_result[8]), .IN2(sub_result[8]), .S(n20), .Q(n743)
         );
  NOR3X0 U622 ( .IN1(n735), .IN2(n559), .IN3(n743), .QN(n515) );
  NOR2X0 U623 ( .IN1(n759), .IN2(n379), .QN(n514) );
  NOR2X0 U624 ( .IN1(n792), .IN2(n380), .QN(n522) );
  NOR2X0 U625 ( .IN1(n791), .IN2(n381), .QN(n516) );
  NAND3X0 U626 ( .IN1(n805), .IN2(n797), .IN3(n516), .QN(n560) );
  NAND4X0 U627 ( .IN1(n633), .IN2(n660), .IN3(n639), .IN4(n654), .QN(n389) );
  OR4X1 U628 ( .IN1(input_factor_02[31]), .IN2(input_factor_02[27]), .IN3(
        input_factor_02[24]), .IN4(input_factor_02[25]), .Q(n388) );
  NAND4X0 U629 ( .IN1(n600), .IN2(n557), .IN3(n594), .IN4(n582), .QN(n387) );
  NOR4X0 U630 ( .IN1(input_factor_02[16]), .IN2(input_factor_02[17]), .IN3(
        input_factor_02[19]), .IN4(input_factor_02[22]), .QN(n385) );
  NOR4X0 U631 ( .IN1(input_factor_02[0]), .IN2(input_factor_02[21]), .IN3(
        input_factor_02[13]), .IN4(input_factor_02[18]), .QN(n384) );
  NOR4X0 U632 ( .IN1(input_factor_02[5]), .IN2(input_factor_02[7]), .IN3(
        input_factor_02[8]), .IN4(input_factor_02[9]), .QN(n383) );
  NOR4X0 U633 ( .IN1(input_factor_02[2]), .IN2(input_factor_02[3]), .IN3(
        input_factor_02[6]), .IN4(input_factor_02[4]), .QN(n382) );
  NAND4X0 U634 ( .IN1(n385), .IN2(n384), .IN3(n383), .IN4(n382), .QN(n386) );
  AO222X1 U635 ( .IN1(input_factor_01[31]), .IN2(n689), .IN3(
        input_factor_01[31]), .IN4(n391), .IN5(n390), .IN6(input_factor_02[31]), .Q(n392) );
  AND2X1 U636 ( .IN1(n560), .IN2(n392), .Q(N211) );
  MUX21X1 U637 ( .IN1(n813), .IN2(n811), .S(add_sub_result_24_), .Q(N226) );
  MUX21X1 U638 ( .IN1(n811), .IN2(n791), .S(add_sub_result_24_), .Q(N227) );
  MUX21X1 U639 ( .IN1(n791), .IN2(n783), .S(add_sub_result_24_), .Q(N228) );
  MUX21X1 U640 ( .IN1(n783), .IN2(n792), .S(add_sub_result_24_), .Q(N229) );
  MUX21X1 U641 ( .IN1(n792), .IN2(n784), .S(add_sub_result_24_), .Q(N230) );
  MUX21X1 U642 ( .IN1(n784), .IN2(n759), .S(add_sub_result_24_), .Q(N231) );
  MUX21X1 U643 ( .IN1(n759), .IN2(n751), .S(add_sub_result_24_), .Q(N232) );
  MUX21X1 U644 ( .IN1(n751), .IN2(n743), .S(add_sub_result_24_), .Q(N233) );
  MUX21X1 U645 ( .IN1(n743), .IN2(n735), .S(add_sub_result_24_), .Q(N234) );
  MUX21X1 U646 ( .IN1(n735), .IN2(n727), .S(add_sub_result_24_), .Q(N235) );
  MUX21X1 U647 ( .IN1(n727), .IN2(n719), .S(add_sub_result_24_), .Q(N236) );
  MUX21X1 U648 ( .IN1(n719), .IN2(n440), .S(add_sub_result_24_), .Q(N237) );
  MUX21X1 U649 ( .IN1(add_result[13]), .IN2(sub_result[13]), .S(n20), .Q(n445)
         );
  MUX21X1 U650 ( .IN1(n440), .IN2(n445), .S(add_sub_result_24_), .Q(N238) );
  MUX21X1 U651 ( .IN1(add_result[14]), .IN2(sub_result[14]), .S(n20), .Q(n499)
         );
  MUX21X1 U652 ( .IN1(n445), .IN2(n499), .S(add_sub_result_24_), .Q(N239) );
  MUX21X1 U653 ( .IN1(add_result[15]), .IN2(sub_result[15]), .S(n20), .Q(n454)
         );
  MUX21X1 U654 ( .IN1(n499), .IN2(n454), .S(add_sub_result_24_), .Q(N240) );
  MUX21X1 U655 ( .IN1(n454), .IN2(n394), .S(add_sub_result_24_), .Q(N241) );
  MUX21X1 U656 ( .IN1(n394), .IN2(n463), .S(add_sub_result_24_), .Q(N242) );
  MUX21X1 U657 ( .IN1(n463), .IN2(n396), .S(add_sub_result_24_), .Q(N243) );
  MUX21X1 U658 ( .IN1(n396), .IN2(n472), .S(add_sub_result_24_), .Q(N244) );
  MUX21X1 U659 ( .IN1(n472), .IN2(n397), .S(add_sub_result_24_), .Q(N245) );
  MUX21X1 U660 ( .IN1(n397), .IN2(n400), .S(add_sub_result_24_), .Q(N246) );
  MUX21X1 U661 ( .IN1(n400), .IN2(n398), .S(add_sub_result_24_), .Q(N247) );
  MUX21X1 U662 ( .IN1(n398), .IN2(n393), .S(add_sub_result_24_), .Q(N248) );
  NAND4X0 U663 ( .IN1(n494), .IN2(n483), .IN3(n487), .IN4(n485), .QN(N256) );
  INVX0 U664 ( .INP(n400), .ZN(n486) );
  NOR2X0 U665 ( .IN1(n486), .IN2(n401), .QN(n417) );
  NAND4X0 U666 ( .IN1(n494), .IN2(n481), .IN3(n487), .IN4(n489), .QN(N257) );
  NAND3X0 U667 ( .IN1(n402), .IN2(n490), .IN3(n472), .QN(n491) );
  NAND4X0 U668 ( .IN1(n494), .IN2(n483), .IN3(n491), .IN4(n481), .QN(N258) );
  NOR2X0 U669 ( .IN1(n805), .IN2(n485), .QN(N260) );
  INVX0 U670 ( .INP(n485), .ZN(n419) );
  AO22X1 U671 ( .IN1(n419), .IN2(n811), .IN3(n417), .IN4(n813), .Q(N261) );
  INVX0 U672 ( .INP(n487), .ZN(n418) );
  AO222X1 U673 ( .IN1(n813), .IN2(n418), .IN3(n811), .IN4(n417), .IN5(n791), 
        .IN6(n419), .Q(N262) );
  OA22X1 U674 ( .IN1(n797), .IN2(n487), .IN3(n805), .IN4(n491), .Q(n404) );
  OA22X1 U675 ( .IN1(n803), .IN2(n489), .IN3(n801), .IN4(n485), .Q(n403) );
  OA22X1 U676 ( .IN1(n781), .IN2(n485), .IN3(n801), .IN4(n489), .Q(n407) );
  OA22X1 U677 ( .IN1(n797), .IN2(n491), .IN3(n805), .IN4(n483), .Q(n406) );
  NAND3X0 U678 ( .IN1(n407), .IN2(n406), .IN3(n405), .QN(N264) );
  OA22X1 U679 ( .IN1(n771), .IN2(n485), .IN3(n801), .IN4(n487), .Q(n411) );
  OA22X1 U680 ( .IN1(n803), .IN2(n491), .IN3(n797), .IN4(n483), .Q(n410) );
  INVX0 U681 ( .INP(n481), .ZN(n412) );
  NAND4X0 U682 ( .IN1(n411), .IN2(n410), .IN3(n409), .IN4(n408), .QN(N265) );
  OA22X1 U683 ( .IN1(n781), .IN2(n487), .IN3(n801), .IN4(n491), .Q(n416) );
  OA22X1 U684 ( .IN1(n772), .IN2(n485), .IN3(n771), .IN4(n489), .Q(n415) );
  OA22X1 U685 ( .IN1(n803), .IN2(n483), .IN3(n805), .IN4(n494), .Q(n414) );
  NAND4X0 U686 ( .IN1(n416), .IN2(n415), .IN3(n414), .IN4(n413), .QN(N266) );
  NOR4X0 U687 ( .IN1(n419), .IN2(n418), .IN3(n417), .IN4(N258), .QN(n561) );
  OA22X1 U688 ( .IN1(n803), .IN2(n481), .IN3(n801), .IN4(n483), .Q(n423) );
  OA22X1 U689 ( .IN1(n764), .IN2(n485), .IN3(n771), .IN4(n487), .Q(n422) );
  OA22X1 U690 ( .IN1(n772), .IN2(n489), .IN3(n781), .IN4(n491), .Q(n421) );
  OA22X1 U691 ( .IN1(n797), .IN2(n494), .IN3(n805), .IN4(n821), .Q(n420) );
  NAND4X0 U692 ( .IN1(n423), .IN2(n422), .IN3(n421), .IN4(n420), .QN(N267) );
  OA22X1 U693 ( .IN1(n781), .IN2(n483), .IN3(n801), .IN4(n481), .Q(n427) );
  OA22X1 U694 ( .IN1(n756), .IN2(n485), .IN3(n772), .IN4(n487), .Q(n426) );
  OA22X1 U695 ( .IN1(n764), .IN2(n489), .IN3(n771), .IN4(n491), .Q(n425) );
  OA22X1 U696 ( .IN1(n803), .IN2(n494), .IN3(n797), .IN4(n821), .Q(n424) );
  NAND4X0 U697 ( .IN1(n427), .IN2(n426), .IN3(n425), .IN4(n424), .QN(N268) );
  OA22X1 U698 ( .IN1(n771), .IN2(n483), .IN3(n781), .IN4(n481), .Q(n431) );
  OA22X1 U699 ( .IN1(n748), .IN2(n485), .IN3(n764), .IN4(n487), .Q(n430) );
  OA22X1 U700 ( .IN1(n756), .IN2(n489), .IN3(n772), .IN4(n491), .Q(n429) );
  OA22X1 U701 ( .IN1(n803), .IN2(n821), .IN3(n801), .IN4(n494), .Q(n428) );
  NAND4X0 U702 ( .IN1(n431), .IN2(n430), .IN3(n429), .IN4(n428), .QN(N269) );
  OA22X1 U703 ( .IN1(n772), .IN2(n483), .IN3(n771), .IN4(n481), .Q(n435) );
  OA22X1 U704 ( .IN1(n756), .IN2(n487), .IN3(n740), .IN4(n485), .Q(n434) );
  OA22X1 U705 ( .IN1(n748), .IN2(n489), .IN3(n764), .IN4(n491), .Q(n433) );
  OA22X1 U706 ( .IN1(n781), .IN2(n494), .IN3(n801), .IN4(n821), .Q(n432) );
  NAND4X0 U707 ( .IN1(n435), .IN2(n434), .IN3(n433), .IN4(n432), .QN(N270) );
  OA22X1 U708 ( .IN1(n764), .IN2(n483), .IN3(n772), .IN4(n481), .Q(n439) );
  OA22X1 U709 ( .IN1(n732), .IN2(n485), .IN3(n748), .IN4(n487), .Q(n438) );
  OA22X1 U710 ( .IN1(n756), .IN2(n491), .IN3(n740), .IN4(n489), .Q(n437) );
  OA22X1 U711 ( .IN1(n771), .IN2(n494), .IN3(n781), .IN4(n821), .Q(n436) );
  NAND4X0 U712 ( .IN1(n439), .IN2(n438), .IN3(n437), .IN4(n436), .QN(N271) );
  OA22X1 U713 ( .IN1(n756), .IN2(n483), .IN3(n764), .IN4(n481), .Q(n444) );
  OA22X1 U714 ( .IN1(n724), .IN2(n485), .IN3(n740), .IN4(n487), .Q(n443) );
  OA22X1 U715 ( .IN1(n732), .IN2(n489), .IN3(n748), .IN4(n491), .Q(n442) );
  OA22X1 U716 ( .IN1(n772), .IN2(n494), .IN3(n771), .IN4(n821), .Q(n441) );
  NAND4X0 U717 ( .IN1(n444), .IN2(n443), .IN3(n442), .IN4(n441), .QN(N272) );
  OA22X1 U718 ( .IN1(n756), .IN2(n481), .IN3(n748), .IN4(n483), .Q(n449) );
  OA22X1 U719 ( .IN1(n732), .IN2(n487), .IN3(n713), .IN4(n485), .Q(n448) );
  OA22X1 U720 ( .IN1(n724), .IN2(n489), .IN3(n740), .IN4(n491), .Q(n447) );
  OA22X1 U721 ( .IN1(n764), .IN2(n494), .IN3(n772), .IN4(n821), .Q(n446) );
  NAND4X0 U722 ( .IN1(n449), .IN2(n448), .IN3(n447), .IN4(n446), .QN(N273) );
  OA22X1 U723 ( .IN1(n740), .IN2(n483), .IN3(n748), .IN4(n481), .Q(n453) );
  INVX0 U724 ( .INP(n499), .ZN(n493) );
  OA22X1 U725 ( .IN1(n493), .IN2(n485), .IN3(n724), .IN4(n487), .Q(n452) );
  OA22X1 U726 ( .IN1(n732), .IN2(n491), .IN3(n713), .IN4(n489), .Q(n451) );
  OA22X1 U727 ( .IN1(n756), .IN2(n494), .IN3(n764), .IN4(n821), .Q(n450) );
  NAND4X0 U728 ( .IN1(n453), .IN2(n452), .IN3(n451), .IN4(n450), .QN(N274) );
  OA22X1 U729 ( .IN1(n732), .IN2(n483), .IN3(n740), .IN4(n481), .Q(n458) );
  OA22X1 U730 ( .IN1(n563), .IN2(n485), .IN3(n713), .IN4(n487), .Q(n457) );
  OA22X1 U731 ( .IN1(n493), .IN2(n489), .IN3(n724), .IN4(n491), .Q(n456) );
  OA22X1 U732 ( .IN1(n756), .IN2(n821), .IN3(n748), .IN4(n494), .Q(n455) );
  NAND4X0 U733 ( .IN1(n458), .IN2(n457), .IN3(n456), .IN4(n455), .QN(N275) );
  OA22X1 U734 ( .IN1(n724), .IN2(n483), .IN3(n732), .IN4(n481), .Q(n462) );
  OA22X1 U735 ( .IN1(n493), .IN2(n487), .IN3(n482), .IN4(n485), .Q(n461) );
  OA22X1 U736 ( .IN1(n563), .IN2(n489), .IN3(n713), .IN4(n491), .Q(n460) );
  OA22X1 U737 ( .IN1(n740), .IN2(n494), .IN3(n748), .IN4(n821), .Q(n459) );
  NAND4X0 U738 ( .IN1(n462), .IN2(n461), .IN3(n460), .IN4(n459), .QN(N276) );
  OA22X1 U739 ( .IN1(n724), .IN2(n481), .IN3(n713), .IN4(n483), .Q(n467) );
  INVX0 U740 ( .INP(n463), .ZN(n484) );
  OA22X1 U741 ( .IN1(n563), .IN2(n487), .IN3(n484), .IN4(n485), .Q(n466) );
  OA22X1 U742 ( .IN1(n493), .IN2(n491), .IN3(n482), .IN4(n489), .Q(n465) );
  OA22X1 U743 ( .IN1(n732), .IN2(n494), .IN3(n740), .IN4(n821), .Q(n464) );
  NAND4X0 U744 ( .IN1(n467), .IN2(n466), .IN3(n465), .IN4(n464), .QN(N277) );
  OA22X1 U745 ( .IN1(n493), .IN2(n483), .IN3(n713), .IN4(n481), .Q(n471) );
  OA22X1 U746 ( .IN1(n492), .IN2(n485), .IN3(n482), .IN4(n487), .Q(n470) );
  OA22X1 U747 ( .IN1(n563), .IN2(n491), .IN3(n484), .IN4(n489), .Q(n469) );
  OA22X1 U748 ( .IN1(n724), .IN2(n494), .IN3(n732), .IN4(n821), .Q(n468) );
  NAND4X0 U749 ( .IN1(n471), .IN2(n470), .IN3(n469), .IN4(n468), .QN(N278) );
  OA22X1 U750 ( .IN1(n563), .IN2(n483), .IN3(n493), .IN4(n481), .Q(n476) );
  INVX0 U751 ( .INP(n472), .ZN(n488) );
  OA22X1 U752 ( .IN1(n484), .IN2(n487), .IN3(n488), .IN4(n485), .Q(n475) );
  OA22X1 U753 ( .IN1(n492), .IN2(n489), .IN3(n482), .IN4(n491), .Q(n474) );
  OA22X1 U754 ( .IN1(n724), .IN2(n821), .IN3(n713), .IN4(n494), .Q(n473) );
  NAND4X0 U755 ( .IN1(n476), .IN2(n475), .IN3(n474), .IN4(n473), .QN(N279) );
  OA22X1 U756 ( .IN1(n563), .IN2(n481), .IN3(n482), .IN4(n483), .Q(n480) );
  OA22X1 U757 ( .IN1(n492), .IN2(n487), .IN3(n490), .IN4(n485), .Q(n479) );
  OA22X1 U758 ( .IN1(n484), .IN2(n491), .IN3(n488), .IN4(n489), .Q(n478) );
  OA22X1 U759 ( .IN1(n493), .IN2(n494), .IN3(n713), .IN4(n821), .Q(n477) );
  NAND4X0 U760 ( .IN1(n480), .IN2(n479), .IN3(n478), .IN4(n477), .QN(N280) );
  OA22X1 U761 ( .IN1(n484), .IN2(n483), .IN3(n482), .IN4(n481), .Q(n498) );
  OA22X1 U762 ( .IN1(n488), .IN2(n487), .IN3(n486), .IN4(n485), .Q(n497) );
  OA22X1 U763 ( .IN1(n492), .IN2(n491), .IN3(n490), .IN4(n489), .Q(n496) );
  OA22X1 U764 ( .IN1(n563), .IN2(n494), .IN3(n493), .IN4(n821), .Q(n495) );
  NAND4X0 U765 ( .IN1(n498), .IN2(n497), .IN3(n496), .IN4(n495), .QN(N281) );
  NAND3X0 U766 ( .IN1(n499), .IN2(n512), .IN3(n563), .QN(n712) );
  AO22X1 U767 ( .IN1(n510), .IN2(add_result[12]), .IN3(n508), .IN4(
        sub_result[12]), .Q(n500) );
  INVX0 U768 ( .INP(n712), .ZN(n506) );
  NOR3X0 U769 ( .IN1(n501), .IN2(add_result[14]), .IN3(add_result[15]), .QN(
        n503) );
  NOR3X0 U770 ( .IN1(sub_result[14]), .IN2(sub_result[15]), .IN3(n21), .QN(
        n502) );
  AO22X1 U771 ( .IN1(n503), .IN2(add_result[13]), .IN3(n502), .IN4(
        sub_result[13]), .Q(n504) );
  NOR2X0 U772 ( .IN1(n506), .IN2(n505), .QN(N308) );
  INVX0 U773 ( .INP(add_result[12]), .ZN(n509) );
  INVX0 U774 ( .INP(sub_result[12]), .ZN(n507) );
  AO22X1 U775 ( .IN1(n510), .IN2(n509), .IN3(n508), .IN4(n507), .Q(n511) );
  NAND3X0 U776 ( .IN1(n512), .IN2(n719), .IN3(n511), .QN(n806) );
  NAND4X0 U777 ( .IN1(N308), .IN2(n806), .IN3(n789), .IN4(n780), .QN(n773) );
  NAND4X0 U778 ( .IN1(n789), .IN2(n712), .IN3(n718), .IN4(n773), .QN(N306) );
  NAND4X0 U779 ( .IN1(n780), .IN2(n711), .IN3(n718), .IN4(n773), .QN(N307) );
  AO22X1 U780 ( .IN1(n698), .IN2(exponent_factor_12[0]), .IN3(n817), .IN4(
        exponent_factor_21[0]), .Q(N34) );
  NAND3X0 U781 ( .IN1(n801), .IN2(n522), .IN3(n791), .QN(n535) );
  NAND3X0 U782 ( .IN1(n771), .IN2(n514), .IN3(n792), .QN(n530) );
  NAND3X0 U783 ( .IN1(n764), .IN2(n515), .IN3(n759), .QN(n531) );
  NAND3X0 U784 ( .IN1(n803), .IN2(n797), .IN3(n801), .QN(n513) );
  AND2X1 U785 ( .IN1(n530), .IN2(n532), .Q(n517) );
  NAND4X0 U786 ( .IN1(n519), .IN2(n517), .IN3(n531), .IN4(n533), .QN(n518) );
  NAND4X0 U787 ( .IN1(n535), .IN2(n530), .IN3(n531), .IN4(n518), .QN(N346) );
  NAND3X0 U788 ( .IN1(n517), .IN2(n534), .IN3(n518), .QN(N347) );
  NOR2X0 U789 ( .IN1(n805), .IN2(n533), .QN(N349) );
  AO22X1 U790 ( .IN1(n698), .IN2(exponent_factor_12[1]), .IN3(n817), .IN4(
        exponent_factor_21[1]), .Q(N35) );
  OAI22X1 U791 ( .IN1(n797), .IN2(n533), .IN3(n805), .IN4(n531), .QN(N350) );
  OAI222X1 U792 ( .IN1(n532), .IN2(n805), .IN3(n531), .IN4(n797), .IN5(n533), 
        .IN6(n803), .QN(N351) );
  OA22X1 U793 ( .IN1(n803), .IN2(n531), .IN3(n801), .IN4(n533), .Q(n521) );
  OA22X1 U794 ( .IN1(n797), .IN2(n532), .IN3(n805), .IN4(n530), .Q(n520) );
  OA22X1 U795 ( .IN1(n781), .IN2(n533), .IN3(n801), .IN4(n531), .Q(n525) );
  OA22X1 U796 ( .IN1(n803), .IN2(n532), .IN3(n797), .IN4(n530), .Q(n524) );
  AND2X1 U797 ( .IN1(n522), .IN2(n783), .Q(n536) );
  NAND3X0 U798 ( .IN1(n525), .IN2(n524), .IN3(n523), .QN(N353) );
  OA22X1 U799 ( .IN1(n771), .IN2(n533), .IN3(n781), .IN4(n531), .Q(n529) );
  OA22X1 U800 ( .IN1(n803), .IN2(n530), .IN3(n805), .IN4(n535), .Q(n528) );
  OR2X1 U801 ( .IN1(n532), .IN2(n801), .Q(n526) );
  NAND4X0 U802 ( .IN1(n529), .IN2(n528), .IN3(n527), .IN4(n526), .QN(N354) );
  OA22X1 U803 ( .IN1(n771), .IN2(n531), .IN3(n801), .IN4(n530), .Q(n540) );
  OA22X1 U804 ( .IN1(n772), .IN2(n533), .IN3(n781), .IN4(n532), .Q(n539) );
  OA22X1 U805 ( .IN1(n797), .IN2(n535), .IN3(n805), .IN4(n534), .Q(n538) );
  NAND4X0 U806 ( .IN1(n540), .IN2(n539), .IN3(n538), .IN4(n537), .QN(N355) );
  AO22X1 U807 ( .IN1(n698), .IN2(exponent_factor_12[2]), .IN3(n817), .IN4(
        exponent_factor_21[2]), .Q(N36) );
  AO22X1 U808 ( .IN1(n698), .IN2(exponent_factor_12[3]), .IN3(n817), .IN4(
        exponent_factor_21[3]), .Q(N37) );
  AO22X1 U809 ( .IN1(n698), .IN2(exponent_factor_12[4]), .IN3(n817), .IN4(
        exponent_factor_21[4]), .Q(N38) );
  NAND4X0 U810 ( .IN1(n542), .IN2(n599), .IN3(n587), .IN4(n541), .QN(n545) );
  INVX0 U811 ( .INP(input_factor_01[23]), .ZN(n556) );
  NAND4X0 U812 ( .IN1(n543), .IN2(n556), .IN3(n593), .IN4(n581), .QN(n544) );
  NOR2X0 U813 ( .IN1(n545), .IN2(n544), .QN(n555) );
  NOR4X0 U814 ( .IN1(input_factor_01[7]), .IN2(input_factor_01[6]), .IN3(
        input_factor_01[5]), .IN4(input_factor_01[4]), .QN(n554) );
  NOR4X0 U815 ( .IN1(input_factor_01[3]), .IN2(input_factor_01[2]), .IN3(
        input_factor_01[1]), .IN4(input_factor_01[0]), .QN(n553) );
  NAND4X0 U816 ( .IN1(n699), .IN2(n692), .IN3(n546), .IN4(n683), .QN(n551) );
  NAND4X0 U817 ( .IN1(n547), .IN2(n677), .IN3(n671), .IN4(n665), .QN(n550) );
  NAND4X0 U818 ( .IN1(n659), .IN2(n653), .IN3(n647), .IN4(n644), .QN(n549) );
  NAND4X0 U819 ( .IN1(n638), .IN2(n632), .IN3(n626), .IN4(n622), .QN(n548) );
  NOR4X0 U820 ( .IN1(n551), .IN2(n550), .IN3(n549), .IN4(n548), .QN(n552) );
  NAND4X0 U821 ( .IN1(n555), .IN2(n554), .IN3(n553), .IN4(n552), .QN(n701) );
  OA22X1 U822 ( .IN1(n557), .IN2(n701), .IN3(n700), .IN4(n556), .Q(n572) );
  INVX0 U823 ( .INP(n773), .ZN(n558) );
  OA21X1 U824 ( .IN1(n756), .IN2(n559), .IN3(n558), .Q(n565) );
  NAND3X0 U825 ( .IN1(n560), .IN2(n700), .IN3(n701), .QN(n567) );
  OA21X1 U826 ( .IN1(n563), .IN2(n562), .IN3(n561), .Q(n564) );
  AOI22X1 U827 ( .IN1(n704), .IN2(add_output_exponent_w3[0]), .IN3(n703), 
        .IN4(add_output_exponent_w2[0]), .QN(n571) );
  INVX0 U828 ( .INP(n567), .ZN(n566) );
  AND4X1 U829 ( .IN1(n568), .IN2(n566), .IN3(n565), .IN4(n564), .Q(n705) );
  NAND4X0 U830 ( .IN1(n572), .IN2(n571), .IN3(n570), .IN4(n569), .QN(N380) );
  INVX0 U831 ( .INP(n701), .ZN(n619) );
  AOI22X1 U832 ( .IN1(input_factor_02[24]), .IN2(n619), .IN3(n689), .IN4(
        input_factor_01[24]), .QN(n576) );
  AOI22X1 U833 ( .IN1(n704), .IN2(add_output_exponent_w3[1]), .IN3(n703), 
        .IN4(add_output_exponent_w2[1]), .QN(n575) );
  NAND4X0 U834 ( .IN1(n576), .IN2(n575), .IN3(n574), .IN4(n573), .QN(N381) );
  AOI22X1 U835 ( .IN1(input_factor_02[25]), .IN2(n619), .IN3(n689), .IN4(
        input_factor_01[25]), .QN(n580) );
  AOI22X1 U836 ( .IN1(n704), .IN2(add_output_exponent_w3[2]), .IN3(n703), 
        .IN4(add_output_exponent_w2[2]), .QN(n579) );
  NAND4X0 U837 ( .IN1(n580), .IN2(n579), .IN3(n578), .IN4(n577), .QN(N382) );
  OA22X1 U838 ( .IN1(n582), .IN2(n701), .IN3(n700), .IN4(n581), .Q(n586) );
  AOI22X1 U839 ( .IN1(n704), .IN2(add_output_exponent_w3[3]), .IN3(n703), 
        .IN4(add_output_exponent_w2[3]), .QN(n585) );
  NAND4X0 U840 ( .IN1(n586), .IN2(n585), .IN3(n584), .IN4(n583), .QN(N383) );
  OA22X1 U841 ( .IN1(n588), .IN2(n701), .IN3(n700), .IN4(n587), .Q(n592) );
  AOI22X1 U842 ( .IN1(n704), .IN2(add_output_exponent_w3[4]), .IN3(n703), 
        .IN4(add_output_exponent_w2[4]), .QN(n591) );
  NAND4X0 U843 ( .IN1(n592), .IN2(n591), .IN3(n590), .IN4(n589), .QN(N384) );
  OA22X1 U844 ( .IN1(n594), .IN2(n701), .IN3(n700), .IN4(n593), .Q(n598) );
  AOI22X1 U845 ( .IN1(n704), .IN2(add_output_exponent_w3[5]), .IN3(n703), 
        .IN4(add_output_exponent_w2[5]), .QN(n597) );
  NAND4X0 U846 ( .IN1(n598), .IN2(n597), .IN3(n596), .IN4(n595), .QN(N385) );
  OA22X1 U847 ( .IN1(n600), .IN2(n701), .IN3(n700), .IN4(n599), .Q(n604) );
  AOI22X1 U848 ( .IN1(n704), .IN2(add_output_exponent_w3[6]), .IN3(n703), 
        .IN4(add_output_exponent_w2[6]), .QN(n603) );
  NAND4X0 U849 ( .IN1(n604), .IN2(n603), .IN3(n602), .IN4(n601), .QN(N386) );
  AO22X1 U851 ( .IN1(n689), .IN2(input_factor_01[30]), .IN3(n706), .IN4(
        add_output_exponent_w1[7]), .Q(n606) );
  AO22X1 U852 ( .IN1(n704), .IN2(add_output_exponent_w3[7]), .IN3(n703), .IN4(
        add_output_exponent_w2[7]), .Q(n605) );
  AO222X1 U853 ( .IN1(input_factor_02[0]), .IN2(n619), .IN3(input_factor_01[0]), .IN4(n689), .IN5(n706), .IN6(pre_sig_res_01[0]), .Q(N388) );
  AO222X1 U854 ( .IN1(n689), .IN2(input_factor_01[1]), .IN3(n703), .IN4(
        pre_sig_res_02[1]), .IN5(pre_sig_res_01[1]), .IN6(n706), .Q(N389) );
  AO22X1 U855 ( .IN1(n698), .IN2(exponent_factor_12[5]), .IN3(n817), .IN4(
        exponent_factor_21[5]), .Q(N39) );
  AOI22X1 U856 ( .IN1(n703), .IN2(pre_sig_res_02[2]), .IN3(n706), .IN4(
        pre_sig_res_01[2]), .QN(n608) );
  AOI22X1 U857 ( .IN1(input_factor_02[2]), .IN2(n619), .IN3(n689), .IN4(
        input_factor_01[2]), .QN(n607) );
  AOI22X1 U858 ( .IN1(n703), .IN2(pre_sig_res_02[3]), .IN3(n706), .IN4(
        pre_sig_res_01[3]), .QN(n610) );
  AOI22X1 U859 ( .IN1(input_factor_02[3]), .IN2(n619), .IN3(n689), .IN4(
        input_factor_01[3]), .QN(n609) );
  AOI22X1 U860 ( .IN1(n703), .IN2(pre_sig_res_02[4]), .IN3(n706), .IN4(
        pre_sig_res_01[4]), .QN(n612) );
  AOI22X1 U861 ( .IN1(input_factor_02[4]), .IN2(n619), .IN3(n689), .IN4(
        input_factor_01[4]), .QN(n611) );
  AOI22X1 U862 ( .IN1(n703), .IN2(pre_sig_res_02[5]), .IN3(n706), .IN4(
        pre_sig_res_01[5]), .QN(n616) );
  OA22X1 U863 ( .IN1(n614), .IN2(n701), .IN3(n700), .IN4(n613), .Q(n615) );
  AOI22X1 U864 ( .IN1(n703), .IN2(pre_sig_res_02[6]), .IN3(n706), .IN4(
        pre_sig_res_01[6]), .QN(n618) );
  AOI22X1 U865 ( .IN1(input_factor_02[6]), .IN2(n619), .IN3(n689), .IN4(
        input_factor_01[6]), .QN(n617) );
  AOI22X1 U866 ( .IN1(n703), .IN2(pre_sig_res_02[7]), .IN3(n706), .IN4(
        pre_sig_res_01[7]), .QN(n621) );
  AOI22X1 U867 ( .IN1(input_factor_02[7]), .IN2(n619), .IN3(n689), .IN4(
        input_factor_01[7]), .QN(n620) );
  AOI22X1 U868 ( .IN1(n703), .IN2(pre_sig_res_02[8]), .IN3(n706), .IN4(
        pre_sig_res_01[8]), .QN(n625) );
  OA22X1 U869 ( .IN1(n623), .IN2(n701), .IN3(n700), .IN4(n622), .Q(n624) );
  OA22X1 U870 ( .IN1(n627), .IN2(n701), .IN3(n700), .IN4(n626), .Q(n631) );
  NAND4X0 U871 ( .IN1(n631), .IN2(n630), .IN3(n629), .IN4(n628), .QN(N397) );
  OA22X1 U872 ( .IN1(n633), .IN2(n701), .IN3(n700), .IN4(n632), .Q(n637) );
  NAND4X0 U873 ( .IN1(n637), .IN2(n636), .IN3(n635), .IN4(n634), .QN(N398) );
  OA22X1 U874 ( .IN1(n639), .IN2(n701), .IN3(n700), .IN4(n638), .Q(n643) );
  NAND4X0 U875 ( .IN1(n643), .IN2(n642), .IN3(n641), .IN4(n640), .QN(N399) );
  AO22X1 U876 ( .IN1(n698), .IN2(exponent_factor_12[6]), .IN3(n817), .IN4(
        exponent_factor_21[6]), .Q(N40) );
  NOR2X0 U877 ( .IN1(n700), .IN2(n644), .QN(n646) );
  AO22X1 U878 ( .IN1(n704), .IN2(pre_sig_res_03[12]), .IN3(n703), .IN4(
        pre_sig_res_02[12]), .Q(n645) );
  OA22X1 U879 ( .IN1(n648), .IN2(n701), .IN3(n700), .IN4(n647), .Q(n652) );
  NAND4X0 U880 ( .IN1(n652), .IN2(n651), .IN3(n650), .IN4(n649), .QN(N401) );
  OA22X1 U881 ( .IN1(n654), .IN2(n701), .IN3(n700), .IN4(n653), .Q(n658) );
  NAND4X0 U882 ( .IN1(n658), .IN2(n657), .IN3(n656), .IN4(n655), .QN(N402) );
  OA22X1 U883 ( .IN1(n660), .IN2(n701), .IN3(n700), .IN4(n659), .Q(n664) );
  NAND4X0 U884 ( .IN1(n664), .IN2(n663), .IN3(n662), .IN4(n661), .QN(N403) );
  OA22X1 U885 ( .IN1(n666), .IN2(n701), .IN3(n700), .IN4(n665), .Q(n670) );
  AOI22X1 U886 ( .IN1(n704), .IN2(pre_sig_res_03[16]), .IN3(n703), .IN4(
        pre_sig_res_02[16]), .QN(n669) );
  NAND4X0 U887 ( .IN1(n670), .IN2(n669), .IN3(n668), .IN4(n667), .QN(N404) );
  OA22X1 U888 ( .IN1(n672), .IN2(n701), .IN3(n700), .IN4(n671), .Q(n676) );
  AOI22X1 U889 ( .IN1(n704), .IN2(pre_sig_res_03[17]), .IN3(n703), .IN4(
        pre_sig_res_02[17]), .QN(n675) );
  NAND4X0 U890 ( .IN1(n676), .IN2(n675), .IN3(n674), .IN4(n673), .QN(N405) );
  OA22X1 U891 ( .IN1(n678), .IN2(n701), .IN3(n700), .IN4(n677), .Q(n682) );
  AOI22X1 U892 ( .IN1(n704), .IN2(pre_sig_res_03[18]), .IN3(n703), .IN4(
        pre_sig_res_02[18]), .QN(n681) );
  NAND4X0 U893 ( .IN1(n682), .IN2(n681), .IN3(n680), .IN4(n679), .QN(N406) );
  OA22X1 U894 ( .IN1(n684), .IN2(n701), .IN3(n700), .IN4(n683), .Q(n688) );
  AOI22X1 U895 ( .IN1(n704), .IN2(pre_sig_res_03[19]), .IN3(n703), .IN4(
        pre_sig_res_02[19]), .QN(n687) );
  NAND4X0 U896 ( .IN1(n688), .IN2(n687), .IN3(n686), .IN4(n685), .QN(N407) );
  AO22X1 U897 ( .IN1(n689), .IN2(input_factor_01[20]), .IN3(n706), .IN4(
        pre_sig_res_01[20]), .Q(n691) );
  AO22X1 U898 ( .IN1(n704), .IN2(pre_sig_res_03[20]), .IN3(n703), .IN4(
        pre_sig_res_02[20]), .Q(n690) );
  OA22X1 U899 ( .IN1(n693), .IN2(n701), .IN3(n700), .IN4(n692), .Q(n697) );
  AOI22X1 U900 ( .IN1(n704), .IN2(pre_sig_res_03[21]), .IN3(n703), .IN4(
        pre_sig_res_02[21]), .QN(n696) );
  NAND4X0 U901 ( .IN1(n697), .IN2(n696), .IN3(n695), .IN4(n694), .QN(N409) );
  AO22X1 U902 ( .IN1(n698), .IN2(exponent_factor_12[7]), .IN3(n817), .IN4(
        exponent_factor_21[7]), .Q(N41) );
  OA22X1 U903 ( .IN1(n702), .IN2(n701), .IN3(n700), .IN4(n699), .Q(n710) );
  AOI22X1 U904 ( .IN1(n704), .IN2(pre_sig_res_03[22]), .IN3(n703), .IN4(
        pre_sig_res_02[22]), .QN(n709) );
  NAND4X0 U905 ( .IN1(n710), .IN2(n709), .IN3(n708), .IN4(n707), .QN(N410) );
  NOR2X0 U906 ( .IN1(n844), .IN2(n711), .QN(n812) );
  NOR2X0 U907 ( .IN1(n712), .IN2(n844), .QN(n814) );
  OA22X1 U908 ( .IN1(n724), .IN2(n802), .IN3(n713), .IN4(n800), .Q(n723) );
  OA22X1 U909 ( .IN1(n740), .IN2(n806), .IN3(n764), .IN4(n773), .Q(n717) );
  INVX0 U910 ( .INP(rst_n), .ZN(n815) );
  NAND3X0 U911 ( .IN1(n715), .IN2(n735), .IN3(n714), .QN(n716) );
  OA22X1 U912 ( .IN1(n844), .IN2(n717), .IN3(n815), .IN4(n716), .Q(n722) );
  NAND4X0 U913 ( .IN1(n723), .IN2(n722), .IN3(n721), .IN4(n720), .QN(n843) );
  OA22X1 U914 ( .IN1(n724), .IN2(n800), .IN3(n732), .IN4(n802), .Q(n731) );
  OA22X1 U915 ( .IN1(n764), .IN2(n780), .IN3(n772), .IN4(n773), .Q(n726) );
  OA22X1 U916 ( .IN1(n756), .IN2(n789), .IN3(n748), .IN4(n806), .Q(n725) );
  AO21X1 U917 ( .IN1(n726), .IN2(n725), .IN3(n844), .Q(n730) );
  NAND4X0 U918 ( .IN1(n731), .IN2(n730), .IN3(n729), .IN4(n728), .QN(n842) );
  OA22X1 U919 ( .IN1(n732), .IN2(n800), .IN3(n740), .IN4(n802), .Q(n739) );
  OA22X1 U920 ( .IN1(n772), .IN2(n780), .IN3(n771), .IN4(n773), .Q(n734) );
  OA22X1 U921 ( .IN1(n756), .IN2(n806), .IN3(n764), .IN4(n789), .Q(n733) );
  AO21X1 U922 ( .IN1(n734), .IN2(n733), .IN3(n844), .Q(n738) );
  NAND4X0 U923 ( .IN1(n739), .IN2(n738), .IN3(n737), .IN4(n736), .QN(n841) );
  OA22X1 U924 ( .IN1(n740), .IN2(n800), .IN3(n748), .IN4(n802), .Q(n747) );
  OA22X1 U925 ( .IN1(n771), .IN2(n780), .IN3(n781), .IN4(n773), .Q(n742) );
  OA22X1 U926 ( .IN1(n764), .IN2(n806), .IN3(n772), .IN4(n789), .Q(n741) );
  AO21X1 U927 ( .IN1(n742), .IN2(n741), .IN3(n844), .Q(n746) );
  NAND4X0 U928 ( .IN1(n747), .IN2(n746), .IN3(n745), .IN4(n744), .QN(n840) );
  OA22X1 U929 ( .IN1(n756), .IN2(n802), .IN3(n748), .IN4(n800), .Q(n755) );
  OA22X1 U930 ( .IN1(n781), .IN2(n780), .IN3(n801), .IN4(n773), .Q(n750) );
  OA22X1 U931 ( .IN1(n772), .IN2(n806), .IN3(n771), .IN4(n789), .Q(n749) );
  AO21X1 U932 ( .IN1(n750), .IN2(n749), .IN3(n844), .Q(n754) );
  NAND4X0 U933 ( .IN1(n755), .IN2(n754), .IN3(n753), .IN4(n752), .QN(n839) );
  OA22X1 U934 ( .IN1(n756), .IN2(n800), .IN3(n764), .IN4(n802), .Q(n763) );
  OA22X1 U935 ( .IN1(n803), .IN2(n773), .IN3(n801), .IN4(n780), .Q(n758) );
  OA22X1 U936 ( .IN1(n771), .IN2(n806), .IN3(n781), .IN4(n789), .Q(n757) );
  AO21X1 U937 ( .IN1(n758), .IN2(n757), .IN3(n844), .Q(n762) );
  NAND4X0 U938 ( .IN1(n763), .IN2(n762), .IN3(n761), .IN4(n760), .QN(n838) );
  OA22X1 U939 ( .IN1(n764), .IN2(n800), .IN3(n772), .IN4(n802), .Q(n770) );
  OA22X1 U940 ( .IN1(n803), .IN2(n780), .IN3(n797), .IN4(n773), .Q(n766) );
  OA22X1 U941 ( .IN1(n781), .IN2(n806), .IN3(n801), .IN4(n789), .Q(n765) );
  AO21X1 U942 ( .IN1(n766), .IN2(n765), .IN3(n844), .Q(n769) );
  NAND4X0 U943 ( .IN1(n770), .IN2(n769), .IN3(n768), .IN4(n767), .QN(n837) );
  OA22X1 U944 ( .IN1(n772), .IN2(n800), .IN3(n771), .IN4(n802), .Q(n779) );
  OA22X1 U945 ( .IN1(n797), .IN2(n780), .IN3(n805), .IN4(n773), .Q(n775) );
  OA22X1 U946 ( .IN1(n803), .IN2(n789), .IN3(n801), .IN4(n806), .Q(n774) );
  AO21X1 U947 ( .IN1(n775), .IN2(n774), .IN3(n844), .Q(n778) );
  NAND4X0 U948 ( .IN1(n779), .IN2(n778), .IN3(n777), .IN4(n776), .QN(n836) );
  OA222X1 U949 ( .IN1(n806), .IN2(n803), .IN3(n780), .IN4(n805), .IN5(n789), 
        .IN6(n797), .Q(n782) );
  OA22X1 U950 ( .IN1(n844), .IN2(n782), .IN3(n781), .IN4(n802), .Q(n788) );
  NAND4X0 U951 ( .IN1(n788), .IN2(n787), .IN3(n786), .IN4(n785), .QN(n835) );
  OA22X1 U952 ( .IN1(n797), .IN2(n806), .IN3(n805), .IN4(n789), .Q(n790) );
  OA22X1 U953 ( .IN1(n801), .IN2(n802), .IN3(n790), .IN4(n815), .Q(n796) );
  NAND4X0 U954 ( .IN1(n796), .IN2(n795), .IN3(n794), .IN4(n793), .QN(n834) );
  AOI22X1 U955 ( .IN1(pre_sig_res_03[11]), .IN2(n815), .IN3(n804), .IN4(n813), 
        .QN(n799) );
  OA22X1 U956 ( .IN1(n803), .IN2(n800), .IN3(n797), .IN4(n802), .Q(n798) );
  OA22X1 U957 ( .IN1(n803), .IN2(n802), .IN3(n801), .IN4(n800), .Q(n810) );
  OR3X1 U958 ( .IN1(n806), .IN2(n815), .IN3(n805), .Q(n808) );
  NAND4X0 U959 ( .IN1(n810), .IN2(n809), .IN3(n808), .IN4(n807), .QN(n832) );
  AO222X1 U960 ( .IN1(n813), .IN2(n812), .IN3(n811), .IN4(n814), .IN5(n815), 
        .IN6(pre_sig_res_03[10]), .Q(n831) );
  AO22X1 U961 ( .IN1(pre_sig_res_03[9]), .IN2(n815), .IN3(n814), .IN4(n813), 
        .Q(n830) );
  AO222X1 U962 ( .IN1(input_factor_02[23]), .IN2(n819), .IN3(
        input_factor_01[23]), .IN4(n818), .IN5(larger_exponent[0]), .IN6(n844), 
        .Q(n829) );
  AO222X1 U963 ( .IN1(input_factor_02[24]), .IN2(n819), .IN3(
        input_factor_01[24]), .IN4(n818), .IN5(n844), .IN6(larger_exponent[1]), 
        .Q(n828) );
  AO222X1 U964 ( .IN1(input_factor_02[25]), .IN2(n819), .IN3(
        input_factor_01[25]), .IN4(n818), .IN5(n844), .IN6(larger_exponent[2]), 
        .Q(n827) );
  AO222X1 U965 ( .IN1(input_factor_02[26]), .IN2(n819), .IN3(
        input_factor_01[26]), .IN4(n818), .IN5(n844), .IN6(larger_exponent[3]), 
        .Q(n826) );
  AO222X1 U966 ( .IN1(input_factor_02[27]), .IN2(n819), .IN3(
        input_factor_01[27]), .IN4(n818), .IN5(n844), .IN6(larger_exponent[4]), 
        .Q(n825) );
  AO222X1 U967 ( .IN1(input_factor_02[28]), .IN2(n819), .IN3(
        input_factor_01[28]), .IN4(n818), .IN5(n844), .IN6(larger_exponent[5]), 
        .Q(n824) );
  AO222X1 U968 ( .IN1(input_factor_02[29]), .IN2(n819), .IN3(
        input_factor_01[29]), .IN4(n818), .IN5(n844), .IN6(larger_exponent[6]), 
        .Q(n823) );
endmodule


module add_257 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_258 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_259 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_260 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_261 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_262 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_263 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_264 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_265 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_266 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_267 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_268 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_269 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_270 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_271 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_272 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_273 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_274 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_275 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_276 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_277 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_278 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_279 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_280 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(b), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(b), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module adder24_5 ( clk, rst_n, a, b, cin, out );
  input [23:0] a;
  input [23:0] b;
  output [24:0] out;
  input clk, rst_n, cin;
  wire   c_tmp;
  wire   [24:0] s;
  wire   [22:0] c;

  add_280 add_01 ( .s(s[0]), .a(a[0]), .b(b[0]), .ci(1'b0), .co(c[0]) );
  add_279 add_02 ( .s(s[1]), .a(a[1]), .b(b[1]), .ci(c[0]), .co(c[1]) );
  add_278 add_03 ( .s(s[2]), .a(a[2]), .b(b[2]), .ci(c[1]), .co(c[2]) );
  add_277 add_04 ( .s(s[3]), .a(a[3]), .b(b[3]), .ci(c[2]), .co(c[3]) );
  add_276 add_05 ( .s(s[4]), .a(a[4]), .b(b[4]), .ci(c[3]), .co(c[4]) );
  add_275 add_06 ( .s(s[5]), .a(a[5]), .b(b[5]), .ci(c[4]), .co(c[5]) );
  add_274 add_07 ( .s(s[6]), .a(a[6]), .b(b[6]), .ci(c[5]), .co(c[6]) );
  add_273 add_08 ( .s(s[7]), .a(a[7]), .b(b[7]), .ci(c[6]), .co(c[7]) );
  add_272 add_09 ( .s(s[8]), .a(a[8]), .b(b[8]), .ci(c[7]), .co(c[8]) );
  add_271 add_10 ( .s(s[9]), .a(a[9]), .b(b[9]), .ci(c[8]), .co(c[9]) );
  add_270 add_11 ( .s(s[10]), .a(a[10]), .b(b[10]), .ci(c[9]), .co(c[10]) );
  add_269 add_12 ( .s(s[11]), .a(a[11]), .b(b[11]), .ci(c_tmp), .co(c[11]) );
  add_268 add_13 ( .s(s[12]), .a(a[12]), .b(b[12]), .ci(c[11]), .co(c[12]) );
  add_267 add_14 ( .s(s[13]), .a(a[13]), .b(b[13]), .ci(c[12]), .co(c[13]) );
  add_266 add_15 ( .s(s[14]), .a(a[14]), .b(b[14]), .ci(c[13]), .co(c[14]) );
  add_265 add_16 ( .s(s[15]), .a(a[15]), .b(b[15]), .ci(c[14]), .co(c[15]) );
  add_264 add_17 ( .s(s[16]), .a(a[16]), .b(b[16]), .ci(c[15]), .co(c[16]) );
  add_263 add_18 ( .s(s[17]), .a(a[17]), .b(b[17]), .ci(c[16]), .co(c[17]) );
  add_262 add_19 ( .s(s[18]), .a(a[18]), .b(b[18]), .ci(c[17]), .co(c[18]) );
  add_261 add_20 ( .s(s[19]), .a(a[19]), .b(b[19]), .ci(c[18]), .co(c[19]) );
  add_260 add_21 ( .s(s[20]), .a(a[20]), .b(b[20]), .ci(c[19]), .co(c[20]) );
  add_259 add_22 ( .s(s[21]), .a(a[21]), .b(b[21]), .ci(c[20]), .co(c[21]) );
  add_258 add_23 ( .s(s[22]), .a(a[22]), .b(b[22]), .ci(c[21]), .co(c[22]) );
  add_257 add_24 ( .s(s[23]), .a(a[23]), .b(b[23]), .ci(c[22]), .co(s[24]) );
  DFFARX1 out_reg_10_ ( .D(s[10]), .CLK(clk), .RSTB(rst_n), .Q(out[10]) );
  DFFARX1 out_reg_9_ ( .D(s[9]), .CLK(clk), .RSTB(rst_n), .Q(out[9]) );
  DFFARX1 out_reg_8_ ( .D(s[8]), .CLK(clk), .RSTB(rst_n), .Q(out[8]) );
  DFFARX1 out_reg_7_ ( .D(s[7]), .CLK(clk), .RSTB(rst_n), .Q(out[7]) );
  DFFARX1 out_reg_6_ ( .D(s[6]), .CLK(clk), .RSTB(rst_n), .Q(out[6]) );
  DFFARX1 out_reg_5_ ( .D(s[5]), .CLK(clk), .RSTB(rst_n), .Q(out[5]) );
  DFFARX1 out_reg_4_ ( .D(s[4]), .CLK(clk), .RSTB(rst_n), .Q(out[4]) );
  DFFARX1 out_reg_3_ ( .D(s[3]), .CLK(clk), .RSTB(rst_n), .Q(out[3]) );
  DFFARX1 out_reg_2_ ( .D(s[2]), .CLK(clk), .RSTB(rst_n), .Q(out[2]) );
  DFFARX1 out_reg_1_ ( .D(s[1]), .CLK(clk), .RSTB(rst_n), .Q(out[1]) );
  DFFARX1 out_reg_0_ ( .D(s[0]), .CLK(clk), .RSTB(rst_n), .Q(out[0]) );
  DFFARX1 c_tmp_reg ( .D(c[10]), .CLK(clk), .RSTB(rst_n), .Q(c_tmp) );
  DFFARX1 out_reg_24_ ( .D(s[24]), .CLK(clk), .RSTB(rst_n), .Q(out[24]) );
  DFFARX1 out_reg_23_ ( .D(s[23]), .CLK(clk), .RSTB(rst_n), .Q(out[23]) );
  DFFARX1 out_reg_22_ ( .D(s[22]), .CLK(clk), .RSTB(rst_n), .Q(out[22]) );
  DFFARX1 out_reg_21_ ( .D(s[21]), .CLK(clk), .RSTB(rst_n), .Q(out[21]) );
  DFFARX1 out_reg_20_ ( .D(s[20]), .CLK(clk), .RSTB(rst_n), .Q(out[20]) );
  DFFARX1 out_reg_19_ ( .D(s[19]), .CLK(clk), .RSTB(rst_n), .Q(out[19]) );
  DFFARX1 out_reg_18_ ( .D(s[18]), .CLK(clk), .RSTB(rst_n), .Q(out[18]) );
  DFFARX1 out_reg_17_ ( .D(s[17]), .CLK(clk), .RSTB(rst_n), .Q(out[17]) );
  DFFARX1 out_reg_16_ ( .D(s[16]), .CLK(clk), .RSTB(rst_n), .Q(out[16]) );
  DFFARX1 out_reg_15_ ( .D(s[15]), .CLK(clk), .RSTB(rst_n), .Q(out[15]) );
  DFFARX1 out_reg_14_ ( .D(s[14]), .CLK(clk), .RSTB(rst_n), .Q(out[14]) );
  DFFARX1 out_reg_13_ ( .D(s[13]), .CLK(clk), .RSTB(rst_n), .Q(out[13]) );
  DFFARX1 out_reg_12_ ( .D(s[12]), .CLK(clk), .RSTB(rst_n), .Q(out[12]) );
  DFFARX1 out_reg_11_ ( .D(s[11]), .CLK(clk), .RSTB(rst_n), .Q(out[11]) );
endmodule


module add_281 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_282 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_283 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_284 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_285 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_286 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_287 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_288 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_289 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_290 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_291 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_292 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_293 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_294 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_295 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_296 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_297 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_298 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_299 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_300 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_301 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_302 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_303 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_304 ( s, a, ci, co, b_BAR );
  input a, ci, b_BAR;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(b_BAR), .IN2(n1), .QN(co) );
  INVX0 U2 ( .INP(a), .ZN(n1) );
  MUX21X1 U3 ( .IN1(a), .IN2(n1), .S(b_BAR), .Q(s) );
endmodule


module adder24_6 ( clk, rst_n, a, b, cin, out );
  input [23:0] a;
  input [23:0] b;
  output [24:0] out;
  input clk, rst_n, cin;
  wire   c_tmp, n_1_net_, n_2_net_, n_3_net_, n_4_net_, n_5_net_, n_6_net_,
         n_7_net_, n_8_net_, n_9_net_, n_10_net_, n_11_net_, n_12_net_,
         n_13_net_, n_14_net_, n_15_net_, n_16_net_, n_17_net_, n_18_net_,
         n_19_net_, n_20_net_, n_21_net_, n_22_net_, n_23_net_;
  wire   [24:0] s;
  wire   [23:0] c;

  add_304 add_01 ( .s(s[0]), .a(a[0]), .ci(1'b1), .co(c[0]), .b_BAR(b[0]) );
  add_303 add_02 ( .s(s[1]), .a(a[1]), .b(n_1_net_), .ci(c[0]), .co(c[1]) );
  add_302 add_03 ( .s(s[2]), .a(a[2]), .b(n_2_net_), .ci(c[1]), .co(c[2]) );
  add_301 add_04 ( .s(s[3]), .a(a[3]), .b(n_3_net_), .ci(c[2]), .co(c[3]) );
  add_300 add_05 ( .s(s[4]), .a(a[4]), .b(n_4_net_), .ci(c[3]), .co(c[4]) );
  add_299 add_06 ( .s(s[5]), .a(a[5]), .b(n_5_net_), .ci(c[4]), .co(c[5]) );
  add_298 add_07 ( .s(s[6]), .a(a[6]), .b(n_6_net_), .ci(c[5]), .co(c[6]) );
  add_297 add_08 ( .s(s[7]), .a(a[7]), .b(n_7_net_), .ci(c[6]), .co(c[7]) );
  add_296 add_09 ( .s(s[8]), .a(a[8]), .b(n_8_net_), .ci(c[7]), .co(c[8]) );
  add_295 add_10 ( .s(s[9]), .a(a[9]), .b(n_9_net_), .ci(c[8]), .co(c[9]) );
  add_294 add_11 ( .s(s[10]), .a(a[10]), .b(n_10_net_), .ci(c[9]), .co(c[10])
         );
  add_293 add_12 ( .s(s[11]), .a(a[11]), .b(n_11_net_), .ci(c_tmp), .co(c[11])
         );
  add_292 add_13 ( .s(s[12]), .a(a[12]), .b(n_12_net_), .ci(c[11]), .co(c[12])
         );
  add_291 add_14 ( .s(s[13]), .a(a[13]), .b(n_13_net_), .ci(c[12]), .co(c[13])
         );
  add_290 add_15 ( .s(s[14]), .a(a[14]), .b(n_14_net_), .ci(c[13]), .co(c[14])
         );
  add_289 add_16 ( .s(s[15]), .a(a[15]), .b(n_15_net_), .ci(c[14]), .co(c[15])
         );
  add_288 add_17 ( .s(s[16]), .a(a[16]), .b(n_16_net_), .ci(c[15]), .co(c[16])
         );
  add_287 add_18 ( .s(s[17]), .a(a[17]), .b(n_17_net_), .ci(c[16]), .co(c[17])
         );
  add_286 add_19 ( .s(s[18]), .a(a[18]), .b(n_18_net_), .ci(c[17]), .co(c[18])
         );
  add_285 add_20 ( .s(s[19]), .a(a[19]), .b(n_19_net_), .ci(c[18]), .co(c[19])
         );
  add_284 add_21 ( .s(s[20]), .a(a[20]), .b(n_20_net_), .ci(c[19]), .co(c[20])
         );
  add_283 add_22 ( .s(s[21]), .a(a[21]), .b(n_21_net_), .ci(c[20]), .co(c[21])
         );
  add_282 add_23 ( .s(s[22]), .a(a[22]), .b(n_22_net_), .ci(c[21]), .co(c[22])
         );
  add_281 add_24 ( .s(s[23]), .a(a[23]), .b(n_23_net_), .ci(c[22]), .co(c[23])
         );
  DFFARX1 out_reg_10_ ( .D(s[10]), .CLK(clk), .RSTB(rst_n), .Q(out[10]) );
  DFFARX1 out_reg_9_ ( .D(s[9]), .CLK(clk), .RSTB(rst_n), .Q(out[9]) );
  DFFARX1 out_reg_8_ ( .D(s[8]), .CLK(clk), .RSTB(rst_n), .Q(out[8]) );
  DFFARX1 out_reg_7_ ( .D(s[7]), .CLK(clk), .RSTB(rst_n), .Q(out[7]) );
  DFFARX1 out_reg_6_ ( .D(s[6]), .CLK(clk), .RSTB(rst_n), .Q(out[6]) );
  DFFARX1 out_reg_5_ ( .D(s[5]), .CLK(clk), .RSTB(rst_n), .Q(out[5]) );
  DFFARX1 out_reg_4_ ( .D(s[4]), .CLK(clk), .RSTB(rst_n), .Q(out[4]) );
  DFFARX1 out_reg_3_ ( .D(s[3]), .CLK(clk), .RSTB(rst_n), .Q(out[3]) );
  DFFARX1 out_reg_2_ ( .D(s[2]), .CLK(clk), .RSTB(rst_n), .Q(out[2]) );
  DFFARX1 out_reg_1_ ( .D(s[1]), .CLK(clk), .RSTB(rst_n), .Q(out[1]) );
  DFFARX1 out_reg_0_ ( .D(s[0]), .CLK(clk), .RSTB(rst_n), .Q(out[0]) );
  DFFARX1 c_tmp_reg ( .D(c[10]), .CLK(clk), .RSTB(rst_n), .Q(c_tmp) );
  DFFARX1 out_reg_24_ ( .D(s[24]), .CLK(clk), .RSTB(rst_n), .Q(out[24]) );
  DFFARX1 out_reg_23_ ( .D(s[23]), .CLK(clk), .RSTB(rst_n), .Q(out[23]) );
  DFFARX1 out_reg_22_ ( .D(s[22]), .CLK(clk), .RSTB(rst_n), .Q(out[22]) );
  DFFARX1 out_reg_21_ ( .D(s[21]), .CLK(clk), .RSTB(rst_n), .Q(out[21]) );
  DFFARX1 out_reg_20_ ( .D(s[20]), .CLK(clk), .RSTB(rst_n), .Q(out[20]) );
  DFFARX1 out_reg_19_ ( .D(s[19]), .CLK(clk), .RSTB(rst_n), .Q(out[19]) );
  DFFARX1 out_reg_18_ ( .D(s[18]), .CLK(clk), .RSTB(rst_n), .Q(out[18]) );
  DFFARX1 out_reg_17_ ( .D(s[17]), .CLK(clk), .RSTB(rst_n), .Q(out[17]) );
  DFFARX1 out_reg_16_ ( .D(s[16]), .CLK(clk), .RSTB(rst_n), .Q(out[16]) );
  DFFARX1 out_reg_15_ ( .D(s[15]), .CLK(clk), .RSTB(rst_n), .Q(out[15]) );
  DFFARX1 out_reg_14_ ( .D(s[14]), .CLK(clk), .RSTB(rst_n), .Q(out[14]) );
  DFFARX1 out_reg_13_ ( .D(s[13]), .CLK(clk), .RSTB(rst_n), .Q(out[13]) );
  DFFARX1 out_reg_12_ ( .D(s[12]), .CLK(clk), .RSTB(rst_n), .Q(out[12]) );
  DFFARX1 out_reg_11_ ( .D(s[11]), .CLK(clk), .RSTB(rst_n), .Q(out[11]) );
  INVX0 U3 ( .INP(b[1]), .ZN(n_1_net_) );
  INVX0 U4 ( .INP(b[2]), .ZN(n_2_net_) );
  INVX0 U5 ( .INP(b[3]), .ZN(n_3_net_) );
  INVX0 U6 ( .INP(b[4]), .ZN(n_4_net_) );
  INVX0 U7 ( .INP(b[5]), .ZN(n_5_net_) );
  INVX0 U8 ( .INP(b[6]), .ZN(n_6_net_) );
  INVX0 U9 ( .INP(b[7]), .ZN(n_7_net_) );
  INVX0 U10 ( .INP(b[8]), .ZN(n_8_net_) );
  INVX0 U11 ( .INP(b[9]), .ZN(n_9_net_) );
  INVX0 U12 ( .INP(b[10]), .ZN(n_10_net_) );
  INVX0 U13 ( .INP(c[23]), .ZN(s[24]) );
  INVX0 U14 ( .INP(b[11]), .ZN(n_11_net_) );
  INVX0 U15 ( .INP(b[12]), .ZN(n_12_net_) );
  INVX0 U16 ( .INP(b[13]), .ZN(n_13_net_) );
  INVX0 U17 ( .INP(b[14]), .ZN(n_14_net_) );
  INVX0 U18 ( .INP(b[15]), .ZN(n_15_net_) );
  INVX0 U19 ( .INP(b[16]), .ZN(n_16_net_) );
  INVX0 U20 ( .INP(b[17]), .ZN(n_17_net_) );
  INVX0 U21 ( .INP(b[18]), .ZN(n_18_net_) );
  INVX0 U22 ( .INP(b[19]), .ZN(n_19_net_) );
  INVX0 U23 ( .INP(b[20]), .ZN(n_20_net_) );
  INVX0 U24 ( .INP(b[21]), .ZN(n_21_net_) );
  INVX0 U25 ( .INP(b[22]), .ZN(n_22_net_) );
  INVX0 U26 ( .INP(b[23]), .ZN(n_23_net_) );
endmodule


module add_225 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  XNOR2X1 U1 ( .IN1(ci), .IN2(a), .Q(s) );
endmodule


module add_226 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_227 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_228 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_229 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_230 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_231 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_232 ( s, a, ci, co, b_BAR );
  input a, ci, b_BAR;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(b_BAR), .IN2(n1), .QN(co) );
  INVX0 U2 ( .INP(a), .ZN(n1) );
  MUX21X1 U3 ( .IN1(a), .IN2(n1), .S(b_BAR), .Q(s) );
endmodule


module adder8_17 ( out, a, b, cin );
  output [7:0] out;
  input [7:0] a;
  input [7:0] b;
  input cin;
  wire   n_1_net_, n_2_net_, n_4_net_;
  wire   [6:0] c;

  add_232 add_01 ( .s(out[0]), .a(a[0]), .ci(1'b1), .co(c[0]), .b_BAR(b[0]) );
  add_231 add_02 ( .s(out[1]), .a(a[1]), .b(n_1_net_), .ci(c[0]), .co(c[1]) );
  add_230 add_03 ( .s(out[2]), .a(a[2]), .b(n_2_net_), .ci(c[1]), .co(c[2]) );
  add_229 add_04 ( .s(out[3]), .a(a[3]), .b(1'b1), .ci(c[2]), .co(c[3]) );
  add_228 add_05 ( .s(out[4]), .a(a[4]), .b(n_4_net_), .ci(c[3]), .co(c[4]) );
  add_227 add_06 ( .s(out[5]), .a(a[5]), .b(1'b1), .ci(c[4]), .co(c[5]) );
  add_226 add_07 ( .s(out[6]), .a(a[6]), .b(1'b1), .ci(c[5]), .co(c[6]) );
  add_225 add_08 ( .s(out[7]), .a(a[7]), .b(1'b1), .ci(c[6]) );
  INVX0 U1 ( .INP(b[1]), .ZN(n_1_net_) );
  INVX0 U2 ( .INP(b[2]), .ZN(n_2_net_) );
  INVX0 U3 ( .INP(b[4]), .ZN(n_4_net_) );
endmodule


module add_233 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  XNOR2X1 U1 ( .IN1(ci), .IN2(a), .Q(s) );
endmodule


module add_234 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_235 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_236 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_237 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_238 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_239 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_240 ( s, a, ci, co, b_BAR );
  input a, ci, b_BAR;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(b_BAR), .IN2(n1), .QN(co) );
  INVX0 U2 ( .INP(a), .ZN(n1) );
  MUX21X1 U3 ( .IN1(a), .IN2(n1), .S(b_BAR), .Q(s) );
endmodule


module adder8_18 ( out, a, b, cin );
  output [7:0] out;
  input [7:0] a;
  input [7:0] b;
  input cin;
  wire   n_1_net_, n_2_net_, n_3_net_;
  wire   [6:0] c;

  add_240 add_01 ( .s(out[0]), .a(a[0]), .ci(1'b1), .co(c[0]), .b_BAR(b[0]) );
  add_239 add_02 ( .s(out[1]), .a(a[1]), .b(n_1_net_), .ci(c[0]), .co(c[1]) );
  add_238 add_03 ( .s(out[2]), .a(a[2]), .b(n_2_net_), .ci(c[1]), .co(c[2]) );
  add_237 add_04 ( .s(out[3]), .a(a[3]), .b(n_3_net_), .ci(c[2]), .co(c[3]) );
  add_236 add_05 ( .s(out[4]), .a(a[4]), .b(1'b1), .ci(c[3]), .co(c[4]) );
  add_235 add_06 ( .s(out[5]), .a(a[5]), .b(1'b1), .ci(c[4]), .co(c[5]) );
  add_234 add_07 ( .s(out[6]), .a(a[6]), .b(1'b1), .ci(c[5]), .co(c[6]) );
  add_233 add_08 ( .s(out[7]), .a(a[7]), .b(1'b1), .ci(c[6]) );
  INVX0 U1 ( .INP(b[1]), .ZN(n_1_net_) );
  INVX0 U2 ( .INP(b[2]), .ZN(n_2_net_) );
  INVX0 U3 ( .INP(b[3]), .ZN(n_3_net_) );
endmodule


module add_241 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  XNOR2X1 U1 ( .IN1(ci), .IN2(a), .Q(s) );
endmodule


module add_242 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_243 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_244 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(n1), .IN2(co), .QN(s) );
  NAND2X0 U2 ( .IN1(a), .IN2(ci), .QN(n1) );
  OR2X1 U3 ( .IN1(ci), .IN2(a), .Q(co) );
endmodule


module add_245 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_246 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_247 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_248 ( s, a, ci, co, b_BAR );
  input a, ci, b_BAR;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(b_BAR), .IN2(n1), .QN(co) );
  INVX0 U2 ( .INP(a), .ZN(n1) );
  MUX21X1 U3 ( .IN1(a), .IN2(n1), .S(b_BAR), .Q(s) );
endmodule


module adder8_19 ( out, a, b, cin );
  output [7:0] out;
  input [7:0] a;
  input [7:0] b;
  input cin;
  wire   n_1_net_, n_2_net_, n_3_net_;
  wire   [6:0] c;

  add_248 add_01 ( .s(out[0]), .a(a[0]), .ci(1'b1), .co(c[0]), .b_BAR(b[0]) );
  add_247 add_02 ( .s(out[1]), .a(a[1]), .b(n_1_net_), .ci(c[0]), .co(c[1]) );
  add_246 add_03 ( .s(out[2]), .a(a[2]), .b(n_2_net_), .ci(c[1]), .co(c[2]) );
  add_245 add_04 ( .s(out[3]), .a(a[3]), .b(n_3_net_), .ci(c[2]), .co(c[3]) );
  add_244 add_05 ( .s(out[4]), .a(a[4]), .b(1'b1), .ci(c[3]), .co(c[4]) );
  add_243 add_06 ( .s(out[5]), .a(a[5]), .b(1'b1), .ci(c[4]), .co(c[5]) );
  add_242 add_07 ( .s(out[6]), .a(a[6]), .b(1'b1), .ci(c[5]), .co(c[6]) );
  add_241 add_08 ( .s(out[7]), .a(a[7]), .b(1'b1), .ci(c[6]) );
  INVX0 U1 ( .INP(b[1]), .ZN(n_1_net_) );
  INVX0 U2 ( .INP(b[2]), .ZN(n_2_net_) );
  INVX0 U3 ( .INP(b[3]), .ZN(n_3_net_) );
endmodule


module add_249 ( s, a, b, co, ci_BAR );
  input a, b, ci_BAR;
  output s, co;


  XNOR2X1 U1 ( .IN1(a), .IN2(ci_BAR), .Q(s) );
endmodule


module add_250 ( s, a, b, ci, co_BAR );
  input a, b, ci;
  output s, co_BAR;


  NAND2X0 U1 ( .IN1(ci), .IN2(a), .QN(co_BAR) );
  OA21X1 U2 ( .IN1(ci), .IN2(a), .IN3(co_BAR), .Q(s) );
endmodule


module add_251 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_252 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_253 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_254 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_255 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_256 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(b), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(b), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module adder8_20 ( out, a, b, cin );
  output [7:0] out;
  input [7:0] a;
  input [7:0] b;
  input cin;

  wire   [6:0] c;

  add_256 add_01 ( .s(out[0]), .a(a[0]), .b(b[0]), .ci(1'b0), .co(c[0]) );
  add_255 add_02 ( .s(out[1]), .a(a[1]), .b(1'b0), .ci(c[0]), .co(c[1]) );
  add_254 add_03 ( .s(out[2]), .a(a[2]), .b(1'b0), .ci(c[1]), .co(c[2]) );
  add_253 add_04 ( .s(out[3]), .a(a[3]), .b(1'b0), .ci(c[2]), .co(c[3]) );
  add_252 add_05 ( .s(out[4]), .a(a[4]), .b(1'b0), .ci(c[3]), .co(c[4]) );
  add_251 add_06 ( .s(out[5]), .a(a[5]), .b(1'b0), .ci(c[4]), .co(c[5]) );
  add_250 add_07 ( .s(out[6]), .a(a[6]), .b(1'b0), .ci(c[5]), .co_BAR(c[6]) );
  add_249 add_08 ( .s(out[7]), .a(a[7]), .b(1'b0), .ci_BAR(c[6]) );
endmodule


module add_305 ( s, a, ci, co, b_BAR );
  input a, ci, b_BAR;
  output s, co;


  XNOR2X1 U1 ( .IN1(ci), .IN2(a), .Q(s) );
endmodule


module add_306 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_307 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_308 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_309 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_310 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_311 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_312 ( s, a, ci, co, b_BAR );
  input a, ci, b_BAR;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(b_BAR), .IN2(n1), .QN(co) );
  INVX0 U2 ( .INP(a), .ZN(n1) );
  MUX21X1 U3 ( .IN1(a), .IN2(n1), .S(b_BAR), .Q(s) );
endmodule


module adder8_21 ( out, a, b, cin );
  output [7:0] out;
  input [7:0] a;
  input [7:0] b;
  input cin;
  wire   n_1_net_, n_2_net_, n_3_net_, n_4_net_, n_5_net_, n_6_net_;
  wire   [6:0] c;

  add_312 add_01 ( .s(out[0]), .a(a[0]), .ci(1'b1), .co(c[0]), .b_BAR(b[0]) );
  add_311 add_02 ( .s(out[1]), .a(a[1]), .b(n_1_net_), .ci(c[0]), .co(c[1]) );
  add_310 add_03 ( .s(out[2]), .a(a[2]), .b(n_2_net_), .ci(c[1]), .co(c[2]) );
  add_309 add_04 ( .s(out[3]), .a(a[3]), .b(n_3_net_), .ci(c[2]), .co(c[3]) );
  add_308 add_05 ( .s(out[4]), .a(a[4]), .b(n_4_net_), .ci(c[3]), .co(c[4]) );
  add_307 add_06 ( .s(out[5]), .a(a[5]), .b(n_5_net_), .ci(c[4]), .co(c[5]) );
  add_306 add_07 ( .s(out[6]), .a(a[6]), .b(n_6_net_), .ci(c[5]), .co(c[6]) );
  add_305 add_08 ( .s(out[7]), .a(a[7]), .ci(c[6]), .b_BAR(1'b0) );
  INVX0 U1 ( .INP(b[1]), .ZN(n_1_net_) );
  INVX0 U2 ( .INP(b[2]), .ZN(n_2_net_) );
  INVX0 U3 ( .INP(b[3]), .ZN(n_3_net_) );
  INVX0 U4 ( .INP(b[4]), .ZN(n_4_net_) );
  INVX0 U5 ( .INP(b[5]), .ZN(n_5_net_) );
  INVX0 U6 ( .INP(b[6]), .ZN(n_6_net_) );
endmodule


module add_313 ( s, a, ci, co, b_BAR );
  input a, ci, b_BAR;
  output s, co;


  XNOR2X1 U1 ( .IN1(b_BAR), .IN2(ci), .Q(s) );
endmodule


module add_314 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_315 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_316 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_317 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_318 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_319 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_320 ( s, a, ci, co, b_BAR );
  input a, ci, b_BAR;
  output s, co;
  wire   n1;

  NAND2X0 U1 ( .IN1(b_BAR), .IN2(n1), .QN(co) );
  INVX0 U2 ( .INP(a), .ZN(n1) );
  MUX21X1 U3 ( .IN1(a), .IN2(n1), .S(b_BAR), .Q(s) );
endmodule


module adder8_22 ( out, a, b, cin );
  output [7:0] out;
  input [7:0] a;
  input [7:0] b;
  input cin;
  wire   n_1_net_, n_2_net_, n_3_net_, n_4_net_, n_5_net_, n_6_net_;
  wire   [6:0] c;

  add_320 add_01 ( .s(out[0]), .a(a[0]), .ci(1'b1), .co(c[0]), .b_BAR(b[0]) );
  add_319 add_02 ( .s(out[1]), .a(a[1]), .b(n_1_net_), .ci(c[0]), .co(c[1]) );
  add_318 add_03 ( .s(out[2]), .a(a[2]), .b(n_2_net_), .ci(c[1]), .co(c[2]) );
  add_317 add_04 ( .s(out[3]), .a(a[3]), .b(n_3_net_), .ci(c[2]), .co(c[3]) );
  add_316 add_05 ( .s(out[4]), .a(a[4]), .b(n_4_net_), .ci(c[3]), .co(c[4]) );
  add_315 add_06 ( .s(out[5]), .a(a[5]), .b(n_5_net_), .ci(c[4]), .co(c[5]) );
  add_314 add_07 ( .s(out[6]), .a(a[6]), .b(n_6_net_), .ci(c[5]), .co(c[6]) );
  add_313 add_08 ( .s(out[7]), .a(1'b0), .ci(c[6]), .b_BAR(b[7]) );
  INVX0 U1 ( .INP(b[1]), .ZN(n_1_net_) );
  INVX0 U2 ( .INP(b[2]), .ZN(n_2_net_) );
  INVX0 U3 ( .INP(b[3]), .ZN(n_3_net_) );
  INVX0 U4 ( .INP(b[4]), .ZN(n_4_net_) );
  INVX0 U5 ( .INP(b[5]), .ZN(n_5_net_) );
  INVX0 U6 ( .INP(b[6]), .ZN(n_6_net_) );
endmodule


module floating_point_adder_3 ( clk, rst_n, input_factor_01, input_factor_02, 
        output_adder );
  input [31:0] input_factor_01;
  input [31:0] input_factor_02;
  output [31:0] output_adder;
  input clk, rst_n;
  wire   N34, N35, N36, N37, N38, N39, N40, N41, N152, N153, N154, N155, N156,
         N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, N167,
         N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178,
         N179, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189,
         N190, N191, N192, N193, N194, N195, N196, N197, N198,
         add_sub_result_24_, N211, shift_temp_01_0_, N226, N227, N228, N229,
         N230, N231, N232, N233, N234, N235, N236, N237, N238, N239, N240,
         N241, N242, N243, N244, N245, N246, N247, N248, N256, N257, N258,
         N260, N261, N262, N263, N264, N265, N266, N267, N268, N269, N270,
         N271, N272, N273, N274, N275, N276, N277, N278, N279, N280, N281,
         N306, N307, N308, N346, N347, N348, N349, N350, N351, N352, N353,
         N354, N355, N380, N381, N382, N383, N384, N385, N386, N387, N388,
         N389, N390, N391, N392, N393, N394, N395, N396, N397, N398, N399,
         N400, N401, N402, N403, N404, N405, N406, N407, N408, N409, N410, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848;
  wire   [7:0] exp_diff_value;
  wire   [7:0] exponent_factor_21;
  wire   [7:0] exponent_factor_12;
  wire   [23:0] shift_smaller_factor;
  wire   [22:0] larger_factor;
  wire   [7:0] larger_exponent;
  wire   [24:0] add_result;
  wire   [24:0] sub_result;
  wire   [22:0] pre_sig_res_01;
  wire   [3:0] shift_temp_02;
  wire   [22:1] pre_sig_res_02;
  wire   [2:0] shift_temp_03;
  wire   [22:9] pre_sig_res_03;
  wire   [4:0] shift_temp_04;
  wire   [22:16] pre_sig_res_04;
  wire   [7:0] add_output_exponent_w1;
  wire   [7:0] add_output_exponent_w2;
  wire   [7:0] add_output_exponent_w3;
  wire   [7:0] add_output_exponent_w4;

  adder8_22 adder8_01 ( .out(exponent_factor_21), .a({1'b0, 
        input_factor_02[29:23]}), .b(input_factor_01[30:23]), .cin(1'b1) );
  adder8_21 adder8_02 ( .out(exponent_factor_12), .a(input_factor_01[30:23]), 
        .b({1'b0, input_factor_02[29:23]}), .cin(1'b1) );
  adder24_6 adder24_01 ( .clk(clk), .rst_n(rst_n), .a({shift_temp_04[4], 
        larger_factor}), .b(shift_smaller_factor), .cin(1'b1), .out(sub_result) );
  adder24_5 adder24_02 ( .clk(clk), .rst_n(rst_n), .a({shift_temp_04[4], 
        larger_factor}), .b(shift_smaller_factor), .cin(1'b0), .out(add_result) );
  adder8_20 adder8_03 ( .out(add_output_exponent_w1), .a(larger_exponent), .b(
        {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, shift_temp_01_0_}), .cin(
        1'b0) );
  adder8_19 adder8_04 ( .out(add_output_exponent_w2), .a(larger_exponent), .b(
        {1'b0, 1'b0, 1'b0, 1'b0, shift_temp_02}), .cin(1'b1) );
  adder8_18 adder8_05 ( .out(add_output_exponent_w3), .a(larger_exponent), .b(
        {1'b0, 1'b0, 1'b0, 1'b0, shift_temp_04[4], shift_temp_03}), .cin(1'b1)
         );
  adder8_17 adder8_06 ( .out(add_output_exponent_w4), .a(larger_exponent), .b(
        {1'b0, 1'b0, 1'b0, shift_temp_04[4], 1'b0, shift_temp_04[2:0]}), .cin(
        1'b1) );
  DFFARX1 exp_diff_value_reg_7_ ( .D(N41), .CLK(clk), .RSTB(rst_n), .Q(
        exp_diff_value[7]) );
  DFFARX1 exp_diff_value_reg_6_ ( .D(N40), .CLK(clk), .RSTB(rst_n), .Q(
        exp_diff_value[6]) );
  DFFARX1 exp_diff_value_reg_5_ ( .D(N39), .CLK(clk), .RSTB(rst_n), .Q(
        exp_diff_value[5]) );
  DFFARX1 exp_diff_value_reg_4_ ( .D(N38), .CLK(clk), .RSTB(rst_n), .Q(
        exp_diff_value[4]) );
  DFFARX1 exp_diff_value_reg_3_ ( .D(N37), .CLK(clk), .RSTB(rst_n), .Q(
        exp_diff_value[3]), .QN(n4) );
  DFFARX1 exp_diff_value_reg_2_ ( .D(N36), .CLK(clk), .RSTB(rst_n), .Q(n2), 
        .QN(n5) );
  DFFARX1 exp_diff_value_reg_1_ ( .D(N35), .CLK(clk), .RSTB(rst_n), .Q(
        exp_diff_value[1]), .QN(n3) );
  DFFARX1 exp_diff_value_reg_0_ ( .D(N34), .CLK(clk), .RSTB(rst_n), .Q(
        exp_diff_value[0]), .QN(n1) );
  DFFARX1 larger_factor_reg_22_ ( .D(N198), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[22]) );
  DFFARX1 larger_factor_reg_21_ ( .D(N197), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[21]) );
  DFFARX1 larger_factor_reg_20_ ( .D(N196), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[20]) );
  DFFARX1 larger_factor_reg_19_ ( .D(N195), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[19]) );
  DFFARX1 larger_factor_reg_18_ ( .D(N194), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[18]) );
  DFFARX1 larger_factor_reg_17_ ( .D(N193), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[17]) );
  DFFARX1 larger_factor_reg_16_ ( .D(N192), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[16]) );
  DFFARX1 larger_factor_reg_15_ ( .D(N191), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[15]) );
  DFFARX1 larger_factor_reg_14_ ( .D(N190), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[14]) );
  DFFARX1 larger_factor_reg_13_ ( .D(N189), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[13]) );
  DFFARX1 larger_factor_reg_12_ ( .D(N188), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[12]) );
  DFFARX1 larger_factor_reg_11_ ( .D(N187), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[11]) );
  DFFARX1 larger_factor_reg_10_ ( .D(N186), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[10]) );
  DFFARX1 larger_factor_reg_9_ ( .D(N185), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[9]) );
  DFFARX1 larger_factor_reg_8_ ( .D(N184), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[8]) );
  DFFARX1 larger_factor_reg_7_ ( .D(N183), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[7]) );
  DFFARX1 larger_factor_reg_6_ ( .D(N182), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[6]) );
  DFFARX1 larger_factor_reg_5_ ( .D(N181), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[5]) );
  DFFARX1 larger_factor_reg_4_ ( .D(N180), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[4]) );
  DFFARX1 larger_factor_reg_3_ ( .D(N179), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[3]) );
  DFFARX1 larger_factor_reg_2_ ( .D(N178), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[2]) );
  DFFARX1 larger_factor_reg_1_ ( .D(N177), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[1]) );
  DFFARX1 larger_factor_reg_0_ ( .D(N176), .CLK(clk), .RSTB(rst_n), .Q(
        larger_factor[0]) );
  DFFARX1 shift_smaller_factor_reg_23_ ( .D(N175), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[23]) );
  DFFARX1 shift_smaller_factor_reg_22_ ( .D(N174), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[22]) );
  DFFARX1 shift_smaller_factor_reg_21_ ( .D(N173), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[21]) );
  DFFARX1 shift_smaller_factor_reg_20_ ( .D(N172), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[20]) );
  DFFARX1 shift_smaller_factor_reg_19_ ( .D(N171), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[19]) );
  DFFARX1 shift_smaller_factor_reg_18_ ( .D(N170), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[18]) );
  DFFARX1 shift_smaller_factor_reg_17_ ( .D(N169), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[17]) );
  DFFARX1 shift_smaller_factor_reg_16_ ( .D(N168), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[16]) );
  DFFARX1 shift_smaller_factor_reg_15_ ( .D(N167), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[15]) );
  DFFARX1 shift_smaller_factor_reg_14_ ( .D(N166), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[14]) );
  DFFARX1 shift_smaller_factor_reg_13_ ( .D(N165), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[13]) );
  DFFARX1 shift_smaller_factor_reg_12_ ( .D(N164), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[12]) );
  DFFARX1 shift_smaller_factor_reg_11_ ( .D(N163), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[11]) );
  DFFARX1 shift_smaller_factor_reg_10_ ( .D(N162), .CLK(clk), .RSTB(rst_n), 
        .Q(shift_smaller_factor[10]) );
  DFFARX1 shift_smaller_factor_reg_9_ ( .D(N161), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[9]) );
  DFFARX1 shift_smaller_factor_reg_8_ ( .D(N160), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[8]) );
  DFFARX1 shift_smaller_factor_reg_7_ ( .D(N159), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[7]) );
  DFFARX1 shift_smaller_factor_reg_6_ ( .D(N158), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[6]) );
  DFFARX1 shift_smaller_factor_reg_5_ ( .D(N157), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[5]) );
  DFFARX1 shift_smaller_factor_reg_4_ ( .D(N156), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[4]) );
  DFFARX1 shift_smaller_factor_reg_3_ ( .D(N155), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[3]) );
  DFFARX1 shift_smaller_factor_reg_2_ ( .D(N154), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[2]) );
  DFFARX1 shift_smaller_factor_reg_1_ ( .D(N153), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[1]) );
  DFFARX1 shift_smaller_factor_reg_0_ ( .D(N152), .CLK(clk), .RSTB(rst_n), .Q(
        shift_smaller_factor[0]) );
  DFFX1 larger_exponent_reg_7_ ( .D(n826), .CLK(clk), .Q(larger_exponent[7])
         );
  DFFX1 larger_exponent_reg_6_ ( .D(n827), .CLK(clk), .Q(larger_exponent[6])
         );
  DFFX1 larger_exponent_reg_5_ ( .D(n828), .CLK(clk), .Q(larger_exponent[5])
         );
  DFFX1 larger_exponent_reg_4_ ( .D(n829), .CLK(clk), .Q(larger_exponent[4])
         );
  DFFX1 larger_exponent_reg_3_ ( .D(n830), .CLK(clk), .Q(larger_exponent[3])
         );
  DFFX1 larger_exponent_reg_2_ ( .D(n831), .CLK(clk), .Q(larger_exponent[2])
         );
  DFFX1 larger_exponent_reg_1_ ( .D(n832), .CLK(clk), .Q(larger_exponent[1])
         );
  DFFX1 larger_exponent_reg_0_ ( .D(n833), .CLK(clk), .Q(larger_exponent[0])
         );
  DFFARX1 shift_temp_04_reg_4_ ( .D(1'b1), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_04[4]) );
  DFFARX1 shift_temp_01_reg_0_ ( .D(add_sub_result_24_), .CLK(clk), .RSTB(
        rst_n), .Q(shift_temp_01_0_) );
  DFFARX1 pre_sig_res_02_reg_1_ ( .D(N260), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[1]) );
  DFFARX1 pre_sig_res_02_reg_2_ ( .D(N261), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[2]) );
  DFFARX1 pre_sig_res_02_reg_3_ ( .D(N262), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[3]) );
  DFFARX1 pre_sig_res_02_reg_4_ ( .D(N263), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[4]) );
  DFFARX1 pre_sig_res_02_reg_5_ ( .D(N264), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[5]) );
  DFFARX1 pre_sig_res_02_reg_6_ ( .D(N265), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[6]) );
  DFFARX1 pre_sig_res_02_reg_7_ ( .D(N266), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[7]) );
  DFFARX1 shift_temp_02_reg_2_ ( .D(N258), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_02[2]) );
  DFFASX1 shift_temp_02_reg_3_ ( .D(n825), .CLK(clk), .SETB(rst_n), .QN(
        shift_temp_02[3]) );
  DFFARX1 pre_sig_res_02_reg_8_ ( .D(N267), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[8]) );
  DFFARX1 pre_sig_res_02_reg_9_ ( .D(N268), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[9]) );
  DFFARX1 pre_sig_res_02_reg_10_ ( .D(N269), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[10]) );
  DFFARX1 pre_sig_res_02_reg_11_ ( .D(N270), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[11]) );
  DFFARX1 pre_sig_res_02_reg_12_ ( .D(N271), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[12]) );
  DFFARX1 pre_sig_res_02_reg_13_ ( .D(N272), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[13]) );
  DFFARX1 pre_sig_res_02_reg_14_ ( .D(N273), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[14]) );
  DFFARX1 pre_sig_res_02_reg_15_ ( .D(N274), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[15]) );
  DFFARX1 pre_sig_res_02_reg_16_ ( .D(N275), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[16]) );
  DFFARX1 pre_sig_res_02_reg_17_ ( .D(N276), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[17]) );
  DFFARX1 pre_sig_res_02_reg_18_ ( .D(N277), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[18]) );
  DFFARX1 pre_sig_res_02_reg_19_ ( .D(N278), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[19]) );
  DFFARX1 pre_sig_res_02_reg_20_ ( .D(N279), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[20]) );
  DFFARX1 pre_sig_res_02_reg_21_ ( .D(N280), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[21]) );
  DFFARX1 pre_sig_res_02_reg_22_ ( .D(N281), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_02[22]) );
  DFFARX1 shift_temp_02_reg_1_ ( .D(N257), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_02[1]) );
  DFFARX1 shift_temp_02_reg_0_ ( .D(N256), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_02[0]) );
  DFFX1 pre_sig_res_03_reg_9_ ( .D(n834), .CLK(clk), .Q(pre_sig_res_03[9]) );
  DFFX1 pre_sig_res_03_reg_10_ ( .D(n835), .CLK(clk), .Q(pre_sig_res_03[10])
         );
  DFFX1 pre_sig_res_03_reg_12_ ( .D(n836), .CLK(clk), .Q(pre_sig_res_03[12])
         );
  DFFX1 pre_sig_res_03_reg_11_ ( .D(n837), .CLK(clk), .Q(pre_sig_res_03[11])
         );
  DFFX1 pre_sig_res_03_reg_13_ ( .D(n838), .CLK(clk), .Q(pre_sig_res_03[13])
         );
  DFFX1 pre_sig_res_03_reg_14_ ( .D(n839), .CLK(clk), .Q(pre_sig_res_03[14])
         );
  DFFARX1 shift_temp_03_reg_2_ ( .D(N308), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_03[2]) );
  DFFARX1 shift_temp_03_reg_0_ ( .D(N306), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_03[0]) );
  DFFARX1 shift_temp_03_reg_1_ ( .D(N307), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_03[1]) );
  DFFX1 pre_sig_res_03_reg_15_ ( .D(n840), .CLK(clk), .Q(pre_sig_res_03[15])
         );
  DFFX1 pre_sig_res_03_reg_16_ ( .D(n841), .CLK(clk), .Q(pre_sig_res_03[16])
         );
  DFFX1 pre_sig_res_03_reg_17_ ( .D(n842), .CLK(clk), .Q(pre_sig_res_03[17])
         );
  DFFX1 pre_sig_res_03_reg_18_ ( .D(n843), .CLK(clk), .Q(pre_sig_res_03[18])
         );
  DFFX1 pre_sig_res_03_reg_19_ ( .D(n844), .CLK(clk), .Q(pre_sig_res_03[19])
         );
  DFFX1 pre_sig_res_03_reg_20_ ( .D(n845), .CLK(clk), .Q(pre_sig_res_03[20])
         );
  DFFX1 pre_sig_res_03_reg_21_ ( .D(n846), .CLK(clk), .Q(pre_sig_res_03[21])
         );
  DFFX1 pre_sig_res_03_reg_22_ ( .D(n847), .CLK(clk), .Q(pre_sig_res_03[22])
         );
  DFFARX1 pre_sig_res_04_reg_16_ ( .D(N349), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_04[16]) );
  DFFARX1 pre_sig_res_04_reg_17_ ( .D(N350), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_04[17]) );
  DFFARX1 pre_sig_res_04_reg_18_ ( .D(N351), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_04[18]) );
  DFFARX1 pre_sig_res_04_reg_19_ ( .D(N352), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_04[19]) );
  DFFARX1 pre_sig_res_04_reg_20_ ( .D(N353), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_04[20]) );
  DFFARX1 pre_sig_res_04_reg_21_ ( .D(N354), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_04[21]) );
  DFFARX1 pre_sig_res_04_reg_22_ ( .D(N355), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_04[22]) );
  DFFARX1 add_output_sign_reg ( .D(N211), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[31]) );
  DFFARX1 pre_sig_res_01_reg_0_ ( .D(N226), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[0]) );
  DFFARX1 pre_sig_res_01_reg_1_ ( .D(N227), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[1]) );
  DFFARX1 pre_sig_res_01_reg_2_ ( .D(N228), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[2]) );
  DFFARX1 pre_sig_res_01_reg_3_ ( .D(N229), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[3]) );
  DFFARX1 pre_sig_res_01_reg_4_ ( .D(N230), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[4]) );
  DFFARX1 pre_sig_res_01_reg_5_ ( .D(N231), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[5]) );
  DFFARX1 pre_sig_res_01_reg_6_ ( .D(N232), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[6]) );
  DFFARX1 pre_sig_res_01_reg_7_ ( .D(N233), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[7]) );
  DFFARX1 pre_sig_res_01_reg_8_ ( .D(N234), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[8]) );
  DFFARX1 pre_sig_res_01_reg_9_ ( .D(N235), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[9]) );
  DFFARX1 pre_sig_res_01_reg_10_ ( .D(N236), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[10]) );
  DFFARX1 pre_sig_res_01_reg_11_ ( .D(N237), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[11]) );
  DFFARX1 pre_sig_res_01_reg_12_ ( .D(N238), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[12]) );
  DFFARX1 pre_sig_res_01_reg_13_ ( .D(N239), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[13]) );
  DFFARX1 pre_sig_res_01_reg_14_ ( .D(N240), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[14]) );
  DFFARX1 pre_sig_res_01_reg_15_ ( .D(N241), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[15]) );
  DFFARX1 pre_sig_res_01_reg_16_ ( .D(N242), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[16]) );
  DFFARX1 pre_sig_res_01_reg_17_ ( .D(N243), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[17]) );
  DFFARX1 pre_sig_res_01_reg_18_ ( .D(N244), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[18]) );
  DFFARX1 pre_sig_res_01_reg_19_ ( .D(N245), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[19]) );
  DFFARX1 pre_sig_res_01_reg_20_ ( .D(N246), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[20]) );
  DFFARX1 pre_sig_res_01_reg_21_ ( .D(N247), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[21]) );
  DFFARX1 pre_sig_res_01_reg_22_ ( .D(N248), .CLK(clk), .RSTB(rst_n), .Q(
        pre_sig_res_01[22]) );
  DFFARX1 shift_temp_04_reg_2_ ( .D(N348), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_04[2]) );
  DFFARX1 shift_temp_04_reg_1_ ( .D(N347), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_04[1]) );
  DFFARX1 shift_temp_04_reg_0_ ( .D(N346), .CLK(clk), .RSTB(rst_n), .Q(
        shift_temp_04[0]) );
  DFFARX1 add_output_exponent_reg_7_ ( .D(N387), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[30]) );
  DFFARX1 add_output_exponent_reg_6_ ( .D(N386), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[29]) );
  DFFARX1 add_output_exponent_reg_5_ ( .D(N385), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[28]) );
  DFFARX1 add_output_exponent_reg_4_ ( .D(N384), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[27]) );
  DFFARX1 add_output_exponent_reg_3_ ( .D(N383), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[26]) );
  DFFARX1 add_output_exponent_reg_2_ ( .D(N382), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[25]) );
  DFFARX1 add_output_exponent_reg_1_ ( .D(N381), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[24]) );
  DFFARX1 add_output_exponent_reg_0_ ( .D(N380), .CLK(clk), .RSTB(rst_n), .Q(
        output_adder[23]) );
  DFFARX1 add_output_significands_reg_22_ ( .D(N410), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[22]) );
  DFFARX1 add_output_significands_reg_21_ ( .D(N409), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[21]) );
  DFFARX1 add_output_significands_reg_20_ ( .D(N408), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[20]) );
  DFFARX1 add_output_significands_reg_19_ ( .D(N407), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[19]) );
  DFFARX1 add_output_significands_reg_18_ ( .D(N406), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[18]) );
  DFFARX1 add_output_significands_reg_17_ ( .D(N405), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[17]) );
  DFFARX1 add_output_significands_reg_16_ ( .D(N404), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[16]) );
  DFFARX1 add_output_significands_reg_15_ ( .D(N403), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[15]) );
  DFFARX1 add_output_significands_reg_14_ ( .D(N402), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[14]) );
  DFFARX1 add_output_significands_reg_13_ ( .D(N401), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[13]) );
  DFFARX1 add_output_significands_reg_12_ ( .D(N400), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[12]) );
  DFFARX1 add_output_significands_reg_11_ ( .D(N399), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[11]) );
  DFFARX1 add_output_significands_reg_10_ ( .D(N398), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[10]) );
  DFFARX1 add_output_significands_reg_9_ ( .D(N397), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[9]) );
  DFFARX1 add_output_significands_reg_8_ ( .D(N396), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[8]) );
  DFFARX1 add_output_significands_reg_7_ ( .D(N395), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[7]) );
  DFFARX1 add_output_significands_reg_6_ ( .D(N394), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[6]) );
  DFFARX1 add_output_significands_reg_5_ ( .D(N393), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[5]) );
  DFFARX1 add_output_significands_reg_4_ ( .D(N392), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[4]) );
  DFFARX1 add_output_significands_reg_3_ ( .D(N391), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[3]) );
  DFFARX1 add_output_significands_reg_2_ ( .D(N390), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[2]) );
  DFFARX1 add_output_significands_reg_1_ ( .D(N389), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[1]) );
  DFFARX1 add_output_significands_reg_0_ ( .D(N388), .CLK(clk), .RSTB(rst_n), 
        .Q(output_adder[0]) );
  INVX1 U5 ( .INP(rst_n), .ZN(n848) );
  NAND2X0 U3 ( .IN1(n484), .IN2(n397), .QN(n559) );
  NAND2X0 U4 ( .IN1(exp_diff_value[4]), .IN2(n118), .QN(n212) );
  NAND2X0 U6 ( .IN1(input_factor_01[16]), .IN2(n372), .QN(n119) );
  NAND2X0 U7 ( .IN1(input_factor_02[17]), .IN2(n684), .QN(n67) );
  NAND2X0 U8 ( .IN1(n352), .IN2(n356), .QN(n545) );
  NAND2X0 U9 ( .IN1(input_factor_02[24]), .IN2(n543), .QN(n37) );
  NAND2X0 U10 ( .IN1(input_factor_01[27]), .IN2(n585), .QN(n33) );
  NAND2X0 U11 ( .IN1(input_factor_01[26]), .IN2(n579), .QN(n34) );
  NAND2X0 U12 ( .IN1(n23), .IN2(input_factor_02[25]), .QN(n36) );
  NAND2X0 U13 ( .IN1(input_factor_01[28]), .IN2(n591), .QN(n44) );
  NAND2X0 U14 ( .IN1(input_factor_02[28]), .IN2(n590), .QN(n48) );
  NAND2X0 U15 ( .IN1(n806), .IN2(n524), .QN(n382) );
  NAND2X0 U16 ( .IN1(n776), .IN2(n516), .QN(n381) );
  NAND2X0 U17 ( .IN1(n769), .IN2(n517), .QN(n380) );
  NAND2X0 U18 ( .IN1(n745), .IN2(n719), .QN(n556) );
  NAND2X0 U19 ( .IN1(n401), .IN2(n494), .QN(n378) );
  NAND2X0 U20 ( .IN1(n492), .IN2(n404), .QN(n377) );
  NAND2X0 U21 ( .IN1(n376), .IN2(n565), .QN(n403) );
  NAND2X0 U22 ( .IN1(n79), .IN2(n77), .QN(n218) );
  NAND2X0 U23 ( .IN1(n83), .IN2(n82), .QN(n219) );
  NAND2X0 U24 ( .IN1(n129), .IN2(n128), .QN(n240) );
  NAND2X0 U25 ( .IN1(n158), .IN2(n157), .QN(n249) );
  NAND2X0 U26 ( .IN1(n156), .IN2(n155), .QN(n250) );
  NAND2X0 U27 ( .IN1(n183), .IN2(n182), .QN(n269) );
  NAND2X0 U28 ( .IN1(exp_diff_value[1]), .IN2(exp_diff_value[0]), .QN(n184) );
  NAND2X0 U29 ( .IN1(n81), .IN2(n80), .QN(n226) );
  NAND2X0 U30 ( .IN1(n133), .IN2(n132), .QN(n236) );
  NAND2X0 U31 ( .IN1(n160), .IN2(n159), .QN(n257) );
  NAND2X0 U32 ( .IN1(n119), .IN2(n120), .QN(n19) );
  NAND2X0 U33 ( .IN1(input_factor_02[21]), .IN2(n700), .QN(n70) );
  NAND2X0 U34 ( .IN1(input_factor_02[27]), .IN2(n584), .QN(n26) );
  NAND2X0 U35 ( .IN1(input_factor_02[26]), .IN2(n578), .QN(n24) );
  NAND2X0 U36 ( .IN1(input_factor_01[23]), .IN2(n383), .QN(n35) );
  NAND2X0 U37 ( .IN1(n3), .IN2(n1), .QN(n207) );
  NAND2X0 U38 ( .IN1(n373), .IN2(n73), .QN(n72) );
  NAND2X0 U39 ( .IN1(n709), .IN2(pre_sig_res_01[9]), .QN(n640) );
  NAND2X0 U40 ( .IN1(n709), .IN2(pre_sig_res_01[10]), .QN(n646) );
  NAND2X0 U41 ( .IN1(n709), .IN2(pre_sig_res_01[11]), .QN(n652) );
  NAND2X0 U42 ( .IN1(n709), .IN2(pre_sig_res_01[12]), .QN(n658) );
  NAND2X0 U43 ( .IN1(n709), .IN2(pre_sig_res_01[13]), .QN(n664) );
  NAND2X0 U44 ( .IN1(n709), .IN2(pre_sig_res_01[14]), .QN(n670) );
  NAND2X0 U45 ( .IN1(n709), .IN2(pre_sig_res_01[15]), .QN(n676) );
  NAND2X0 U46 ( .IN1(n709), .IN2(pre_sig_res_01[16]), .QN(n680) );
  NAND2X0 U47 ( .IN1(n709), .IN2(pre_sig_res_01[17]), .QN(n686) );
  NAND2X0 U48 ( .IN1(n709), .IN2(pre_sig_res_01[20]), .QN(n696) );
  NAND2X0 U49 ( .IN1(n709), .IN2(pre_sig_res_01[21]), .QN(n704) );
  NAND2X0 U50 ( .IN1(n709), .IN2(add_output_exponent_w1[0]), .QN(n566) );
  NAND2X0 U51 ( .IN1(n709), .IN2(add_output_exponent_w1[1]), .QN(n570) );
  NAND2X0 U52 ( .IN1(n709), .IN2(add_output_exponent_w1[2]), .QN(n574) );
  NAND2X0 U53 ( .IN1(n709), .IN2(add_output_exponent_w1[3]), .QN(n580) );
  NAND2X0 U54 ( .IN1(n709), .IN2(add_output_exponent_w1[4]), .QN(n586) );
  NAND2X0 U55 ( .IN1(n709), .IN2(add_output_exponent_w1[5]), .QN(n592) );
  NAND2X0 U56 ( .IN1(n709), .IN2(add_output_exponent_w1[6]), .QN(n598) );
  NAND2X0 U57 ( .IN1(n518), .IN2(n816), .QN(n536) );
  NAND2X0 U58 ( .IN1(n515), .IN2(n524), .QN(n521) );
  NAND2X0 U59 ( .IN1(n72), .IN2(n367), .QN(n393) );
  NAND2X0 U60 ( .IN1(n516), .IN2(n789), .QN(n534) );
  NAND2X0 U61 ( .IN1(n517), .IN2(n756), .QN(n535) );
  NAND2X0 U62 ( .IN1(n761), .IN2(n745), .QN(n720) );
  NAND2X0 U63 ( .IN1(n719), .IN2(n732), .QN(n794) );
  NAND2X0 U64 ( .IN1(n514), .IN2(n502), .QN(n723) );
  NAND2X0 U65 ( .IN1(n514), .IN2(n506), .QN(n716) );
  NAND2X0 U66 ( .IN1(n397), .IN2(n396), .QN(n496) );
  NAND2X0 U67 ( .IN1(n414), .IN2(n818), .QN(n411) );
  NAND2X0 U68 ( .IN1(n401), .IN2(n398), .QN(n485) );
  NAND2X0 U69 ( .IN1(n404), .IN2(n399), .QN(n489) );
  NAND2X0 U70 ( .IN1(n400), .IN2(n565), .QN(n487) );
  NAND2X0 U71 ( .IN1(n76), .IN2(n75), .QN(n84) );
  NAND2X0 U72 ( .IN1(n135), .IN2(n134), .QN(n136) );
  NAND2X0 U73 ( .IN1(n162), .IN2(n161), .QN(n163) );
  NAND2X0 U74 ( .IN1(n708), .IN2(n370), .QN(n223) );
  NAND2X0 U75 ( .IN1(n370), .IN2(n821), .QN(n199) );
  NAND2X0 U76 ( .IN1(n186), .IN2(n185), .QN(n187) );
  NAND2X0 U77 ( .IN1(n708), .IN2(n122), .QN(n235) );
  NAND2X0 U78 ( .IN1(n821), .IN2(n122), .QN(n208) );
  NAND2X0 U79 ( .IN1(n220), .IN2(n222), .QN(n17) );
  NAND2X0 U80 ( .IN1(n280), .IN2(n240), .QN(n241) );
  NAND2X0 U81 ( .IN1(n131), .IN2(n130), .QN(n244) );
  NAND2X0 U82 ( .IN1(n821), .IN2(n266), .QN(n253) );
  NAND2X0 U83 ( .IN1(n708), .IN2(n266), .QN(n254) );
  NAND2X0 U84 ( .IN1(n271), .IN2(n272), .QN(n15) );
  NAND2X0 U85 ( .IN1(n270), .IN2(n269), .QN(n271) );
  NAND2X0 U86 ( .IN1(n181), .IN2(n180), .QN(n279) );
  NAND2X0 U87 ( .IN1(exp_diff_value[3]), .IN2(n216), .QN(n336) );
  NAND2X0 U88 ( .IN1(exp_diff_value[1]), .IN2(n1), .QN(n310) );
  NAND2X0 U89 ( .IN1(n323), .IN2(n5), .QN(n325) );
  NAND2X0 U90 ( .IN1(n337), .IN2(n336), .QN(n338) );
  NAND2X0 U91 ( .IN1(n4), .IN2(n216), .QN(n354) );
  NAND2X0 U92 ( .IN1(n311), .IN2(n310), .QN(n358) );
  NAND2X0 U93 ( .IN1(n74), .IN2(n123), .QN(n367) );
  NAND2X0 U94 ( .IN1(n371), .IN2(n216), .QN(n364) );
  NAND2X0 U95 ( .IN1(exp_diff_value[0]), .IN2(n3), .QN(n326) );
  NAND2X0 U96 ( .IN1(n607), .IN2(n606), .QN(N389) );
  NAND2X0 U97 ( .IN1(n611), .IN2(n610), .QN(N390) );
  NAND2X0 U98 ( .IN1(n615), .IN2(n614), .QN(N391) );
  NAND2X0 U99 ( .IN1(n619), .IN2(n618), .QN(N392) );
  NAND2X0 U100 ( .IN1(n623), .IN2(n622), .QN(N393) );
  NAND2X0 U101 ( .IN1(n627), .IN2(n626), .QN(N394) );
  NAND2X0 U102 ( .IN1(n631), .IN2(n630), .QN(N395) );
  NAND2X0 U103 ( .IN1(n635), .IN2(n634), .QN(N396) );
  NAND2X0 U104 ( .IN1(n712), .IN2(pre_sig_res_03[9]), .QN(n638) );
  NAND2X0 U105 ( .IN1(n711), .IN2(pre_sig_res_02[9]), .QN(n639) );
  NAND2X0 U106 ( .IN1(n712), .IN2(pre_sig_res_03[10]), .QN(n644) );
  NAND2X0 U107 ( .IN1(n711), .IN2(pre_sig_res_02[10]), .QN(n645) );
  NAND2X0 U108 ( .IN1(n712), .IN2(pre_sig_res_03[11]), .QN(n650) );
  NAND2X0 U109 ( .IN1(n711), .IN2(pre_sig_res_02[11]), .QN(n651) );
  NAND2X0 U110 ( .IN1(n712), .IN2(pre_sig_res_03[12]), .QN(n656) );
  NAND2X0 U111 ( .IN1(n711), .IN2(pre_sig_res_02[12]), .QN(n657) );
  NAND2X0 U112 ( .IN1(n712), .IN2(pre_sig_res_03[13]), .QN(n662) );
  NAND2X0 U113 ( .IN1(n711), .IN2(pre_sig_res_02[13]), .QN(n663) );
  NAND2X0 U114 ( .IN1(n712), .IN2(pre_sig_res_03[14]), .QN(n668) );
  NAND2X0 U115 ( .IN1(n711), .IN2(pre_sig_res_02[14]), .QN(n669) );
  NAND2X0 U116 ( .IN1(n712), .IN2(pre_sig_res_03[15]), .QN(n674) );
  NAND2X0 U117 ( .IN1(n711), .IN2(pre_sig_res_02[15]), .QN(n675) );
  NAND2X0 U118 ( .IN1(n714), .IN2(pre_sig_res_04[16]), .QN(n681) );
  NAND2X0 U119 ( .IN1(n714), .IN2(pre_sig_res_04[17]), .QN(n687) );
  NAND2X0 U120 ( .IN1(n10), .IN2(n11), .QN(N406) );
  NAND2X0 U121 ( .IN1(n714), .IN2(pre_sig_res_04[18]), .QN(n11) );
  NAND2X0 U122 ( .IN1(n8), .IN2(n9), .QN(N407) );
  NAND2X0 U123 ( .IN1(n714), .IN2(pre_sig_res_04[19]), .QN(n9) );
  NAND2X0 U124 ( .IN1(n714), .IN2(pre_sig_res_04[20]), .QN(n697) );
  NAND2X0 U125 ( .IN1(n714), .IN2(pre_sig_res_04[21]), .QN(n705) );
  NAND2X0 U126 ( .IN1(n6), .IN2(n7), .QN(N410) );
  NAND2X0 U127 ( .IN1(n714), .IN2(pre_sig_res_04[22]), .QN(n7) );
  NAND2X0 U128 ( .IN1(n714), .IN2(add_output_exponent_w4[0]), .QN(n567) );
  NAND2X0 U129 ( .IN1(n714), .IN2(add_output_exponent_w4[1]), .QN(n571) );
  NAND2X0 U130 ( .IN1(n714), .IN2(add_output_exponent_w4[2]), .QN(n575) );
  NAND2X0 U131 ( .IN1(n714), .IN2(add_output_exponent_w4[3]), .QN(n581) );
  NAND2X0 U132 ( .IN1(n714), .IN2(add_output_exponent_w4[4]), .QN(n587) );
  NAND2X0 U133 ( .IN1(n714), .IN2(add_output_exponent_w4[5]), .QN(n593) );
  NAND2X0 U134 ( .IN1(n714), .IN2(add_output_exponent_w4[6]), .QN(n599) );
  NAND2X0 U135 ( .IN1(n12), .IN2(n13), .QN(N387) );
  NAND2X0 U136 ( .IN1(n714), .IN2(add_output_exponent_w4[7]), .QN(n13) );
  NAND2X0 U137 ( .IN1(n521), .IN2(n520), .QN(N348) );
  NAND2X0 U138 ( .IN1(n538), .IN2(n796), .QN(n539) );
  NAND2X0 U139 ( .IN1(n538), .IN2(n816), .QN(n529) );
  NAND2X0 U140 ( .IN1(n538), .IN2(n818), .QN(n525) );
  NAND2X0 U141 ( .IN1(n523), .IN2(n522), .QN(N352) );
  NAND2X0 U142 ( .IN1(pre_sig_res_03[22]), .IN2(n820), .QN(n725) );
  NAND2X0 U143 ( .IN1(n809), .IN2(n724), .QN(n726) );
  NAND2X0 U144 ( .IN1(pre_sig_res_03[21]), .IN2(n820), .QN(n733) );
  NAND2X0 U145 ( .IN1(n809), .IN2(n732), .QN(n734) );
  NAND2X0 U146 ( .IN1(pre_sig_res_03[20]), .IN2(n820), .QN(n741) );
  NAND2X0 U147 ( .IN1(n809), .IN2(n740), .QN(n742) );
  NAND2X0 U148 ( .IN1(pre_sig_res_03[19]), .IN2(n820), .QN(n749) );
  NAND2X0 U149 ( .IN1(n809), .IN2(n748), .QN(n750) );
  NAND2X0 U150 ( .IN1(pre_sig_res_03[18]), .IN2(n820), .QN(n757) );
  NAND2X0 U151 ( .IN1(n809), .IN2(n756), .QN(n758) );
  NAND2X0 U152 ( .IN1(pre_sig_res_03[17]), .IN2(n820), .QN(n765) );
  NAND2X0 U153 ( .IN1(n809), .IN2(n764), .QN(n766) );
  NAND2X0 U154 ( .IN1(pre_sig_res_03[16]), .IN2(n820), .QN(n772) );
  NAND2X0 U155 ( .IN1(n809), .IN2(n789), .QN(n773) );
  NAND2X0 U156 ( .IN1(pre_sig_res_03[15]), .IN2(n820), .QN(n781) );
  NAND2X0 U157 ( .IN1(n809), .IN2(n797), .QN(n782) );
  NAND2X0 U158 ( .IN1(n716), .IN2(n723), .QN(n507) );
  NAND2X0 U159 ( .IN1(pre_sig_res_03[14]), .IN2(n848), .QN(n791) );
  NAND2X0 U160 ( .IN1(n819), .IN2(n789), .QN(n790) );
  NAND2X0 U161 ( .IN1(n809), .IN2(n788), .QN(n792) );
  NAND2X0 U162 ( .IN1(pre_sig_res_03[13]), .IN2(n820), .QN(n799) );
  NAND2X0 U163 ( .IN1(n819), .IN2(n797), .QN(n798) );
  NAND2X0 U164 ( .IN1(n809), .IN2(n796), .QN(n800) );
  NAND2X0 U165 ( .IN1(n804), .IN2(n803), .QN(n837) );
  NAND2X0 U166 ( .IN1(pre_sig_res_03[12]), .IN2(n820), .QN(n812) );
  NAND2X0 U167 ( .IN1(n809), .IN2(n816), .QN(n814) );
  NAND2X0 U168 ( .IN1(n414), .IN2(n816), .QN(n415) );
  NAND2X0 U169 ( .IN1(n419), .IN2(n797), .QN(n410) );
  NAND2X0 U170 ( .IN1(n420), .IN2(n796), .QN(n407) );
  NAND2X0 U171 ( .IN1(n406), .IN2(n405), .QN(N263) );
  NAND2X0 U172 ( .IN1(n323), .IN2(n312), .QN(n227) );
  NAND2X0 U173 ( .IN1(n270), .IN2(n244), .QN(n245) );
  NAND2X0 U174 ( .IN1(n313), .IN2(n312), .QN(n314) );
  NAND2X0 U175 ( .IN1(n345), .IN2(n344), .QN(N168) );
  NAND2X0 U176 ( .IN1(n349), .IN2(n348), .QN(N169) );
  NAND2X0 U177 ( .IN1(n361), .IN2(n360), .QN(N172) );
  NAND2X0 U178 ( .IN1(n369), .IN2(n368), .QN(N173) );
  NAND2X0 U179 ( .IN1(n374), .IN2(n373), .QN(N175) );
  INVX0 U180 ( .INP(n393), .ZN(n392) );
  INVX0 U181 ( .INP(n558), .ZN(n825) );
  INVX0 U182 ( .INP(n419), .ZN(n491) );
  NOR2X0 U183 ( .IN1(n821), .IN2(n848), .QN(n822) );
  NOR2X0 U184 ( .IN1(n723), .IN2(n820), .QN(n809) );
  INVX0 U185 ( .INP(n817), .ZN(n807) );
  INVX0 U186 ( .INP(n796), .ZN(n808) );
  INVX0 U187 ( .INP(n797), .ZN(n786) );
  INVX0 U188 ( .INP(n764), .ZN(n777) );
  NOR2X0 U189 ( .IN1(n561), .IN2(n564), .QN(n711) );
  NOR2X0 U190 ( .IN1(n562), .IN2(n564), .QN(n712) );
  INVX0 U191 ( .INP(n740), .ZN(n753) );
  INVX0 U192 ( .INP(n456), .ZN(n560) );
  INVX0 U193 ( .INP(n559), .ZN(n514) );
  INVX0 U194 ( .INP(n748), .ZN(n761) );
  NOR2X0 U195 ( .IN1(n565), .IN2(n564), .QN(n709) );
  NAND4X0 U196 ( .IN1(n554), .IN2(n553), .IN3(n552), .IN4(n551), .QN(n702) );
  INVX0 U197 ( .INP(n710), .ZN(n701) );
  INVX0 U198 ( .INP(n310), .ZN(n203) );
  INVX0 U199 ( .INP(n207), .ZN(n372) );
  NOR2X0 U200 ( .IN1(n74), .IN2(n73), .QN(n821) );
  INVX0 U201 ( .INP(n313), .ZN(n362) );
  INVX0 U202 ( .INP(n72), .ZN(n708) );
  INVX0 U203 ( .INP(n398), .ZN(n494) );
  NOR2X0 U204 ( .IN1(add_sub_result_24_), .IN2(n395), .QN(n565) );
  MUX21X1 U205 ( .IN1(add_result[24]), .IN2(sub_result[24]), .S(n20), .Q(
        add_sub_result_24_) );
  INVX0 U206 ( .INP(n396), .ZN(n484) );
  INVX0 U207 ( .INP(n21), .ZN(n20) );
  INVX0 U208 ( .INP(n503), .ZN(n21) );
  INVX0 U209 ( .INP(n732), .ZN(n745) );
  INVX0 U210 ( .INP(n756), .ZN(n769) );
  INVX0 U211 ( .INP(n789), .ZN(n776) );
  INVX0 U212 ( .INP(n788), .ZN(n806) );
  INVX0 U213 ( .INP(n816), .ZN(n802) );
  INVX0 U214 ( .INP(n818), .ZN(n810) );
  MUX21X1 U215 ( .IN1(input_factor_01[31]), .IN2(n375), .S(input_factor_02[31]), .Q(n503) );
  NAND2X0 U216 ( .IN1(input_factor_02[29]), .IN2(n596), .QN(n49) );
  INVX0 U217 ( .INP(input_factor_02[29]), .ZN(n597) );
  INVX0 U218 ( .INP(input_factor_01[31]), .ZN(n375) );
  NAND4X0 U219 ( .IN1(n32), .IN2(n31), .IN3(n30), .IN4(n35), .QN(n373) );
  INVX0 U220 ( .INP(n447), .ZN(n718) );
  INVX0 U221 ( .INP(n442), .ZN(n729) );
  INVX0 U222 ( .INP(n724), .ZN(n737) );
  INVX0 U223 ( .INP(n819), .ZN(n805) );
  NOR2X0 U224 ( .IN1(n14), .IN2(n15), .QN(n284) );
  NOR2X0 U225 ( .IN1(n336), .IN2(n334), .QN(n14) );
  NOR2X0 U226 ( .IN1(n715), .IN2(n713), .QN(n6) );
  NOR2X0 U227 ( .IN1(n603), .IN2(n602), .QN(n12) );
  NOR2X0 U228 ( .IN1(n693), .IN2(n692), .QN(n8) );
  NOR2X0 U229 ( .IN1(n691), .IN2(n690), .QN(n10) );
  NAND3X0 U230 ( .IN1(n494), .IN2(n401), .IN3(n465), .QN(n483) );
  OR2X1 U231 ( .IN1(n556), .IN2(n753), .Q(n785) );
  NOR2X0 U232 ( .IN1(n16), .IN2(n17), .QN(n228) );
  NOR2X0 U233 ( .IN1(n364), .IN2(n221), .QN(n16) );
  NOR2X0 U234 ( .IN1(n18), .IN2(n19), .QN(n214) );
  NOR2X0 U235 ( .IN1(n356), .IN2(n184), .QN(n18) );
  INVX0 U236 ( .INP(n184), .ZN(n204) );
  INVX0 U237 ( .INP(n326), .ZN(n202) );
  NOR4X0 U238 ( .IN1(n391), .IN2(n390), .IN3(n389), .IN4(n388), .QN(n710) );
  MUX21X1 U239 ( .IN1(add_result[1]), .IN2(sub_result[1]), .S(n503), .Q(n816)
         );
  INVX0 U240 ( .INP(input_factor_02[12]), .ZN(n655) );
  INVX0 U241 ( .INP(input_factor_02[13]), .ZN(n661) );
  INVX0 U242 ( .INP(input_factor_02[14]), .ZN(n667) );
  INVX0 U243 ( .INP(n702), .ZN(n22) );
  INVX0 U244 ( .INP(input_factor_01[29]), .ZN(n596) );
  INVX0 U245 ( .INP(input_factor_02[23]), .ZN(n383) );
  OA222X1 U246 ( .IN1(input_factor_02[29]), .IN2(n596), .IN3(n597), .IN4(
        input_factor_01[29]), .IN5(input_factor_01[23]), .IN6(n383), .Q(n32)
         );
  INVX0 U247 ( .INP(input_factor_01[25]), .ZN(n23) );
  INVX0 U248 ( .INP(n36), .ZN(n29) );
  NOR2X0 U249 ( .IN1(input_factor_02[25]), .IN2(n23), .QN(n41) );
  INVX0 U250 ( .INP(input_factor_02[28]), .ZN(n591) );
  INVX0 U251 ( .INP(input_factor_02[26]), .ZN(n579) );
  INVX0 U252 ( .INP(input_factor_01[28]), .ZN(n590) );
  INVX0 U253 ( .INP(input_factor_01[26]), .ZN(n578) );
  NAND4X0 U254 ( .IN1(n44), .IN2(n34), .IN3(n48), .IN4(n24), .QN(n28) );
  INVX0 U255 ( .INP(input_factor_01[27]), .ZN(n584) );
  INVX0 U256 ( .INP(input_factor_02[27]), .ZN(n585) );
  INVX0 U257 ( .INP(input_factor_01[24]), .ZN(n543) );
  NOR2X0 U258 ( .IN1(n543), .IN2(input_factor_02[24]), .QN(n39) );
  INVX0 U259 ( .INP(n39), .ZN(n25) );
  NAND4X0 U260 ( .IN1(n26), .IN2(n33), .IN3(n37), .IN4(n25), .QN(n27) );
  NOR4X0 U261 ( .IN1(n29), .IN2(n41), .IN3(n28), .IN4(n27), .QN(n31) );
  INVX0 U262 ( .INP(input_factor_01[30]), .ZN(n30) );
  INVX0 U263 ( .INP(n33), .ZN(n47) );
  INVX0 U264 ( .INP(n34), .ZN(n43) );
  INVX0 U265 ( .INP(n35), .ZN(n38) );
  OA221X1 U266 ( .IN1(n39), .IN2(n38), .IN3(n39), .IN4(n37), .IN5(n36), .Q(n40) );
  OA22X1 U267 ( .IN1(n41), .IN2(n40), .IN3(input_factor_01[26]), .IN4(n579), 
        .Q(n42) );
  OA22X1 U268 ( .IN1(n43), .IN2(n42), .IN3(input_factor_01[27]), .IN4(n585), 
        .Q(n46) );
  INVX0 U269 ( .INP(n44), .ZN(n45) );
  AO221X1 U270 ( .IN1(n48), .IN2(n47), .IN3(n48), .IN4(n46), .IN5(n45), .Q(n50) );
  AO221X1 U271 ( .IN1(n50), .IN2(n49), .IN3(n597), .IN4(input_factor_01[29]), 
        .IN5(input_factor_01[30]), .Q(n73) );
  INVX0 U272 ( .INP(n373), .ZN(n74) );
  INVX0 U273 ( .INP(input_factor_02[20]), .ZN(n695) );
  INVX0 U274 ( .INP(input_factor_02[16]), .ZN(n679) );
  INVX0 U275 ( .INP(input_factor_02[15]), .ZN(n673) );
  INVX0 U276 ( .INP(input_factor_02[11]), .ZN(n649) );
  INVX0 U277 ( .INP(input_factor_02[10]), .ZN(n643) );
  INVX0 U278 ( .INP(input_factor_02[9]), .ZN(n637) );
  INVX0 U279 ( .INP(input_factor_02[8]), .ZN(n633) );
  INVX0 U280 ( .INP(input_factor_02[7]), .ZN(n629) );
  INVX0 U281 ( .INP(input_factor_02[6]), .ZN(n625) );
  INVX0 U282 ( .INP(input_factor_02[5]), .ZN(n621) );
  INVX0 U283 ( .INP(input_factor_02[4]), .ZN(n617) );
  INVX0 U284 ( .INP(input_factor_02[3]), .ZN(n613) );
  INVX0 U285 ( .INP(input_factor_02[2]), .ZN(n609) );
  INVX0 U286 ( .INP(input_factor_01[0]), .ZN(n546) );
  NOR2X0 U287 ( .IN1(input_factor_02[0]), .IN2(n546), .QN(n51) );
  INVX0 U288 ( .INP(input_factor_02[1]), .ZN(n605) );
  AO222X1 U289 ( .IN1(input_factor_01[1]), .IN2(n51), .IN3(input_factor_01[1]), 
        .IN4(n605), .IN5(n51), .IN6(n605), .Q(n52) );
  AO222X1 U290 ( .IN1(input_factor_01[2]), .IN2(n609), .IN3(input_factor_01[2]), .IN4(n52), .IN5(n609), .IN6(n52), .Q(n53) );
  AO222X1 U291 ( .IN1(input_factor_01[3]), .IN2(n613), .IN3(input_factor_01[3]), .IN4(n53), .IN5(n613), .IN6(n53), .Q(n54) );
  AO222X1 U292 ( .IN1(input_factor_01[4]), .IN2(n617), .IN3(input_factor_01[4]), .IN4(n54), .IN5(n617), .IN6(n54), .Q(n55) );
  AO222X1 U293 ( .IN1(input_factor_01[5]), .IN2(n621), .IN3(input_factor_01[5]), .IN4(n55), .IN5(n621), .IN6(n55), .Q(n56) );
  AO222X1 U294 ( .IN1(input_factor_01[6]), .IN2(n625), .IN3(input_factor_01[6]), .IN4(n56), .IN5(n625), .IN6(n56), .Q(n57) );
  AO222X1 U295 ( .IN1(input_factor_01[7]), .IN2(n629), .IN3(input_factor_01[7]), .IN4(n57), .IN5(n629), .IN6(n57), .Q(n58) );
  AO222X1 U296 ( .IN1(input_factor_01[8]), .IN2(n633), .IN3(input_factor_01[8]), .IN4(n58), .IN5(n633), .IN6(n58), .Q(n59) );
  AO222X1 U297 ( .IN1(input_factor_01[9]), .IN2(n637), .IN3(input_factor_01[9]), .IN4(n59), .IN5(n637), .IN6(n59), .Q(n60) );
  AO222X1 U298 ( .IN1(input_factor_01[10]), .IN2(n643), .IN3(
        input_factor_01[10]), .IN4(n60), .IN5(n643), .IN6(n60), .Q(n61) );
  AO222X1 U299 ( .IN1(input_factor_01[11]), .IN2(n649), .IN3(
        input_factor_01[11]), .IN4(n61), .IN5(n649), .IN6(n61), .Q(n62) );
  AO222X1 U300 ( .IN1(input_factor_01[12]), .IN2(n655), .IN3(
        input_factor_01[12]), .IN4(n62), .IN5(n655), .IN6(n62), .Q(n63) );
  AO222X1 U301 ( .IN1(input_factor_01[13]), .IN2(n661), .IN3(
        input_factor_01[13]), .IN4(n63), .IN5(n661), .IN6(n63), .Q(n64) );
  AO222X1 U302 ( .IN1(input_factor_01[14]), .IN2(n667), .IN3(
        input_factor_01[14]), .IN4(n64), .IN5(n667), .IN6(n64), .Q(n65) );
  AO222X1 U303 ( .IN1(input_factor_01[15]), .IN2(n673), .IN3(
        input_factor_01[15]), .IN4(n65), .IN5(n673), .IN6(n65), .Q(n66) );
  AO222X1 U304 ( .IN1(input_factor_01[16]), .IN2(n679), .IN3(
        input_factor_01[16]), .IN4(n66), .IN5(n679), .IN6(n66), .Q(n68) );
  INVX0 U305 ( .INP(input_factor_01[17]), .ZN(n684) );
  INVX0 U306 ( .INP(input_factor_02[17]), .ZN(n685) );
  INVX0 U307 ( .INP(input_factor_01[18]), .ZN(n352) );
  INVX0 U308 ( .INP(input_factor_01[19]), .ZN(n356) );
  AO221X1 U309 ( .IN1(n68), .IN2(n67), .IN3(n685), .IN4(input_factor_01[17]), 
        .IN5(n545), .Q(n69) );
  AO222X1 U310 ( .IN1(input_factor_01[20]), .IN2(n695), .IN3(
        input_factor_01[20]), .IN4(n69), .IN5(n695), .IN6(n69), .Q(n71) );
  INVX0 U311 ( .INP(input_factor_01[21]), .ZN(n700) );
  INVX0 U312 ( .INP(input_factor_02[21]), .ZN(n703) );
  AO221X1 U313 ( .IN1(n71), .IN2(n70), .IN3(n703), .IN4(input_factor_01[21]), 
        .IN5(input_factor_01[22]), .Q(n123) );
  NOR2X0 U314 ( .IN1(n392), .IN2(n352), .QN(N194) );
  NOR2X0 U315 ( .IN1(n392), .IN2(n356), .QN(N195) );
  INVX0 U316 ( .INP(input_factor_01[22]), .ZN(n121) );
  NOR2X0 U317 ( .IN1(n392), .IN2(n121), .QN(N198) );
  AO22X1 U318 ( .IN1(input_factor_01[30]), .IN2(rst_n), .IN3(n848), .IN4(
        larger_exponent[7]), .Q(n826) );
  NOR4X0 U319 ( .IN1(exp_diff_value[4]), .IN2(exp_diff_value[5]), .IN3(
        exp_diff_value[6]), .IN4(exp_diff_value[7]), .QN(n370) );
  NOR2X0 U320 ( .IN1(exp_diff_value[3]), .IN2(n2), .QN(n371) );
  INVX0 U321 ( .INP(n371), .ZN(n213) );
  NOR2X0 U322 ( .IN1(n223), .IN2(n213), .QN(n280) );
  INVX0 U323 ( .INP(n280), .ZN(n357) );
  AO21X1 U324 ( .IN1(n121), .IN2(n1), .IN3(exp_diff_value[1]), .Q(n329) );
  INVX0 U325 ( .INP(n199), .ZN(n216) );
  OAI22X1 U326 ( .IN1(n326), .IN2(n357), .IN3(n329), .IN4(n364), .QN(N174) );
  INVX0 U328 ( .INP(input_factor_02[0]), .ZN(n124) );
  OA22X1 U329 ( .IN1(n605), .IN2(n326), .IN3(n124), .IN4(n207), .Q(n76) );
  OA22X1 U330 ( .IN1(n609), .IN2(n310), .IN3(n613), .IN4(n184), .Q(n75) );
  OA22X1 U331 ( .IN1(n633), .IN2(n207), .IN3(n637), .IN4(n326), .Q(n79) );
  OA22X1 U332 ( .IN1(n643), .IN2(n310), .IN3(n649), .IN4(n184), .Q(n77) );
  OA22X1 U333 ( .IN1(n655), .IN2(n207), .IN3(n661), .IN4(n326), .Q(n81) );
  OA22X1 U334 ( .IN1(n673), .IN2(n184), .IN3(n667), .IN4(n310), .Q(n80) );
  MUX21X1 U335 ( .IN1(n218), .IN2(n226), .S(n2), .Q(n285) );
  OA22X1 U336 ( .IN1(n617), .IN2(n207), .IN3(n621), .IN4(n326), .Q(n83) );
  OA22X1 U337 ( .IN1(n625), .IN2(n310), .IN3(n629), .IN4(n184), .Q(n82) );
  NOR2X0 U338 ( .IN1(exp_diff_value[3]), .IN2(n5), .QN(n188) );
  AOI222X1 U339 ( .IN1(n84), .IN2(n371), .IN3(n285), .IN4(exp_diff_value[3]), 
        .IN5(n219), .IN6(n188), .QN(n117) );
  AO22X1 U340 ( .IN1(input_factor_01[9]), .IN2(n202), .IN3(input_factor_01[8]), 
        .IN4(n372), .Q(n86) );
  AO22X1 U341 ( .IN1(input_factor_01[11]), .IN2(n204), .IN3(
        input_factor_01[10]), .IN4(n203), .Q(n85) );
  NOR2X0 U342 ( .IN1(n86), .IN2(n85), .QN(n217) );
  AO22X1 U343 ( .IN1(input_factor_01[13]), .IN2(n202), .IN3(
        input_factor_01[12]), .IN4(n372), .Q(n88) );
  AO22X1 U344 ( .IN1(input_factor_01[15]), .IN2(n204), .IN3(
        input_factor_01[14]), .IN4(n203), .Q(n87) );
  NOR2X0 U345 ( .IN1(n88), .IN2(n87), .QN(n215) );
  MUX21X1 U346 ( .IN1(n217), .IN2(n215), .S(n2), .Q(n287) );
  INVX0 U347 ( .INP(n188), .ZN(n198) );
  AO22X1 U348 ( .IN1(input_factor_01[5]), .IN2(n202), .IN3(input_factor_01[4]), 
        .IN4(n372), .Q(n90) );
  AO22X1 U349 ( .IN1(input_factor_01[7]), .IN2(n204), .IN3(input_factor_01[6]), 
        .IN4(n203), .Q(n89) );
  NOR2X0 U350 ( .IN1(n90), .IN2(n89), .QN(n221) );
  AO22X1 U351 ( .IN1(input_factor_01[0]), .IN2(n372), .IN3(input_factor_01[1]), 
        .IN4(n202), .Q(n92) );
  AO22X1 U352 ( .IN1(input_factor_01[3]), .IN2(n204), .IN3(input_factor_01[2]), 
        .IN4(n203), .Q(n91) );
  NOR2X0 U353 ( .IN1(n92), .IN2(n91), .QN(n93) );
  OA222X1 U354 ( .IN1(n4), .IN2(n287), .IN3(n198), .IN4(n221), .IN5(n213), 
        .IN6(n93), .Q(n116) );
  OA22X1 U355 ( .IN1(n117), .IN2(n223), .IN3(n116), .IN4(n199), .Q(n127) );
  AO221X1 U356 ( .IN1(exp_diff_value[0]), .IN2(n685), .IN3(n1), .IN4(n679), 
        .IN5(exp_diff_value[1]), .Q(n224) );
  OA22X1 U357 ( .IN1(input_factor_02[21]), .IN2(n326), .IN3(
        input_factor_02[20]), .IN4(exp_diff_value[0]), .Q(n311) );
  MUX21X1 U358 ( .IN1(n224), .IN2(n358), .S(n2), .Q(n343) );
  NOR3X0 U359 ( .IN1(exp_diff_value[5]), .IN2(exp_diff_value[6]), .IN3(
        exp_diff_value[7]), .QN(n118) );
  NOR2X0 U360 ( .IN1(exp_diff_value[3]), .IN2(n212), .QN(n122) );
  OA22X1 U361 ( .IN1(n352), .IN2(n310), .IN3(n684), .IN4(n326), .Q(n120) );
  INVX0 U362 ( .INP(input_factor_01[20]), .ZN(n694) );
  AO222X1 U363 ( .IN1(n203), .IN2(n121), .IN3(n202), .IN4(n700), .IN5(n372), 
        .IN6(n694), .Q(n359) );
  MUX21X1 U364 ( .IN1(n214), .IN2(n359), .S(n2), .Q(n342) );
  OA22X1 U365 ( .IN1(n343), .IN2(n235), .IN3(n342), .IN4(n208), .Q(n126) );
  OR2X1 U366 ( .IN1(n373), .IN2(n123), .Q(n366) );
  OA22X1 U367 ( .IN1(n124), .IN2(n367), .IN3(n546), .IN4(n366), .Q(n125) );
  NAND3X0 U368 ( .IN1(n127), .IN2(n126), .IN3(n125), .QN(N152) );
  OA22X1 U369 ( .IN1(n621), .IN2(n207), .IN3(n625), .IN4(n326), .Q(n129) );
  OA22X1 U370 ( .IN1(n633), .IN2(n184), .IN3(n629), .IN4(n310), .Q(n128) );
  OA22X1 U371 ( .IN1(n637), .IN2(n207), .IN3(n643), .IN4(n326), .Q(n131) );
  OA22X1 U372 ( .IN1(n655), .IN2(n184), .IN3(n649), .IN4(n310), .Q(n130) );
  OA22X1 U373 ( .IN1(n661), .IN2(n207), .IN3(n667), .IN4(n326), .Q(n133) );
  OA22X1 U374 ( .IN1(n673), .IN2(n310), .IN3(n679), .IN4(n184), .Q(n132) );
  MUX21X1 U375 ( .IN1(n244), .IN2(n236), .S(n2), .Q(n291) );
  OA22X1 U376 ( .IN1(n605), .IN2(n207), .IN3(n609), .IN4(n326), .Q(n135) );
  OA22X1 U377 ( .IN1(n613), .IN2(n310), .IN3(n617), .IN4(n184), .Q(n134) );
  AOI222X1 U378 ( .IN1(n240), .IN2(n188), .IN3(exp_diff_value[3]), .IN4(n291), 
        .IN5(n136), .IN6(n371), .QN(n148) );
  AO22X1 U379 ( .IN1(input_factor_01[10]), .IN2(n202), .IN3(input_factor_01[9]), .IN4(n372), .Q(n139) );
  AO22X1 U380 ( .IN1(input_factor_01[12]), .IN2(n204), .IN3(
        input_factor_01[11]), .IN4(n203), .Q(n137) );
  NOR2X0 U381 ( .IN1(n139), .IN2(n137), .QN(n239) );
  AO22X1 U382 ( .IN1(input_factor_01[14]), .IN2(n202), .IN3(
        input_factor_01[13]), .IN4(n372), .Q(n141) );
  AO22X1 U383 ( .IN1(input_factor_01[16]), .IN2(n204), .IN3(
        input_factor_01[15]), .IN4(n203), .Q(n140) );
  NOR2X0 U384 ( .IN1(n141), .IN2(n140), .QN(n232) );
  MUX21X1 U385 ( .IN1(n239), .IN2(n232), .S(n2), .Q(n293) );
  AO22X1 U386 ( .IN1(input_factor_01[6]), .IN2(n202), .IN3(input_factor_01[5]), 
        .IN4(n372), .Q(n143) );
  AO22X1 U387 ( .IN1(input_factor_01[8]), .IN2(n204), .IN3(input_factor_01[7]), 
        .IN4(n203), .Q(n142) );
  NOR2X0 U388 ( .IN1(n143), .IN2(n142), .QN(n233) );
  AO22X1 U389 ( .IN1(input_factor_01[2]), .IN2(n202), .IN3(input_factor_01[1]), 
        .IN4(n372), .Q(n145) );
  AO22X1 U390 ( .IN1(input_factor_01[4]), .IN2(n204), .IN3(input_factor_01[3]), 
        .IN4(n203), .Q(n144) );
  NOR2X0 U391 ( .IN1(n145), .IN2(n144), .QN(n146) );
  OA222X1 U392 ( .IN1(n4), .IN2(n293), .IN3(n198), .IN4(n233), .IN5(n213), 
        .IN6(n146), .Q(n147) );
  OA22X1 U393 ( .IN1(n148), .IN2(n223), .IN3(n147), .IN4(n199), .Q(n154) );
  AO22X1 U394 ( .IN1(input_factor_01[18]), .IN2(n202), .IN3(
        input_factor_01[17]), .IN4(n372), .Q(n150) );
  AO22X1 U395 ( .IN1(input_factor_01[20]), .IN2(n204), .IN3(
        input_factor_01[19]), .IN4(n203), .Q(n149) );
  NOR2X0 U396 ( .IN1(n150), .IN2(n149), .QN(n231) );
  AO22X1 U397 ( .IN1(input_factor_01[22]), .IN2(n202), .IN3(
        input_factor_01[21]), .IN4(n1), .Q(n151) );
  NOR2X0 U398 ( .IN1(n203), .IN2(n151), .QN(n365) );
  MUX21X1 U399 ( .IN1(n231), .IN2(n365), .S(n2), .Q(n347) );
  OA22X1 U400 ( .IN1(n685), .IN2(n207), .IN3(n695), .IN4(n184), .Q(n237) );
  AO21X1 U401 ( .IN1(n703), .IN2(n3), .IN3(exp_diff_value[0]), .Q(n234) );
  MUX21X1 U402 ( .IN1(n237), .IN2(n234), .S(n2), .Q(n346) );
  OA22X1 U403 ( .IN1(n208), .IN2(n347), .IN3(n235), .IN4(n346), .Q(n153) );
  INVX0 U404 ( .INP(input_factor_01[1]), .ZN(n604) );
  OA22X1 U405 ( .IN1(n605), .IN2(n367), .IN3(n604), .IN4(n366), .Q(n152) );
  NAND3X0 U406 ( .IN1(n154), .IN2(n153), .IN3(n152), .QN(N153) );
  OA22X1 U407 ( .IN1(n625), .IN2(n207), .IN3(n629), .IN4(n326), .Q(n156) );
  OA22X1 U408 ( .IN1(n633), .IN2(n310), .IN3(n637), .IN4(n184), .Q(n155) );
  OA22X1 U409 ( .IN1(n643), .IN2(n207), .IN3(n649), .IN4(n326), .Q(n158) );
  OA22X1 U410 ( .IN1(n655), .IN2(n310), .IN3(n661), .IN4(n184), .Q(n157) );
  OA22X1 U411 ( .IN1(n673), .IN2(n326), .IN3(n667), .IN4(n207), .Q(n160) );
  OA22X1 U412 ( .IN1(n679), .IN2(n310), .IN3(n685), .IN4(n184), .Q(n159) );
  MUX21X1 U413 ( .IN1(n249), .IN2(n257), .S(n2), .Q(n297) );
  OA22X1 U414 ( .IN1(n609), .IN2(n207), .IN3(n613), .IN4(n326), .Q(n162) );
  OA22X1 U415 ( .IN1(n617), .IN2(n310), .IN3(n621), .IN4(n184), .Q(n161) );
  AOI222X1 U416 ( .IN1(n250), .IN2(n188), .IN3(exp_diff_value[3]), .IN4(n297), 
        .IN5(n163), .IN6(n371), .QN(n174) );
  AO22X1 U417 ( .IN1(input_factor_01[11]), .IN2(n202), .IN3(
        input_factor_01[10]), .IN4(n372), .Q(n165) );
  AO22X1 U418 ( .IN1(input_factor_01[13]), .IN2(n204), .IN3(
        input_factor_01[12]), .IN4(n203), .Q(n164) );
  NOR2X0 U419 ( .IN1(n165), .IN2(n164), .QN(n261) );
  AO22X1 U420 ( .IN1(input_factor_01[15]), .IN2(n202), .IN3(
        input_factor_01[14]), .IN4(n372), .Q(n167) );
  AO22X1 U421 ( .IN1(input_factor_01[17]), .IN2(n204), .IN3(
        input_factor_01[16]), .IN4(n203), .Q(n166) );
  NOR2X0 U422 ( .IN1(n167), .IN2(n166), .QN(n256) );
  MUX21X1 U423 ( .IN1(n261), .IN2(n256), .S(n2), .Q(n299) );
  AO22X1 U424 ( .IN1(input_factor_01[7]), .IN2(n202), .IN3(input_factor_01[6]), 
        .IN4(n372), .Q(n169) );
  AO22X1 U425 ( .IN1(input_factor_01[9]), .IN2(n204), .IN3(input_factor_01[8]), 
        .IN4(n203), .Q(n168) );
  NOR2X0 U426 ( .IN1(n169), .IN2(n168), .QN(n252) );
  AO22X1 U427 ( .IN1(input_factor_01[3]), .IN2(n202), .IN3(input_factor_01[2]), 
        .IN4(n372), .Q(n171) );
  AO22X1 U428 ( .IN1(input_factor_01[5]), .IN2(n204), .IN3(input_factor_01[4]), 
        .IN4(n203), .Q(n170) );
  NOR2X0 U429 ( .IN1(n171), .IN2(n170), .QN(n172) );
  OA222X1 U430 ( .IN1(n4), .IN2(n299), .IN3(n198), .IN4(n252), .IN5(n213), 
        .IN6(n172), .Q(n173) );
  OA22X1 U431 ( .IN1(n174), .IN2(n223), .IN3(n173), .IN4(n199), .Q(n179) );
  AO22X1 U432 ( .IN1(input_factor_01[18]), .IN2(n372), .IN3(
        input_factor_01[19]), .IN4(n202), .Q(n176) );
  AO22X1 U433 ( .IN1(input_factor_01[21]), .IN2(n204), .IN3(
        input_factor_01[20]), .IN4(n203), .Q(n175) );
  NOR2X0 U434 ( .IN1(n176), .IN2(n175), .QN(n255) );
  MUX21X1 U435 ( .IN1(n255), .IN2(n329), .S(n2), .Q(n350) );
  OA22X1 U436 ( .IN1(n695), .IN2(n310), .IN3(n703), .IN4(n184), .Q(n258) );
  MUX21X1 U437 ( .IN1(n258), .IN2(n326), .S(n2), .Q(n351) );
  OA22X1 U438 ( .IN1(n350), .IN2(n208), .IN3(n351), .IN4(n235), .Q(n178) );
  INVX0 U439 ( .INP(input_factor_01[2]), .ZN(n608) );
  OA22X1 U440 ( .IN1(n609), .IN2(n367), .IN3(n608), .IN4(n366), .Q(n177) );
  NAND3X0 U441 ( .IN1(n179), .IN2(n178), .IN3(n177), .QN(N154) );
  OA22X1 U442 ( .IN1(n633), .IN2(n326), .IN3(n629), .IN4(n207), .Q(n181) );
  OA22X1 U443 ( .IN1(n637), .IN2(n310), .IN3(n643), .IN4(n184), .Q(n180) );
  OA22X1 U444 ( .IN1(n655), .IN2(n326), .IN3(n649), .IN4(n207), .Q(n183) );
  OA22X1 U445 ( .IN1(n661), .IN2(n310), .IN3(n667), .IN4(n184), .Q(n182) );
  AO222X1 U446 ( .IN1(input_factor_02[15]), .IN2(n372), .IN3(
        input_factor_02[17]), .IN4(n203), .IN5(input_factor_02[16]), .IN6(n202), .Q(n278) );
  MUX21X1 U447 ( .IN1(n269), .IN2(n278), .S(n2), .Q(n303) );
  OA22X1 U448 ( .IN1(n613), .IN2(n207), .IN3(n617), .IN4(n326), .Q(n186) );
  OA22X1 U449 ( .IN1(n621), .IN2(n310), .IN3(n625), .IN4(n184), .Q(n185) );
  AOI222X1 U450 ( .IN1(n279), .IN2(n188), .IN3(exp_diff_value[3]), .IN4(n303), 
        .IN5(n187), .IN6(n371), .QN(n201) );
  AO22X1 U451 ( .IN1(input_factor_01[12]), .IN2(n202), .IN3(
        input_factor_01[11]), .IN4(n372), .Q(n190) );
  AO22X1 U452 ( .IN1(input_factor_01[14]), .IN2(n204), .IN3(
        input_factor_01[13]), .IN4(n203), .Q(n189) );
  NOR2X0 U453 ( .IN1(n190), .IN2(n189), .QN(n274) );
  AO22X1 U454 ( .IN1(input_factor_01[16]), .IN2(n202), .IN3(
        input_factor_01[15]), .IN4(n372), .Q(n192) );
  AO22X1 U455 ( .IN1(input_factor_01[18]), .IN2(n204), .IN3(
        input_factor_01[17]), .IN4(n203), .Q(n191) );
  NOR2X0 U456 ( .IN1(n192), .IN2(n191), .QN(n268) );
  MUX21X1 U457 ( .IN1(n274), .IN2(n268), .S(n2), .Q(n305) );
  AO22X1 U458 ( .IN1(input_factor_01[8]), .IN2(n202), .IN3(input_factor_01[7]), 
        .IN4(n372), .Q(n194) );
  AO22X1 U459 ( .IN1(input_factor_01[10]), .IN2(n204), .IN3(input_factor_01[9]), .IN4(n203), .Q(n193) );
  NOR2X0 U460 ( .IN1(n194), .IN2(n193), .QN(n275) );
  AO22X1 U461 ( .IN1(input_factor_01[4]), .IN2(n202), .IN3(input_factor_01[3]), 
        .IN4(n372), .Q(n196) );
  AO22X1 U462 ( .IN1(input_factor_01[6]), .IN2(n204), .IN3(input_factor_01[5]), 
        .IN4(n203), .Q(n195) );
  NOR2X0 U463 ( .IN1(n196), .IN2(n195), .QN(n197) );
  OA222X1 U464 ( .IN1(n4), .IN2(n305), .IN3(n198), .IN4(n275), .IN5(n213), 
        .IN6(n197), .Q(n200) );
  OA22X1 U465 ( .IN1(n201), .IN2(n223), .IN3(n200), .IN4(n199), .Q(n211) );
  AO22X1 U466 ( .IN1(input_factor_01[20]), .IN2(n202), .IN3(
        input_factor_01[19]), .IN4(n372), .Q(n206) );
  AO22X1 U467 ( .IN1(input_factor_01[22]), .IN2(n204), .IN3(
        input_factor_01[21]), .IN4(n203), .Q(n205) );
  NOR2X0 U468 ( .IN1(n206), .IN2(n205), .QN(n267) );
  MUX21X1 U469 ( .IN1(n267), .IN2(n207), .S(n2), .Q(n353) );
  OA22X1 U470 ( .IN1(n695), .IN2(n326), .IN3(n703), .IN4(n310), .Q(n276) );
  MUX21X1 U471 ( .IN1(n276), .IN2(n207), .S(n2), .Q(n355) );
  OA22X1 U472 ( .IN1(n353), .IN2(n208), .IN3(n355), .IN4(n235), .Q(n210) );
  INVX0 U473 ( .INP(input_factor_01[3]), .ZN(n612) );
  OA22X1 U474 ( .IN1(n613), .IN2(n367), .IN3(n612), .IN4(n366), .Q(n209) );
  NAND3X0 U475 ( .IN1(n211), .IN2(n210), .IN3(n209), .QN(N155) );
  NOR2X0 U476 ( .IN1(n213), .IN2(n212), .QN(n266) );
  OA22X1 U477 ( .IN1(n359), .IN2(n253), .IN3(n358), .IN4(n254), .Q(n230) );
  OR2X1 U478 ( .IN1(n5), .IN2(n354), .Q(n273) );
  MUX21X1 U479 ( .IN1(n215), .IN2(n214), .S(n2), .Q(n309) );
  OA22X1 U480 ( .IN1(n217), .IN2(n273), .IN3(n309), .IN4(n336), .Q(n229) );
  NOR2X0 U481 ( .IN1(n223), .IN2(exp_diff_value[3]), .QN(n313) );
  NOR2X0 U482 ( .IN1(n5), .IN2(n362), .QN(n270) );
  AOI22X1 U483 ( .IN1(n280), .IN2(n219), .IN3(n270), .IN4(n218), .QN(n222) );
  INVX0 U484 ( .INP(input_factor_01[4]), .ZN(n616) );
  OA22X1 U485 ( .IN1(n617), .IN2(n367), .IN3(n616), .IN4(n366), .Q(n220) );
  NOR2X0 U486 ( .IN1(n223), .IN2(n4), .QN(n323) );
  INVX0 U487 ( .INP(n224), .ZN(n225) );
  MUX21X1 U488 ( .IN1(n226), .IN2(n225), .S(n2), .Q(n312) );
  NAND4X0 U489 ( .IN1(n230), .IN2(n229), .IN3(n228), .IN4(n227), .QN(N156) );
  MUX21X1 U490 ( .IN1(n232), .IN2(n231), .S(n2), .Q(n318) );
  OA22X1 U491 ( .IN1(n233), .IN2(n364), .IN3(n318), .IN4(n336), .Q(n248) );
  OR2X1 U492 ( .IN1(n2), .IN2(n234), .Q(n363) );
  OA22X1 U493 ( .IN1(n365), .IN2(n253), .IN3(n235), .IN4(n363), .Q(n243) );
  INVX0 U494 ( .INP(n236), .ZN(n238) );
  MUX21X1 U495 ( .IN1(n238), .IN2(n237), .S(n2), .Q(n319) );
  INVX0 U496 ( .INP(n323), .ZN(n337) );
  OA22X1 U497 ( .IN1(n239), .IN2(n273), .IN3(n319), .IN4(n337), .Q(n242) );
  AND3X1 U498 ( .IN1(n243), .IN2(n242), .IN3(n241), .Q(n247) );
  INVX0 U499 ( .INP(input_factor_01[5]), .ZN(n620) );
  OA22X1 U500 ( .IN1(n621), .IN2(n367), .IN3(n620), .IN4(n366), .Q(n246) );
  NAND4X0 U501 ( .IN1(n248), .IN2(n247), .IN3(n246), .IN4(n245), .QN(N157) );
  AOI22X1 U502 ( .IN1(n280), .IN2(n250), .IN3(n270), .IN4(n249), .QN(n251) );
  OA21X1 U503 ( .IN1(n252), .IN2(n364), .IN3(n251), .Q(n265) );
  OA22X1 U504 ( .IN1(n326), .IN2(n254), .IN3(n329), .IN4(n253), .Q(n264) );
  MUX21X1 U505 ( .IN1(n256), .IN2(n255), .S(n2), .Q(n327) );
  INVX0 U506 ( .INP(n257), .ZN(n259) );
  MUX21X1 U507 ( .IN1(n259), .IN2(n258), .S(n2), .Q(n324) );
  OA22X1 U508 ( .IN1(n336), .IN2(n327), .IN3(n337), .IN4(n324), .Q(n260) );
  OA21X1 U509 ( .IN1(n261), .IN2(n273), .IN3(n260), .Q(n263) );
  INVX0 U510 ( .INP(input_factor_01[6]), .ZN(n624) );
  OA22X1 U511 ( .IN1(n625), .IN2(n367), .IN3(n624), .IN4(n366), .Q(n262) );
  NAND4X0 U512 ( .IN1(n265), .IN2(n264), .IN3(n263), .IN4(n262), .QN(N158) );
  NAND3X0 U513 ( .IN1(n372), .IN2(n266), .IN3(n373), .QN(n272) );
  MUX21X1 U514 ( .IN1(n268), .IN2(n267), .S(n2), .Q(n334) );
  OA22X1 U515 ( .IN1(n275), .IN2(n364), .IN3(n274), .IN4(n273), .Q(n283) );
  INVX0 U516 ( .INP(n276), .ZN(n277) );
  MUX21X1 U517 ( .IN1(n278), .IN2(n277), .S(n2), .Q(n333) );
  AOI22X1 U518 ( .IN1(n333), .IN2(n323), .IN3(n280), .IN4(n279), .QN(n282) );
  INVX0 U519 ( .INP(input_factor_01[7]), .ZN(n628) );
  OA22X1 U520 ( .IN1(n629), .IN2(n367), .IN3(n628), .IN4(n366), .Q(n281) );
  NAND4X0 U521 ( .IN1(n284), .IN2(n283), .IN3(n282), .IN4(n281), .QN(N159) );
  INVX0 U522 ( .INP(n285), .ZN(n286) );
  OA22X1 U523 ( .IN1(n342), .IN2(n336), .IN3(n286), .IN4(n362), .Q(n290) );
  OA22X1 U524 ( .IN1(n343), .IN2(n337), .IN3(n287), .IN4(n354), .Q(n289) );
  INVX0 U525 ( .INP(input_factor_01[8]), .ZN(n632) );
  OA22X1 U526 ( .IN1(n633), .IN2(n367), .IN3(n632), .IN4(n366), .Q(n288) );
  NAND3X0 U527 ( .IN1(n290), .IN2(n289), .IN3(n288), .QN(N160) );
  INVX0 U528 ( .INP(n291), .ZN(n292) );
  OA22X1 U529 ( .IN1(n292), .IN2(n362), .IN3(n347), .IN4(n336), .Q(n296) );
  OA22X1 U530 ( .IN1(n293), .IN2(n354), .IN3(n346), .IN4(n337), .Q(n295) );
  INVX0 U531 ( .INP(input_factor_01[9]), .ZN(n636) );
  OA22X1 U532 ( .IN1(n637), .IN2(n367), .IN3(n636), .IN4(n366), .Q(n294) );
  NAND3X0 U533 ( .IN1(n296), .IN2(n295), .IN3(n294), .QN(N161) );
  INVX0 U534 ( .INP(n297), .ZN(n298) );
  OA22X1 U535 ( .IN1(n350), .IN2(n336), .IN3(n298), .IN4(n362), .Q(n302) );
  OA22X1 U536 ( .IN1(n351), .IN2(n337), .IN3(n299), .IN4(n354), .Q(n301) );
  INVX0 U537 ( .INP(input_factor_01[10]), .ZN(n642) );
  OA22X1 U538 ( .IN1(n643), .IN2(n367), .IN3(n642), .IN4(n366), .Q(n300) );
  NAND3X0 U539 ( .IN1(n302), .IN2(n301), .IN3(n300), .QN(N162) );
  INVX0 U540 ( .INP(n303), .ZN(n304) );
  OA22X1 U541 ( .IN1(n353), .IN2(n336), .IN3(n304), .IN4(n362), .Q(n308) );
  OA22X1 U542 ( .IN1(n355), .IN2(n337), .IN3(n305), .IN4(n354), .Q(n307) );
  INVX0 U543 ( .INP(input_factor_01[11]), .ZN(n648) );
  OA22X1 U544 ( .IN1(n649), .IN2(n367), .IN3(n648), .IN4(n366), .Q(n306) );
  NAND3X0 U545 ( .IN1(n308), .IN2(n307), .IN3(n306), .QN(N163) );
  OR2X1 U546 ( .IN1(n336), .IN2(n2), .Q(n328) );
  OA22X1 U547 ( .IN1(n359), .IN2(n328), .IN3(n354), .IN4(n309), .Q(n317) );
  INVX0 U548 ( .INP(input_factor_01[12]), .ZN(n654) );
  OA22X1 U549 ( .IN1(n655), .IN2(n367), .IN3(n654), .IN4(n366), .Q(n316) );
  NAND4X0 U550 ( .IN1(n311), .IN2(n323), .IN3(n5), .IN4(n310), .QN(n315) );
  NAND4X0 U551 ( .IN1(n317), .IN2(n316), .IN3(n315), .IN4(n314), .QN(N164) );
  OA22X1 U552 ( .IN1(n362), .IN2(n319), .IN3(n354), .IN4(n318), .Q(n322) );
  OA22X1 U553 ( .IN1(n365), .IN2(n328), .IN3(n363), .IN4(n337), .Q(n321) );
  INVX0 U554 ( .INP(input_factor_01[13]), .ZN(n660) );
  OA22X1 U555 ( .IN1(n661), .IN2(n367), .IN3(n660), .IN4(n366), .Q(n320) );
  NAND3X0 U556 ( .IN1(n322), .IN2(n321), .IN3(n320), .QN(N165) );
  OA22X1 U557 ( .IN1(n326), .IN2(n325), .IN3(n362), .IN4(n324), .Q(n332) );
  OA22X1 U558 ( .IN1(n329), .IN2(n328), .IN3(n354), .IN4(n327), .Q(n331) );
  INVX0 U559 ( .INP(input_factor_01[14]), .ZN(n666) );
  OA22X1 U560 ( .IN1(n667), .IN2(n367), .IN3(n666), .IN4(n366), .Q(n330) );
  NAND3X0 U561 ( .IN1(n332), .IN2(n331), .IN3(n330), .QN(N166) );
  INVX0 U562 ( .INP(n333), .ZN(n335) );
  OA22X1 U563 ( .IN1(n362), .IN2(n335), .IN3(n354), .IN4(n334), .Q(n341) );
  INVX0 U564 ( .INP(input_factor_01[15]), .ZN(n672) );
  OA22X1 U565 ( .IN1(n673), .IN2(n367), .IN3(n672), .IN4(n366), .Q(n340) );
  NAND3X0 U566 ( .IN1(n338), .IN2(n5), .IN3(n372), .QN(n339) );
  NAND3X0 U567 ( .IN1(n341), .IN2(n340), .IN3(n339), .QN(N167) );
  OA22X1 U568 ( .IN1(n343), .IN2(n362), .IN3(n342), .IN4(n354), .Q(n345) );
  INVX0 U569 ( .INP(input_factor_01[16]), .ZN(n678) );
  OA22X1 U570 ( .IN1(n679), .IN2(n367), .IN3(n678), .IN4(n366), .Q(n344) );
  OA22X1 U571 ( .IN1(n347), .IN2(n354), .IN3(n346), .IN4(n362), .Q(n349) );
  OA22X1 U572 ( .IN1(n685), .IN2(n367), .IN3(n684), .IN4(n366), .Q(n348) );
  OAI222X1 U573 ( .IN1(n366), .IN2(n352), .IN3(n362), .IN4(n351), .IN5(n354), 
        .IN6(n350), .QN(N170) );
  OAI222X1 U574 ( .IN1(n366), .IN2(n356), .IN3(n362), .IN4(n355), .IN5(n354), 
        .IN6(n353), .QN(N171) );
  OA22X1 U575 ( .IN1(n359), .IN2(n364), .IN3(n358), .IN4(n357), .Q(n361) );
  OA22X1 U576 ( .IN1(n695), .IN2(n367), .IN3(n694), .IN4(n366), .Q(n360) );
  OA22X1 U577 ( .IN1(n365), .IN2(n364), .IN3(n363), .IN4(n362), .Q(n369) );
  OA22X1 U578 ( .IN1(n703), .IN2(n367), .IN3(n700), .IN4(n366), .Q(n368) );
  NAND3X0 U579 ( .IN1(n372), .IN2(n371), .IN3(n370), .QN(n374) );
  MUX21X1 U580 ( .IN1(input_factor_01[0]), .IN2(input_factor_02[0]), .S(n392), 
        .Q(N176) );
  MUX21X1 U581 ( .IN1(input_factor_01[1]), .IN2(input_factor_02[1]), .S(n392), 
        .Q(N177) );
  MUX21X1 U582 ( .IN1(input_factor_01[2]), .IN2(input_factor_02[2]), .S(n392), 
        .Q(N178) );
  MUX21X1 U583 ( .IN1(input_factor_01[3]), .IN2(input_factor_02[3]), .S(n392), 
        .Q(N179) );
  MUX21X1 U584 ( .IN1(input_factor_01[4]), .IN2(input_factor_02[4]), .S(n392), 
        .Q(N180) );
  MUX21X1 U585 ( .IN1(input_factor_01[5]), .IN2(input_factor_02[5]), .S(n392), 
        .Q(N181) );
  MUX21X1 U586 ( .IN1(input_factor_01[6]), .IN2(input_factor_02[6]), .S(n392), 
        .Q(N182) );
  MUX21X1 U587 ( .IN1(input_factor_01[7]), .IN2(input_factor_02[7]), .S(n392), 
        .Q(N183) );
  MUX21X1 U588 ( .IN1(input_factor_01[8]), .IN2(input_factor_02[8]), .S(n392), 
        .Q(N184) );
  MUX21X1 U589 ( .IN1(input_factor_01[9]), .IN2(input_factor_02[9]), .S(n392), 
        .Q(N185) );
  MUX21X1 U590 ( .IN1(input_factor_01[10]), .IN2(input_factor_02[10]), .S(n392), .Q(N186) );
  MUX21X1 U591 ( .IN1(input_factor_01[11]), .IN2(input_factor_02[11]), .S(n392), .Q(N187) );
  MUX21X1 U592 ( .IN1(input_factor_01[12]), .IN2(input_factor_02[12]), .S(n392), .Q(N188) );
  MUX21X1 U593 ( .IN1(input_factor_01[13]), .IN2(input_factor_02[13]), .S(n392), .Q(N189) );
  MUX21X1 U594 ( .IN1(input_factor_01[14]), .IN2(input_factor_02[14]), .S(n392), .Q(N190) );
  MUX21X1 U595 ( .IN1(input_factor_01[15]), .IN2(input_factor_02[15]), .S(n392), .Q(N191) );
  MUX21X1 U596 ( .IN1(input_factor_01[16]), .IN2(input_factor_02[16]), .S(n392), .Q(N192) );
  MUX21X1 U597 ( .IN1(input_factor_01[17]), .IN2(input_factor_02[17]), .S(n392), .Q(N193) );
  MUX21X1 U598 ( .IN1(input_factor_01[20]), .IN2(input_factor_02[20]), .S(n392), .Q(N196) );
  MUX21X1 U599 ( .IN1(input_factor_01[21]), .IN2(input_factor_02[21]), .S(n392), .Q(N197) );
  MUX21X1 U600 ( .IN1(add_result[0]), .IN2(sub_result[0]), .S(n503), .Q(n818)
         );
  MUX21X1 U601 ( .IN1(add_result[2]), .IN2(sub_result[2]), .S(n503), .Q(n796)
         );
  MUX21X1 U602 ( .IN1(add_result[3]), .IN2(sub_result[3]), .S(n503), .Q(n788)
         );
  MUX21X1 U603 ( .IN1(add_result[4]), .IN2(sub_result[4]), .S(n503), .Q(n797)
         );
  MUX21X1 U604 ( .IN1(add_result[5]), .IN2(sub_result[5]), .S(n503), .Q(n789)
         );
  MUX21X1 U605 ( .IN1(add_result[6]), .IN2(sub_result[6]), .S(n503), .Q(n764)
         );
  MUX21X1 U606 ( .IN1(add_result[7]), .IN2(sub_result[7]), .S(n503), .Q(n756)
         );
  MUX21X1 U607 ( .IN1(add_result[9]), .IN2(sub_result[9]), .S(n503), .Q(n740)
         );
  MUX21X1 U608 ( .IN1(add_result[10]), .IN2(sub_result[10]), .S(n503), .Q(n732) );
  NOR4X0 U609 ( .IN1(n503), .IN2(add_result[14]), .IN3(add_result[15]), .IN4(
        add_result[13]), .QN(n512) );
  NOR4X0 U610 ( .IN1(sub_result[15]), .IN2(sub_result[14]), .IN3(
        sub_result[13]), .IN4(n21), .QN(n510) );
  NOR2X0 U611 ( .IN1(n512), .IN2(n510), .QN(n379) );
  MUX21X1 U612 ( .IN1(add_result[11]), .IN2(sub_result[11]), .S(n503), .Q(n724) );
  MUX21X1 U613 ( .IN1(add_result[16]), .IN2(sub_result[16]), .S(n20), .Q(n396)
         );
  MUX21X1 U614 ( .IN1(add_result[17]), .IN2(sub_result[17]), .S(n20), .Q(n465)
         );
  MUX21X1 U615 ( .IN1(add_result[20]), .IN2(sub_result[20]), .S(n20), .Q(n399)
         );
  INVX0 U616 ( .INP(n399), .ZN(n492) );
  MUX21X1 U617 ( .IN1(add_result[22]), .IN2(sub_result[22]), .S(n20), .Q(n400)
         );
  INVX0 U618 ( .INP(n400), .ZN(n376) );
  MUX21X1 U619 ( .IN1(add_result[23]), .IN2(sub_result[23]), .S(n20), .Q(n395)
         );
  MUX21X1 U620 ( .IN1(add_result[21]), .IN2(sub_result[21]), .S(n20), .Q(n402)
         );
  NOR2X0 U621 ( .IN1(n403), .IN2(n402), .QN(n404) );
  MUX21X1 U622 ( .IN1(add_result[19]), .IN2(sub_result[19]), .S(n20), .Q(n474)
         );
  NOR2X0 U623 ( .IN1(n377), .IN2(n474), .QN(n401) );
  MUX21X1 U624 ( .IN1(add_result[18]), .IN2(sub_result[18]), .S(n20), .Q(n398)
         );
  NOR2X0 U625 ( .IN1(n465), .IN2(n378), .QN(n397) );
  MUX21X1 U626 ( .IN1(add_result[12]), .IN2(sub_result[12]), .S(n20), .Q(n442)
         );
  NOR4X0 U627 ( .IN1(n379), .IN2(n724), .IN3(n559), .IN4(n442), .QN(n719) );
  MUX21X1 U628 ( .IN1(add_result[8]), .IN2(sub_result[8]), .S(n20), .Q(n748)
         );
  NOR3X0 U629 ( .IN1(n740), .IN2(n556), .IN3(n748), .QN(n517) );
  NOR2X0 U630 ( .IN1(n764), .IN2(n380), .QN(n516) );
  NOR2X0 U631 ( .IN1(n797), .IN2(n381), .QN(n524) );
  NOR2X0 U632 ( .IN1(n796), .IN2(n382), .QN(n518) );
  NAND3X0 U633 ( .IN1(n810), .IN2(n802), .IN3(n518), .QN(n557) );
  NAND4X0 U634 ( .IN1(n655), .IN2(n673), .IN3(n661), .IN4(n667), .QN(n391) );
  OR4X1 U635 ( .IN1(input_factor_02[31]), .IN2(input_factor_02[27]), .IN3(
        input_factor_02[24]), .IN4(input_factor_02[25]), .Q(n390) );
  NAND4X0 U636 ( .IN1(n597), .IN2(n383), .IN3(n591), .IN4(n579), .QN(n389) );
  NOR4X0 U637 ( .IN1(input_factor_02[1]), .IN2(input_factor_02[0]), .IN3(
        input_factor_02[2]), .IN4(input_factor_02[3]), .QN(n387) );
  NOR4X0 U638 ( .IN1(input_factor_02[16]), .IN2(input_factor_02[17]), .IN3(
        input_factor_02[20]), .IN4(input_factor_02[21]), .QN(n386) );
  NOR4X0 U639 ( .IN1(input_factor_02[7]), .IN2(input_factor_02[9]), .IN3(
        input_factor_02[10]), .IN4(input_factor_02[11]), .QN(n385) );
  NOR4X0 U640 ( .IN1(input_factor_02[4]), .IN2(input_factor_02[5]), .IN3(
        input_factor_02[8]), .IN4(input_factor_02[6]), .QN(n384) );
  NAND4X0 U641 ( .IN1(n387), .IN2(n386), .IN3(n385), .IN4(n384), .QN(n388) );
  AO222X1 U642 ( .IN1(input_factor_01[31]), .IN2(n710), .IN3(
        input_factor_01[31]), .IN4(n393), .IN5(n392), .IN6(input_factor_02[31]), .Q(n394) );
  AND2X1 U643 ( .IN1(n557), .IN2(n394), .Q(N211) );
  MUX21X1 U644 ( .IN1(n818), .IN2(n816), .S(add_sub_result_24_), .Q(N226) );
  MUX21X1 U645 ( .IN1(n816), .IN2(n796), .S(add_sub_result_24_), .Q(N227) );
  MUX21X1 U646 ( .IN1(n796), .IN2(n788), .S(add_sub_result_24_), .Q(N228) );
  MUX21X1 U647 ( .IN1(n788), .IN2(n797), .S(add_sub_result_24_), .Q(N229) );
  MUX21X1 U648 ( .IN1(n797), .IN2(n789), .S(add_sub_result_24_), .Q(N230) );
  MUX21X1 U649 ( .IN1(n789), .IN2(n764), .S(add_sub_result_24_), .Q(N231) );
  MUX21X1 U650 ( .IN1(n764), .IN2(n756), .S(add_sub_result_24_), .Q(N232) );
  MUX21X1 U651 ( .IN1(n756), .IN2(n748), .S(add_sub_result_24_), .Q(N233) );
  MUX21X1 U652 ( .IN1(n748), .IN2(n740), .S(add_sub_result_24_), .Q(N234) );
  MUX21X1 U653 ( .IN1(n740), .IN2(n732), .S(add_sub_result_24_), .Q(N235) );
  MUX21X1 U654 ( .IN1(n732), .IN2(n724), .S(add_sub_result_24_), .Q(N236) );
  MUX21X1 U655 ( .IN1(n724), .IN2(n442), .S(add_sub_result_24_), .Q(N237) );
  MUX21X1 U656 ( .IN1(add_result[13]), .IN2(sub_result[13]), .S(n20), .Q(n447)
         );
  MUX21X1 U657 ( .IN1(n442), .IN2(n447), .S(add_sub_result_24_), .Q(N238) );
  MUX21X1 U658 ( .IN1(add_result[14]), .IN2(sub_result[14]), .S(n20), .Q(n501)
         );
  MUX21X1 U659 ( .IN1(n447), .IN2(n501), .S(add_sub_result_24_), .Q(N239) );
  MUX21X1 U660 ( .IN1(add_result[15]), .IN2(sub_result[15]), .S(n20), .Q(n456)
         );
  MUX21X1 U661 ( .IN1(n501), .IN2(n456), .S(add_sub_result_24_), .Q(N240) );
  MUX21X1 U662 ( .IN1(n456), .IN2(n396), .S(add_sub_result_24_), .Q(N241) );
  MUX21X1 U663 ( .IN1(n396), .IN2(n465), .S(add_sub_result_24_), .Q(N242) );
  MUX21X1 U664 ( .IN1(n465), .IN2(n398), .S(add_sub_result_24_), .Q(N243) );
  MUX21X1 U665 ( .IN1(n398), .IN2(n474), .S(add_sub_result_24_), .Q(N244) );
  MUX21X1 U666 ( .IN1(n474), .IN2(n399), .S(add_sub_result_24_), .Q(N245) );
  MUX21X1 U667 ( .IN1(n399), .IN2(n402), .S(add_sub_result_24_), .Q(N246) );
  MUX21X1 U668 ( .IN1(n402), .IN2(n400), .S(add_sub_result_24_), .Q(N247) );
  MUX21X1 U669 ( .IN1(n400), .IN2(n395), .S(add_sub_result_24_), .Q(N248) );
  NAND4X0 U670 ( .IN1(n496), .IN2(n485), .IN3(n489), .IN4(n487), .QN(N256) );
  INVX0 U671 ( .INP(n402), .ZN(n488) );
  NOR2X0 U672 ( .IN1(n488), .IN2(n403), .QN(n419) );
  NAND4X0 U673 ( .IN1(n496), .IN2(n483), .IN3(n489), .IN4(n491), .QN(N257) );
  NAND3X0 U674 ( .IN1(n404), .IN2(n492), .IN3(n474), .QN(n493) );
  NAND4X0 U675 ( .IN1(n496), .IN2(n485), .IN3(n493), .IN4(n483), .QN(N258) );
  NOR2X0 U676 ( .IN1(n810), .IN2(n487), .QN(N260) );
  INVX0 U677 ( .INP(n487), .ZN(n421) );
  AO22X1 U678 ( .IN1(n421), .IN2(n816), .IN3(n419), .IN4(n818), .Q(N261) );
  INVX0 U679 ( .INP(n489), .ZN(n420) );
  AO222X1 U680 ( .IN1(n818), .IN2(n420), .IN3(n816), .IN4(n419), .IN5(n796), 
        .IN6(n421), .Q(N262) );
  OA22X1 U681 ( .IN1(n802), .IN2(n489), .IN3(n810), .IN4(n493), .Q(n406) );
  OA22X1 U682 ( .IN1(n808), .IN2(n491), .IN3(n806), .IN4(n487), .Q(n405) );
  OA22X1 U683 ( .IN1(n786), .IN2(n487), .IN3(n806), .IN4(n491), .Q(n409) );
  OA22X1 U684 ( .IN1(n802), .IN2(n493), .IN3(n810), .IN4(n485), .Q(n408) );
  NAND3X0 U685 ( .IN1(n409), .IN2(n408), .IN3(n407), .QN(N264) );
  OA22X1 U686 ( .IN1(n776), .IN2(n487), .IN3(n806), .IN4(n489), .Q(n413) );
  OA22X1 U687 ( .IN1(n808), .IN2(n493), .IN3(n802), .IN4(n485), .Q(n412) );
  INVX0 U688 ( .INP(n483), .ZN(n414) );
  NAND4X0 U689 ( .IN1(n413), .IN2(n412), .IN3(n411), .IN4(n410), .QN(N265) );
  OA22X1 U690 ( .IN1(n786), .IN2(n489), .IN3(n806), .IN4(n493), .Q(n418) );
  OA22X1 U691 ( .IN1(n777), .IN2(n487), .IN3(n776), .IN4(n491), .Q(n417) );
  OA22X1 U692 ( .IN1(n808), .IN2(n485), .IN3(n810), .IN4(n496), .Q(n416) );
  NAND4X0 U693 ( .IN1(n418), .IN2(n417), .IN3(n416), .IN4(n415), .QN(N266) );
  NOR4X0 U694 ( .IN1(n421), .IN2(n420), .IN3(n419), .IN4(N258), .QN(n558) );
  OA22X1 U695 ( .IN1(n808), .IN2(n483), .IN3(n806), .IN4(n485), .Q(n425) );
  OA22X1 U696 ( .IN1(n769), .IN2(n487), .IN3(n776), .IN4(n489), .Q(n424) );
  OA22X1 U697 ( .IN1(n777), .IN2(n491), .IN3(n786), .IN4(n493), .Q(n423) );
  OA22X1 U698 ( .IN1(n802), .IN2(n496), .IN3(n810), .IN4(n825), .Q(n422) );
  NAND4X0 U699 ( .IN1(n425), .IN2(n424), .IN3(n423), .IN4(n422), .QN(N267) );
  OA22X1 U700 ( .IN1(n786), .IN2(n485), .IN3(n806), .IN4(n483), .Q(n429) );
  OA22X1 U701 ( .IN1(n761), .IN2(n487), .IN3(n777), .IN4(n489), .Q(n428) );
  OA22X1 U702 ( .IN1(n769), .IN2(n491), .IN3(n776), .IN4(n493), .Q(n427) );
  OA22X1 U703 ( .IN1(n808), .IN2(n496), .IN3(n802), .IN4(n825), .Q(n426) );
  NAND4X0 U704 ( .IN1(n429), .IN2(n428), .IN3(n427), .IN4(n426), .QN(N268) );
  OA22X1 U705 ( .IN1(n776), .IN2(n485), .IN3(n786), .IN4(n483), .Q(n433) );
  OA22X1 U706 ( .IN1(n753), .IN2(n487), .IN3(n769), .IN4(n489), .Q(n432) );
  OA22X1 U707 ( .IN1(n761), .IN2(n491), .IN3(n777), .IN4(n493), .Q(n431) );
  OA22X1 U708 ( .IN1(n808), .IN2(n825), .IN3(n806), .IN4(n496), .Q(n430) );
  NAND4X0 U709 ( .IN1(n433), .IN2(n432), .IN3(n431), .IN4(n430), .QN(N269) );
  OA22X1 U710 ( .IN1(n777), .IN2(n485), .IN3(n776), .IN4(n483), .Q(n437) );
  OA22X1 U711 ( .IN1(n761), .IN2(n489), .IN3(n745), .IN4(n487), .Q(n436) );
  OA22X1 U712 ( .IN1(n753), .IN2(n491), .IN3(n769), .IN4(n493), .Q(n435) );
  OA22X1 U713 ( .IN1(n786), .IN2(n496), .IN3(n806), .IN4(n825), .Q(n434) );
  NAND4X0 U714 ( .IN1(n437), .IN2(n436), .IN3(n435), .IN4(n434), .QN(N270) );
  OA22X1 U715 ( .IN1(n769), .IN2(n485), .IN3(n777), .IN4(n483), .Q(n441) );
  OA22X1 U716 ( .IN1(n737), .IN2(n487), .IN3(n753), .IN4(n489), .Q(n440) );
  OA22X1 U717 ( .IN1(n761), .IN2(n493), .IN3(n745), .IN4(n491), .Q(n439) );
  OA22X1 U718 ( .IN1(n776), .IN2(n496), .IN3(n786), .IN4(n825), .Q(n438) );
  NAND4X0 U719 ( .IN1(n441), .IN2(n440), .IN3(n439), .IN4(n438), .QN(N271) );
  OA22X1 U720 ( .IN1(n761), .IN2(n485), .IN3(n769), .IN4(n483), .Q(n446) );
  OA22X1 U721 ( .IN1(n729), .IN2(n487), .IN3(n745), .IN4(n489), .Q(n445) );
  OA22X1 U722 ( .IN1(n737), .IN2(n491), .IN3(n753), .IN4(n493), .Q(n444) );
  OA22X1 U723 ( .IN1(n777), .IN2(n496), .IN3(n776), .IN4(n825), .Q(n443) );
  NAND4X0 U724 ( .IN1(n446), .IN2(n445), .IN3(n444), .IN4(n443), .QN(N272) );
  OA22X1 U725 ( .IN1(n761), .IN2(n483), .IN3(n753), .IN4(n485), .Q(n451) );
  OA22X1 U726 ( .IN1(n737), .IN2(n489), .IN3(n718), .IN4(n487), .Q(n450) );
  OA22X1 U727 ( .IN1(n729), .IN2(n491), .IN3(n745), .IN4(n493), .Q(n449) );
  OA22X1 U728 ( .IN1(n769), .IN2(n496), .IN3(n777), .IN4(n825), .Q(n448) );
  NAND4X0 U729 ( .IN1(n451), .IN2(n450), .IN3(n449), .IN4(n448), .QN(N273) );
  OA22X1 U730 ( .IN1(n745), .IN2(n485), .IN3(n753), .IN4(n483), .Q(n455) );
  INVX0 U731 ( .INP(n501), .ZN(n495) );
  OA22X1 U732 ( .IN1(n495), .IN2(n487), .IN3(n729), .IN4(n489), .Q(n454) );
  OA22X1 U733 ( .IN1(n737), .IN2(n493), .IN3(n718), .IN4(n491), .Q(n453) );
  OA22X1 U734 ( .IN1(n761), .IN2(n496), .IN3(n769), .IN4(n825), .Q(n452) );
  NAND4X0 U735 ( .IN1(n455), .IN2(n454), .IN3(n453), .IN4(n452), .QN(N274) );
  OA22X1 U736 ( .IN1(n737), .IN2(n485), .IN3(n745), .IN4(n483), .Q(n460) );
  OA22X1 U737 ( .IN1(n560), .IN2(n487), .IN3(n718), .IN4(n489), .Q(n459) );
  OA22X1 U738 ( .IN1(n495), .IN2(n491), .IN3(n729), .IN4(n493), .Q(n458) );
  OA22X1 U739 ( .IN1(n761), .IN2(n825), .IN3(n753), .IN4(n496), .Q(n457) );
  NAND4X0 U740 ( .IN1(n460), .IN2(n459), .IN3(n458), .IN4(n457), .QN(N275) );
  OA22X1 U741 ( .IN1(n729), .IN2(n485), .IN3(n737), .IN4(n483), .Q(n464) );
  OA22X1 U742 ( .IN1(n495), .IN2(n489), .IN3(n484), .IN4(n487), .Q(n463) );
  OA22X1 U743 ( .IN1(n560), .IN2(n491), .IN3(n718), .IN4(n493), .Q(n462) );
  OA22X1 U744 ( .IN1(n745), .IN2(n496), .IN3(n753), .IN4(n825), .Q(n461) );
  NAND4X0 U745 ( .IN1(n464), .IN2(n463), .IN3(n462), .IN4(n461), .QN(N276) );
  OA22X1 U746 ( .IN1(n729), .IN2(n483), .IN3(n718), .IN4(n485), .Q(n469) );
  INVX0 U747 ( .INP(n465), .ZN(n486) );
  OA22X1 U748 ( .IN1(n560), .IN2(n489), .IN3(n486), .IN4(n487), .Q(n468) );
  OA22X1 U749 ( .IN1(n495), .IN2(n493), .IN3(n484), .IN4(n491), .Q(n467) );
  OA22X1 U750 ( .IN1(n737), .IN2(n496), .IN3(n745), .IN4(n825), .Q(n466) );
  NAND4X0 U751 ( .IN1(n469), .IN2(n468), .IN3(n467), .IN4(n466), .QN(N277) );
  OA22X1 U752 ( .IN1(n495), .IN2(n485), .IN3(n718), .IN4(n483), .Q(n473) );
  OA22X1 U753 ( .IN1(n494), .IN2(n487), .IN3(n484), .IN4(n489), .Q(n472) );
  OA22X1 U754 ( .IN1(n560), .IN2(n493), .IN3(n486), .IN4(n491), .Q(n471) );
  OA22X1 U755 ( .IN1(n729), .IN2(n496), .IN3(n737), .IN4(n825), .Q(n470) );
  NAND4X0 U756 ( .IN1(n473), .IN2(n472), .IN3(n471), .IN4(n470), .QN(N278) );
  OA22X1 U757 ( .IN1(n560), .IN2(n485), .IN3(n495), .IN4(n483), .Q(n478) );
  INVX0 U758 ( .INP(n474), .ZN(n490) );
  OA22X1 U759 ( .IN1(n486), .IN2(n489), .IN3(n490), .IN4(n487), .Q(n477) );
  OA22X1 U760 ( .IN1(n494), .IN2(n491), .IN3(n484), .IN4(n493), .Q(n476) );
  OA22X1 U761 ( .IN1(n729), .IN2(n825), .IN3(n718), .IN4(n496), .Q(n475) );
  NAND4X0 U762 ( .IN1(n478), .IN2(n477), .IN3(n476), .IN4(n475), .QN(N279) );
  OA22X1 U763 ( .IN1(n560), .IN2(n483), .IN3(n484), .IN4(n485), .Q(n482) );
  OA22X1 U764 ( .IN1(n494), .IN2(n489), .IN3(n492), .IN4(n487), .Q(n481) );
  OA22X1 U765 ( .IN1(n486), .IN2(n493), .IN3(n490), .IN4(n491), .Q(n480) );
  OA22X1 U766 ( .IN1(n495), .IN2(n496), .IN3(n718), .IN4(n825), .Q(n479) );
  NAND4X0 U767 ( .IN1(n482), .IN2(n481), .IN3(n480), .IN4(n479), .QN(N280) );
  OA22X1 U768 ( .IN1(n486), .IN2(n485), .IN3(n484), .IN4(n483), .Q(n500) );
  OA22X1 U769 ( .IN1(n490), .IN2(n489), .IN3(n488), .IN4(n487), .Q(n499) );
  OA22X1 U770 ( .IN1(n494), .IN2(n493), .IN3(n492), .IN4(n491), .Q(n498) );
  OA22X1 U771 ( .IN1(n560), .IN2(n496), .IN3(n495), .IN4(n825), .Q(n497) );
  NAND4X0 U772 ( .IN1(n500), .IN2(n499), .IN3(n498), .IN4(n497), .QN(N281) );
  NAND3X0 U773 ( .IN1(n501), .IN2(n514), .IN3(n560), .QN(n717) );
  AO22X1 U774 ( .IN1(n512), .IN2(add_result[12]), .IN3(n510), .IN4(
        sub_result[12]), .Q(n502) );
  INVX0 U775 ( .INP(n717), .ZN(n508) );
  NOR3X0 U776 ( .IN1(n503), .IN2(add_result[14]), .IN3(add_result[15]), .QN(
        n505) );
  NOR3X0 U777 ( .IN1(sub_result[14]), .IN2(sub_result[15]), .IN3(n21), .QN(
        n504) );
  AO22X1 U778 ( .IN1(n505), .IN2(add_result[13]), .IN3(n504), .IN4(
        sub_result[13]), .Q(n506) );
  NOR2X0 U779 ( .IN1(n508), .IN2(n507), .QN(N308) );
  INVX0 U780 ( .INP(add_result[12]), .ZN(n511) );
  INVX0 U781 ( .INP(sub_result[12]), .ZN(n509) );
  AO22X1 U782 ( .IN1(n512), .IN2(n511), .IN3(n510), .IN4(n509), .Q(n513) );
  NAND3X0 U783 ( .IN1(n514), .IN2(n724), .IN3(n513), .QN(n811) );
  NAND4X0 U784 ( .IN1(N308), .IN2(n811), .IN3(n794), .IN4(n785), .QN(n778) );
  NAND4X0 U785 ( .IN1(n794), .IN2(n717), .IN3(n723), .IN4(n778), .QN(N306) );
  NAND4X0 U786 ( .IN1(n785), .IN2(n716), .IN3(n723), .IN4(n778), .QN(N307) );
  AO22X1 U787 ( .IN1(n708), .IN2(exponent_factor_12[0]), .IN3(n821), .IN4(
        exponent_factor_21[0]), .Q(N34) );
  NAND3X0 U788 ( .IN1(n806), .IN2(n524), .IN3(n796), .QN(n537) );
  NAND3X0 U789 ( .IN1(n776), .IN2(n516), .IN3(n797), .QN(n532) );
  NAND3X0 U790 ( .IN1(n769), .IN2(n517), .IN3(n764), .QN(n533) );
  NAND3X0 U791 ( .IN1(n808), .IN2(n802), .IN3(n806), .QN(n515) );
  AND2X1 U792 ( .IN1(n532), .IN2(n534), .Q(n519) );
  NAND4X0 U793 ( .IN1(n521), .IN2(n519), .IN3(n533), .IN4(n535), .QN(n520) );
  NAND4X0 U794 ( .IN1(n537), .IN2(n532), .IN3(n533), .IN4(n520), .QN(N346) );
  NAND3X0 U795 ( .IN1(n519), .IN2(n536), .IN3(n520), .QN(N347) );
  NOR2X0 U796 ( .IN1(n810), .IN2(n535), .QN(N349) );
  AO22X1 U797 ( .IN1(n708), .IN2(exponent_factor_12[1]), .IN3(n821), .IN4(
        exponent_factor_21[1]), .Q(N35) );
  OAI22X1 U798 ( .IN1(n802), .IN2(n535), .IN3(n810), .IN4(n533), .QN(N350) );
  OAI222X1 U799 ( .IN1(n534), .IN2(n810), .IN3(n533), .IN4(n802), .IN5(n535), 
        .IN6(n808), .QN(N351) );
  OA22X1 U800 ( .IN1(n808), .IN2(n533), .IN3(n806), .IN4(n535), .Q(n523) );
  OA22X1 U801 ( .IN1(n802), .IN2(n534), .IN3(n810), .IN4(n532), .Q(n522) );
  OA22X1 U802 ( .IN1(n786), .IN2(n535), .IN3(n806), .IN4(n533), .Q(n527) );
  OA22X1 U803 ( .IN1(n808), .IN2(n534), .IN3(n802), .IN4(n532), .Q(n526) );
  AND2X1 U804 ( .IN1(n524), .IN2(n788), .Q(n538) );
  NAND3X0 U805 ( .IN1(n527), .IN2(n526), .IN3(n525), .QN(N353) );
  OA22X1 U806 ( .IN1(n776), .IN2(n535), .IN3(n786), .IN4(n533), .Q(n531) );
  OA22X1 U807 ( .IN1(n808), .IN2(n532), .IN3(n810), .IN4(n537), .Q(n530) );
  OR2X1 U808 ( .IN1(n534), .IN2(n806), .Q(n528) );
  NAND4X0 U809 ( .IN1(n531), .IN2(n530), .IN3(n529), .IN4(n528), .QN(N354) );
  OA22X1 U810 ( .IN1(n776), .IN2(n533), .IN3(n806), .IN4(n532), .Q(n542) );
  OA22X1 U811 ( .IN1(n777), .IN2(n535), .IN3(n786), .IN4(n534), .Q(n541) );
  OA22X1 U812 ( .IN1(n802), .IN2(n537), .IN3(n810), .IN4(n536), .Q(n540) );
  NAND4X0 U813 ( .IN1(n542), .IN2(n541), .IN3(n540), .IN4(n539), .QN(N355) );
  AO22X1 U814 ( .IN1(n708), .IN2(exponent_factor_12[2]), .IN3(n821), .IN4(
        exponent_factor_21[2]), .Q(N36) );
  AO22X1 U815 ( .IN1(n708), .IN2(exponent_factor_12[3]), .IN3(n821), .IN4(
        exponent_factor_21[3]), .Q(N37) );
  AO22X1 U816 ( .IN1(n708), .IN2(exponent_factor_12[4]), .IN3(n821), .IN4(
        exponent_factor_21[4]), .Q(N38) );
  NAND4X0 U817 ( .IN1(n590), .IN2(n578), .IN3(n584), .IN4(n543), .QN(n544) );
  NOR4X0 U818 ( .IN1(input_factor_01[30]), .IN2(input_factor_01[23]), .IN3(
        n545), .IN4(n544), .QN(n554) );
  NOR4X0 U819 ( .IN1(input_factor_01[22]), .IN2(input_factor_01[21]), .IN3(
        input_factor_01[20]), .IN4(input_factor_01[17]), .QN(n553) );
  NOR4X0 U820 ( .IN1(input_factor_01[31]), .IN2(input_factor_01[25]), .IN3(
        input_factor_01[29]), .IN4(input_factor_01[16]), .QN(n552) );
  NAND4X0 U821 ( .IN1(n628), .IN2(n624), .IN3(n620), .IN4(n616), .QN(n550) );
  NAND4X0 U822 ( .IN1(n612), .IN2(n608), .IN3(n546), .IN4(n604), .QN(n549) );
  NAND4X0 U823 ( .IN1(n672), .IN2(n666), .IN3(n660), .IN4(n654), .QN(n548) );
  NAND4X0 U824 ( .IN1(n648), .IN2(n642), .IN3(n636), .IN4(n632), .QN(n547) );
  NOR4X0 U825 ( .IN1(n550), .IN2(n549), .IN3(n548), .IN4(n547), .QN(n551) );
  AOI22X1 U826 ( .IN1(input_factor_02[23]), .IN2(n22), .IN3(n710), .IN4(
        input_factor_01[23]), .QN(n569) );
  INVX0 U827 ( .INP(n778), .ZN(n555) );
  OA21X1 U828 ( .IN1(n761), .IN2(n556), .IN3(n555), .Q(n562) );
  NAND3X0 U829 ( .IN1(n557), .IN2(n701), .IN3(n702), .QN(n564) );
  OA21X1 U830 ( .IN1(n560), .IN2(n559), .IN3(n558), .Q(n561) );
  AOI22X1 U831 ( .IN1(n712), .IN2(add_output_exponent_w3[0]), .IN3(n711), 
        .IN4(add_output_exponent_w2[0]), .QN(n568) );
  INVX0 U832 ( .INP(n564), .ZN(n563) );
  AND4X1 U833 ( .IN1(n565), .IN2(n563), .IN3(n562), .IN4(n561), .Q(n714) );
  NAND4X0 U834 ( .IN1(n569), .IN2(n568), .IN3(n567), .IN4(n566), .QN(N380) );
  AOI22X1 U835 ( .IN1(input_factor_02[24]), .IN2(n22), .IN3(n710), .IN4(
        input_factor_01[24]), .QN(n573) );
  AOI22X1 U836 ( .IN1(n712), .IN2(add_output_exponent_w3[1]), .IN3(n711), 
        .IN4(add_output_exponent_w2[1]), .QN(n572) );
  NAND4X0 U837 ( .IN1(n573), .IN2(n572), .IN3(n571), .IN4(n570), .QN(N381) );
  AOI22X1 U838 ( .IN1(input_factor_02[25]), .IN2(n22), .IN3(n710), .IN4(
        input_factor_01[25]), .QN(n577) );
  AOI22X1 U839 ( .IN1(n712), .IN2(add_output_exponent_w3[2]), .IN3(n711), 
        .IN4(add_output_exponent_w2[2]), .QN(n576) );
  NAND4X0 U840 ( .IN1(n577), .IN2(n576), .IN3(n575), .IN4(n574), .QN(N382) );
  OA22X1 U841 ( .IN1(n579), .IN2(n702), .IN3(n701), .IN4(n578), .Q(n583) );
  AOI22X1 U842 ( .IN1(n712), .IN2(add_output_exponent_w3[3]), .IN3(n711), 
        .IN4(add_output_exponent_w2[3]), .QN(n582) );
  NAND4X0 U843 ( .IN1(n583), .IN2(n582), .IN3(n581), .IN4(n580), .QN(N383) );
  OA22X1 U844 ( .IN1(n585), .IN2(n702), .IN3(n701), .IN4(n584), .Q(n589) );
  AOI22X1 U845 ( .IN1(n712), .IN2(add_output_exponent_w3[4]), .IN3(n711), 
        .IN4(add_output_exponent_w2[4]), .QN(n588) );
  NAND4X0 U846 ( .IN1(n589), .IN2(n588), .IN3(n587), .IN4(n586), .QN(N384) );
  OA22X1 U847 ( .IN1(n591), .IN2(n702), .IN3(n701), .IN4(n590), .Q(n595) );
  AOI22X1 U848 ( .IN1(n712), .IN2(add_output_exponent_w3[5]), .IN3(n711), 
        .IN4(add_output_exponent_w2[5]), .QN(n594) );
  NAND4X0 U849 ( .IN1(n595), .IN2(n594), .IN3(n593), .IN4(n592), .QN(N385) );
  OA22X1 U850 ( .IN1(n597), .IN2(n702), .IN3(n701), .IN4(n596), .Q(n601) );
  AOI22X1 U851 ( .IN1(n712), .IN2(add_output_exponent_w3[6]), .IN3(n711), 
        .IN4(add_output_exponent_w2[6]), .QN(n600) );
  NAND4X0 U852 ( .IN1(n601), .IN2(n600), .IN3(n599), .IN4(n598), .QN(N386) );
  AO22X1 U854 ( .IN1(n710), .IN2(input_factor_01[30]), .IN3(n709), .IN4(
        add_output_exponent_w1[7]), .Q(n603) );
  AO22X1 U855 ( .IN1(n712), .IN2(add_output_exponent_w3[7]), .IN3(n711), .IN4(
        add_output_exponent_w2[7]), .Q(n602) );
  AO222X1 U856 ( .IN1(input_factor_02[0]), .IN2(n22), .IN3(input_factor_01[0]), 
        .IN4(n710), .IN5(n709), .IN6(pre_sig_res_01[0]), .Q(N388) );
  AOI22X1 U857 ( .IN1(n711), .IN2(pre_sig_res_02[1]), .IN3(n709), .IN4(
        pre_sig_res_01[1]), .QN(n607) );
  OA22X1 U858 ( .IN1(n605), .IN2(n702), .IN3(n701), .IN4(n604), .Q(n606) );
  AO22X1 U859 ( .IN1(n708), .IN2(exponent_factor_12[5]), .IN3(n821), .IN4(
        exponent_factor_21[5]), .Q(N39) );
  AOI22X1 U860 ( .IN1(n711), .IN2(pre_sig_res_02[2]), .IN3(n709), .IN4(
        pre_sig_res_01[2]), .QN(n611) );
  OA22X1 U861 ( .IN1(n609), .IN2(n702), .IN3(n701), .IN4(n608), .Q(n610) );
  AOI22X1 U862 ( .IN1(n711), .IN2(pre_sig_res_02[3]), .IN3(n709), .IN4(
        pre_sig_res_01[3]), .QN(n615) );
  OA22X1 U863 ( .IN1(n613), .IN2(n702), .IN3(n701), .IN4(n612), .Q(n614) );
  AOI22X1 U864 ( .IN1(n711), .IN2(pre_sig_res_02[4]), .IN3(n709), .IN4(
        pre_sig_res_01[4]), .QN(n619) );
  OA22X1 U865 ( .IN1(n617), .IN2(n702), .IN3(n701), .IN4(n616), .Q(n618) );
  AOI22X1 U866 ( .IN1(n711), .IN2(pre_sig_res_02[5]), .IN3(n709), .IN4(
        pre_sig_res_01[5]), .QN(n623) );
  OA22X1 U867 ( .IN1(n621), .IN2(n702), .IN3(n701), .IN4(n620), .Q(n622) );
  AOI22X1 U868 ( .IN1(n711), .IN2(pre_sig_res_02[6]), .IN3(n709), .IN4(
        pre_sig_res_01[6]), .QN(n627) );
  OA22X1 U869 ( .IN1(n625), .IN2(n702), .IN3(n701), .IN4(n624), .Q(n626) );
  AOI22X1 U870 ( .IN1(n711), .IN2(pre_sig_res_02[7]), .IN3(n709), .IN4(
        pre_sig_res_01[7]), .QN(n631) );
  OA22X1 U871 ( .IN1(n629), .IN2(n702), .IN3(n701), .IN4(n628), .Q(n630) );
  AOI22X1 U872 ( .IN1(n711), .IN2(pre_sig_res_02[8]), .IN3(n709), .IN4(
        pre_sig_res_01[8]), .QN(n635) );
  OA22X1 U873 ( .IN1(n633), .IN2(n702), .IN3(n701), .IN4(n632), .Q(n634) );
  OA22X1 U874 ( .IN1(n637), .IN2(n702), .IN3(n701), .IN4(n636), .Q(n641) );
  NAND4X0 U875 ( .IN1(n641), .IN2(n640), .IN3(n639), .IN4(n638), .QN(N397) );
  OA22X1 U876 ( .IN1(n643), .IN2(n702), .IN3(n701), .IN4(n642), .Q(n647) );
  NAND4X0 U877 ( .IN1(n647), .IN2(n646), .IN3(n645), .IN4(n644), .QN(N398) );
  OA22X1 U878 ( .IN1(n649), .IN2(n702), .IN3(n701), .IN4(n648), .Q(n653) );
  NAND4X0 U879 ( .IN1(n653), .IN2(n652), .IN3(n651), .IN4(n650), .QN(N399) );
  AO22X1 U880 ( .IN1(n708), .IN2(exponent_factor_12[6]), .IN3(n821), .IN4(
        exponent_factor_21[6]), .Q(N40) );
  OA22X1 U881 ( .IN1(n655), .IN2(n702), .IN3(n701), .IN4(n654), .Q(n659) );
  NAND4X0 U882 ( .IN1(n659), .IN2(n658), .IN3(n657), .IN4(n656), .QN(N400) );
  OA22X1 U883 ( .IN1(n661), .IN2(n702), .IN3(n701), .IN4(n660), .Q(n665) );
  NAND4X0 U884 ( .IN1(n665), .IN2(n664), .IN3(n663), .IN4(n662), .QN(N401) );
  OA22X1 U885 ( .IN1(n667), .IN2(n702), .IN3(n701), .IN4(n666), .Q(n671) );
  NAND4X0 U886 ( .IN1(n671), .IN2(n670), .IN3(n669), .IN4(n668), .QN(N402) );
  OA22X1 U887 ( .IN1(n673), .IN2(n702), .IN3(n701), .IN4(n672), .Q(n677) );
  NAND4X0 U888 ( .IN1(n677), .IN2(n676), .IN3(n675), .IN4(n674), .QN(N403) );
  OA22X1 U889 ( .IN1(n679), .IN2(n702), .IN3(n701), .IN4(n678), .Q(n683) );
  AOI22X1 U890 ( .IN1(n712), .IN2(pre_sig_res_03[16]), .IN3(n711), .IN4(
        pre_sig_res_02[16]), .QN(n682) );
  NAND4X0 U891 ( .IN1(n683), .IN2(n682), .IN3(n681), .IN4(n680), .QN(N404) );
  OA22X1 U892 ( .IN1(n685), .IN2(n702), .IN3(n701), .IN4(n684), .Q(n689) );
  AOI22X1 U893 ( .IN1(n712), .IN2(pre_sig_res_03[17]), .IN3(n711), .IN4(
        pre_sig_res_02[17]), .QN(n688) );
  NAND4X0 U894 ( .IN1(n689), .IN2(n688), .IN3(n687), .IN4(n686), .QN(N405) );
  AO22X1 U895 ( .IN1(n710), .IN2(input_factor_01[18]), .IN3(n709), .IN4(
        pre_sig_res_01[18]), .Q(n691) );
  AO22X1 U896 ( .IN1(n712), .IN2(pre_sig_res_03[18]), .IN3(n711), .IN4(
        pre_sig_res_02[18]), .Q(n690) );
  AO22X1 U897 ( .IN1(n710), .IN2(input_factor_01[19]), .IN3(n709), .IN4(
        pre_sig_res_01[19]), .Q(n693) );
  AO22X1 U898 ( .IN1(n712), .IN2(pre_sig_res_03[19]), .IN3(n711), .IN4(
        pre_sig_res_02[19]), .Q(n692) );
  OA22X1 U899 ( .IN1(n695), .IN2(n702), .IN3(n701), .IN4(n694), .Q(n699) );
  AOI22X1 U900 ( .IN1(n712), .IN2(pre_sig_res_03[20]), .IN3(n711), .IN4(
        pre_sig_res_02[20]), .QN(n698) );
  NAND4X0 U901 ( .IN1(n699), .IN2(n698), .IN3(n697), .IN4(n696), .QN(N408) );
  OA22X1 U902 ( .IN1(n703), .IN2(n702), .IN3(n701), .IN4(n700), .Q(n707) );
  AOI22X1 U903 ( .IN1(n712), .IN2(pre_sig_res_03[21]), .IN3(n711), .IN4(
        pre_sig_res_02[21]), .QN(n706) );
  NAND4X0 U904 ( .IN1(n707), .IN2(n706), .IN3(n705), .IN4(n704), .QN(N409) );
  AO22X1 U905 ( .IN1(n708), .IN2(exponent_factor_12[7]), .IN3(n821), .IN4(
        exponent_factor_21[7]), .Q(N41) );
  AO22X1 U906 ( .IN1(n710), .IN2(input_factor_01[22]), .IN3(n709), .IN4(
        pre_sig_res_01[22]), .Q(n715) );
  AO22X1 U907 ( .IN1(n712), .IN2(pre_sig_res_03[22]), .IN3(n711), .IN4(
        pre_sig_res_02[22]), .Q(n713) );
  NOR2X0 U908 ( .IN1(n848), .IN2(n716), .QN(n817) );
  NOR2X0 U909 ( .IN1(n717), .IN2(n848), .QN(n819) );
  OA22X1 U910 ( .IN1(n729), .IN2(n807), .IN3(n718), .IN4(n805), .Q(n728) );
  OA22X1 U911 ( .IN1(n745), .IN2(n811), .IN3(n769), .IN4(n778), .Q(n722) );
  INVX0 U912 ( .INP(rst_n), .ZN(n820) );
  NAND3X0 U913 ( .IN1(n720), .IN2(n740), .IN3(n719), .QN(n721) );
  OA22X1 U914 ( .IN1(n848), .IN2(n722), .IN3(n820), .IN4(n721), .Q(n727) );
  NAND4X0 U915 ( .IN1(n728), .IN2(n727), .IN3(n726), .IN4(n725), .QN(n847) );
  OA22X1 U916 ( .IN1(n729), .IN2(n805), .IN3(n737), .IN4(n807), .Q(n736) );
  OA22X1 U917 ( .IN1(n769), .IN2(n785), .IN3(n777), .IN4(n778), .Q(n731) );
  OA22X1 U918 ( .IN1(n761), .IN2(n794), .IN3(n753), .IN4(n811), .Q(n730) );
  AO21X1 U919 ( .IN1(n731), .IN2(n730), .IN3(n848), .Q(n735) );
  NAND4X0 U920 ( .IN1(n736), .IN2(n735), .IN3(n734), .IN4(n733), .QN(n846) );
  OA22X1 U921 ( .IN1(n737), .IN2(n805), .IN3(n745), .IN4(n807), .Q(n744) );
  OA22X1 U922 ( .IN1(n777), .IN2(n785), .IN3(n776), .IN4(n778), .Q(n739) );
  OA22X1 U923 ( .IN1(n761), .IN2(n811), .IN3(n769), .IN4(n794), .Q(n738) );
  AO21X1 U924 ( .IN1(n739), .IN2(n738), .IN3(n848), .Q(n743) );
  NAND4X0 U925 ( .IN1(n744), .IN2(n743), .IN3(n742), .IN4(n741), .QN(n845) );
  OA22X1 U926 ( .IN1(n745), .IN2(n805), .IN3(n753), .IN4(n807), .Q(n752) );
  OA22X1 U927 ( .IN1(n776), .IN2(n785), .IN3(n786), .IN4(n778), .Q(n747) );
  OA22X1 U928 ( .IN1(n769), .IN2(n811), .IN3(n777), .IN4(n794), .Q(n746) );
  AO21X1 U929 ( .IN1(n747), .IN2(n746), .IN3(n848), .Q(n751) );
  NAND4X0 U930 ( .IN1(n752), .IN2(n751), .IN3(n750), .IN4(n749), .QN(n844) );
  OA22X1 U931 ( .IN1(n761), .IN2(n807), .IN3(n753), .IN4(n805), .Q(n760) );
  OA22X1 U932 ( .IN1(n786), .IN2(n785), .IN3(n806), .IN4(n778), .Q(n755) );
  OA22X1 U933 ( .IN1(n777), .IN2(n811), .IN3(n776), .IN4(n794), .Q(n754) );
  AO21X1 U934 ( .IN1(n755), .IN2(n754), .IN3(n848), .Q(n759) );
  NAND4X0 U935 ( .IN1(n760), .IN2(n759), .IN3(n758), .IN4(n757), .QN(n843) );
  OA22X1 U936 ( .IN1(n761), .IN2(n805), .IN3(n769), .IN4(n807), .Q(n768) );
  OA22X1 U937 ( .IN1(n808), .IN2(n778), .IN3(n806), .IN4(n785), .Q(n763) );
  OA22X1 U938 ( .IN1(n776), .IN2(n811), .IN3(n786), .IN4(n794), .Q(n762) );
  AO21X1 U939 ( .IN1(n763), .IN2(n762), .IN3(n848), .Q(n767) );
  NAND4X0 U940 ( .IN1(n768), .IN2(n767), .IN3(n766), .IN4(n765), .QN(n842) );
  OA22X1 U941 ( .IN1(n769), .IN2(n805), .IN3(n777), .IN4(n807), .Q(n775) );
  OA22X1 U942 ( .IN1(n808), .IN2(n785), .IN3(n802), .IN4(n778), .Q(n771) );
  OA22X1 U943 ( .IN1(n786), .IN2(n811), .IN3(n806), .IN4(n794), .Q(n770) );
  AO21X1 U944 ( .IN1(n771), .IN2(n770), .IN3(n848), .Q(n774) );
  NAND4X0 U945 ( .IN1(n775), .IN2(n774), .IN3(n773), .IN4(n772), .QN(n841) );
  OA22X1 U946 ( .IN1(n777), .IN2(n805), .IN3(n776), .IN4(n807), .Q(n784) );
  OA22X1 U947 ( .IN1(n802), .IN2(n785), .IN3(n810), .IN4(n778), .Q(n780) );
  OA22X1 U948 ( .IN1(n808), .IN2(n794), .IN3(n806), .IN4(n811), .Q(n779) );
  AO21X1 U949 ( .IN1(n780), .IN2(n779), .IN3(n848), .Q(n783) );
  NAND4X0 U950 ( .IN1(n784), .IN2(n783), .IN3(n782), .IN4(n781), .QN(n840) );
  OA222X1 U951 ( .IN1(n811), .IN2(n808), .IN3(n785), .IN4(n810), .IN5(n794), 
        .IN6(n802), .Q(n787) );
  OA22X1 U952 ( .IN1(n848), .IN2(n787), .IN3(n786), .IN4(n807), .Q(n793) );
  NAND4X0 U953 ( .IN1(n793), .IN2(n792), .IN3(n791), .IN4(n790), .QN(n839) );
  OA22X1 U954 ( .IN1(n802), .IN2(n811), .IN3(n810), .IN4(n794), .Q(n795) );
  OA22X1 U955 ( .IN1(n806), .IN2(n807), .IN3(n795), .IN4(n820), .Q(n801) );
  NAND4X0 U956 ( .IN1(n801), .IN2(n800), .IN3(n799), .IN4(n798), .QN(n838) );
  AOI22X1 U957 ( .IN1(pre_sig_res_03[11]), .IN2(n820), .IN3(n809), .IN4(n818), 
        .QN(n804) );
  OA22X1 U958 ( .IN1(n808), .IN2(n805), .IN3(n802), .IN4(n807), .Q(n803) );
  OA22X1 U959 ( .IN1(n808), .IN2(n807), .IN3(n806), .IN4(n805), .Q(n815) );
  OR3X1 U960 ( .IN1(n811), .IN2(n820), .IN3(n810), .Q(n813) );
  NAND4X0 U961 ( .IN1(n815), .IN2(n814), .IN3(n813), .IN4(n812), .QN(n836) );
  AO222X1 U962 ( .IN1(n818), .IN2(n817), .IN3(n816), .IN4(n819), .IN5(n820), 
        .IN6(pre_sig_res_03[10]), .Q(n835) );
  AO22X1 U963 ( .IN1(pre_sig_res_03[9]), .IN2(n820), .IN3(n819), .IN4(n818), 
        .Q(n834) );
  AND2X1 U964 ( .IN1(n821), .IN2(rst_n), .Q(n823) );
  AO222X1 U965 ( .IN1(input_factor_02[23]), .IN2(n823), .IN3(
        input_factor_01[23]), .IN4(n822), .IN5(larger_exponent[0]), .IN6(n848), 
        .Q(n833) );
  AO222X1 U966 ( .IN1(input_factor_02[24]), .IN2(n823), .IN3(
        input_factor_01[24]), .IN4(n822), .IN5(n848), .IN6(larger_exponent[1]), 
        .Q(n832) );
  AO222X1 U967 ( .IN1(input_factor_02[25]), .IN2(n823), .IN3(
        input_factor_01[25]), .IN4(n822), .IN5(n848), .IN6(larger_exponent[2]), 
        .Q(n831) );
  AO222X1 U968 ( .IN1(input_factor_02[26]), .IN2(n823), .IN3(
        input_factor_01[26]), .IN4(n822), .IN5(n848), .IN6(larger_exponent[3]), 
        .Q(n830) );
  AO222X1 U969 ( .IN1(input_factor_02[27]), .IN2(n823), .IN3(
        input_factor_01[27]), .IN4(n822), .IN5(n848), .IN6(larger_exponent[4]), 
        .Q(n829) );
  AO222X1 U970 ( .IN1(input_factor_02[28]), .IN2(n823), .IN3(
        input_factor_01[28]), .IN4(n822), .IN5(n848), .IN6(larger_exponent[5]), 
        .Q(n828) );
  AO222X1 U971 ( .IN1(input_factor_02[29]), .IN2(n823), .IN3(
        input_factor_01[29]), .IN4(n822), .IN5(n848), .IN6(larger_exponent[6]), 
        .Q(n827) );
endmodule


module cla51squ_1 ( out, a, b );
  output [50:0] out;
  input [50:0] a;
  input [50:0] b;
  wire   intadd_1_CI, intadd_1_n24, intadd_1_n23, intadd_1_n22, intadd_1_n21,
         intadd_1_n20, intadd_1_n19, intadd_1_n18, intadd_1_n17, intadd_1_n16,
         intadd_1_n15, intadd_1_n14, intadd_1_n13, intadd_1_n12, intadd_1_n11,
         intadd_1_n10, intadd_1_n9, intadd_1_n8, intadd_1_n7, intadd_1_n6,
         intadd_1_n5, intadd_1_n4, intadd_1_n3, intadd_1_n2, intadd_1_n1, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14;

  FADDX1 intadd_1_U25 ( .A(b[23]), .B(a[23]), .CI(intadd_1_CI), .CO(
        intadd_1_n24), .S(out[23]) );
  FADDX1 intadd_1_U24 ( .A(b[24]), .B(a[24]), .CI(intadd_1_n24), .CO(
        intadd_1_n23), .S(out[24]) );
  FADDX1 intadd_1_U23 ( .A(b[25]), .B(a[25]), .CI(intadd_1_n23), .CO(
        intadd_1_n22), .S(out[25]) );
  FADDX1 intadd_1_U22 ( .A(b[26]), .B(a[26]), .CI(intadd_1_n22), .CO(
        intadd_1_n21), .S(out[26]) );
  FADDX1 intadd_1_U21 ( .A(b[27]), .B(a[27]), .CI(intadd_1_n21), .CO(
        intadd_1_n20), .S(out[27]) );
  FADDX1 intadd_1_U20 ( .A(b[28]), .B(a[28]), .CI(intadd_1_n20), .CO(
        intadd_1_n19), .S(out[28]) );
  FADDX1 intadd_1_U19 ( .A(b[29]), .B(a[29]), .CI(intadd_1_n19), .CO(
        intadd_1_n18), .S(out[29]) );
  FADDX1 intadd_1_U18 ( .A(b[30]), .B(a[30]), .CI(intadd_1_n18), .CO(
        intadd_1_n17), .S(out[30]) );
  FADDX1 intadd_1_U17 ( .A(b[31]), .B(a[31]), .CI(intadd_1_n17), .CO(
        intadd_1_n16), .S(out[31]) );
  FADDX1 intadd_1_U16 ( .A(b[32]), .B(a[32]), .CI(intadd_1_n16), .CO(
        intadd_1_n15), .S(out[32]) );
  FADDX1 intadd_1_U15 ( .A(b[33]), .B(a[33]), .CI(intadd_1_n15), .CO(
        intadd_1_n14), .S(out[33]) );
  FADDX1 intadd_1_U14 ( .A(b[34]), .B(a[34]), .CI(intadd_1_n14), .CO(
        intadd_1_n13), .S(out[34]) );
  FADDX1 intadd_1_U13 ( .A(b[35]), .B(a[35]), .CI(intadd_1_n13), .CO(
        intadd_1_n12), .S(out[35]) );
  FADDX1 intadd_1_U12 ( .A(b[36]), .B(a[36]), .CI(intadd_1_n12), .CO(
        intadd_1_n11), .S(out[36]) );
  FADDX1 intadd_1_U11 ( .A(b[37]), .B(a[37]), .CI(intadd_1_n11), .CO(
        intadd_1_n10), .S(out[37]) );
  FADDX1 intadd_1_U10 ( .A(b[38]), .B(a[38]), .CI(intadd_1_n10), .CO(
        intadd_1_n9), .S(out[38]) );
  FADDX1 intadd_1_U9 ( .A(b[39]), .B(a[39]), .CI(intadd_1_n9), .CO(intadd_1_n8), .S(out[39]) );
  FADDX1 intadd_1_U8 ( .A(b[40]), .B(a[40]), .CI(intadd_1_n8), .CO(intadd_1_n7), .S(out[40]) );
  FADDX1 intadd_1_U7 ( .A(b[41]), .B(a[41]), .CI(intadd_1_n7), .CO(intadd_1_n6), .S(out[41]) );
  FADDX1 intadd_1_U6 ( .A(b[42]), .B(a[42]), .CI(intadd_1_n6), .CO(intadd_1_n5), .S(out[42]) );
  FADDX1 intadd_1_U5 ( .A(b[43]), .B(a[43]), .CI(intadd_1_n5), .CO(intadd_1_n4), .S(out[43]) );
  FADDX1 intadd_1_U4 ( .A(b[44]), .B(a[44]), .CI(intadd_1_n4), .CO(intadd_1_n3), .S(out[44]) );
  FADDX1 intadd_1_U3 ( .A(b[45]), .B(a[45]), .CI(intadd_1_n3), .CO(intadd_1_n2), .S(out[45]) );
  FADDX1 intadd_1_U2 ( .A(b[46]), .B(a[46]), .CI(intadd_1_n2), .CO(intadd_1_n1), .S(out[46]) );
  OA21X1 U2 ( .IN1(b[9]), .IN2(a[9]), .IN3(a[8]), .Q(n1) );
  AO22X1 U3 ( .IN1(b[9]), .IN2(a[9]), .IN3(b[8]), .IN4(n1), .Q(n2) );
  AO222X1 U4 ( .IN1(b[10]), .IN2(a[10]), .IN3(b[10]), .IN4(n2), .IN5(a[10]), 
        .IN6(n2), .Q(n3) );
  AO222X1 U5 ( .IN1(b[11]), .IN2(a[11]), .IN3(b[11]), .IN4(n3), .IN5(a[11]), 
        .IN6(n3), .Q(n4) );
  AO222X1 U6 ( .IN1(b[12]), .IN2(a[12]), .IN3(b[12]), .IN4(n4), .IN5(a[12]), 
        .IN6(n4), .Q(n5) );
  AO222X1 U7 ( .IN1(b[13]), .IN2(a[13]), .IN3(b[13]), .IN4(n5), .IN5(a[13]), 
        .IN6(n5), .Q(n6) );
  AO222X1 U8 ( .IN1(b[14]), .IN2(a[14]), .IN3(b[14]), .IN4(n6), .IN5(a[14]), 
        .IN6(n6), .Q(n7) );
  AO222X1 U9 ( .IN1(b[15]), .IN2(a[15]), .IN3(b[15]), .IN4(n7), .IN5(a[15]), 
        .IN6(n7), .Q(n8) );
  AO222X1 U10 ( .IN1(b[16]), .IN2(a[16]), .IN3(b[16]), .IN4(n8), .IN5(a[16]), 
        .IN6(n8), .Q(n9) );
  AO222X1 U11 ( .IN1(b[17]), .IN2(a[17]), .IN3(b[17]), .IN4(n9), .IN5(a[17]), 
        .IN6(n9), .Q(n10) );
  AO222X1 U12 ( .IN1(b[18]), .IN2(a[18]), .IN3(b[18]), .IN4(n10), .IN5(a[18]), 
        .IN6(n10), .Q(n11) );
  AO222X1 U13 ( .IN1(b[19]), .IN2(a[19]), .IN3(b[19]), .IN4(n11), .IN5(a[19]), 
        .IN6(n11), .Q(n12) );
  AO222X1 U14 ( .IN1(b[20]), .IN2(a[20]), .IN3(b[20]), .IN4(n12), .IN5(a[20]), 
        .IN6(n12), .Q(n13) );
  AO222X1 U15 ( .IN1(b[21]), .IN2(a[21]), .IN3(b[21]), .IN4(n13), .IN5(a[21]), 
        .IN6(n13), .Q(n14) );
  AO222X1 U16 ( .IN1(b[22]), .IN2(a[22]), .IN3(b[22]), .IN4(n14), .IN5(a[22]), 
        .IN6(n14), .Q(intadd_1_CI) );
  XOR3X1 U17 ( .IN1(intadd_1_n1), .IN2(a[47]), .IN3(b[47]), .Q(out[47]) );
endmodule


module csa51squ_1 ( sumout, in1, in2, in3, cout_50_, cout_49_, cout_48_, 
        cout_47_, cout_46_, cout_44_, cout_42_, cout_40_, cout_38_, cout_36_, 
        cout_34_, cout_32_, cout_30_, cout_28_, cout_27_, cout_7__BAR, cout_6_, 
        cout_5_, cout_4_, cout_3_, cout_2_, cout_1_, cout_0_, cout_8__BAR, 
        cout_9__BAR, cout_10__BAR, cout_11__BAR, cout_12__BAR, cout_13__BAR, 
        cout_14__BAR, cout_15__BAR, cout_16__BAR, cout_17__BAR, cout_18__BAR, 
        cout_19__BAR, cout_20__BAR, cout_21__BAR, cout_22__BAR, cout_23__BAR, 
        cout_24__BAR, cout_25__BAR, cout_26__BAR, cout_29__BAR, cout_31__BAR, 
        cout_33__BAR, cout_35__BAR, cout_37__BAR, cout_39__BAR, cout_41__BAR, 
        cout_43__BAR, cout_45__BAR );
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  output cout_50_, cout_49_, cout_48_, cout_47_, cout_46_, cout_44_, cout_42_,
         cout_40_, cout_38_, cout_36_, cout_34_, cout_32_, cout_30_, cout_28_,
         cout_27_, cout_7__BAR, cout_6_, cout_5_, cout_4_, cout_3_, cout_2_,
         cout_1_, cout_0_, cout_8__BAR, cout_9__BAR, cout_10__BAR,
         cout_11__BAR, cout_12__BAR, cout_13__BAR, cout_14__BAR, cout_15__BAR,
         cout_16__BAR, cout_17__BAR, cout_18__BAR, cout_19__BAR, cout_20__BAR,
         cout_21__BAR, cout_22__BAR, cout_23__BAR, cout_24__BAR, cout_25__BAR,
         cout_26__BAR, cout_29__BAR, cout_31__BAR, cout_33__BAR, cout_35__BAR,
         cout_37__BAR, cout_39__BAR, cout_41__BAR, cout_43__BAR, cout_45__BAR;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11;

  NAND2X0 U1 ( .IN1(in2[8]), .IN2(in1[8]), .QN(cout_8__BAR) );
  NAND2X0 U2 ( .IN1(in2[9]), .IN2(in1[9]), .QN(cout_9__BAR) );
  NAND2X0 U3 ( .IN1(in2[10]), .IN2(in1[10]), .QN(cout_10__BAR) );
  NAND2X0 U4 ( .IN1(in2[11]), .IN2(in1[11]), .QN(cout_11__BAR) );
  NAND2X0 U5 ( .IN1(in2[12]), .IN2(in1[12]), .QN(cout_12__BAR) );
  NAND2X0 U6 ( .IN1(in2[13]), .IN2(in1[13]), .QN(cout_13__BAR) );
  NAND2X0 U7 ( .IN1(in2[14]), .IN2(in1[14]), .QN(cout_14__BAR) );
  NAND2X0 U8 ( .IN1(in2[15]), .IN2(in1[15]), .QN(cout_15__BAR) );
  NAND2X0 U9 ( .IN1(in2[16]), .IN2(in1[16]), .QN(cout_16__BAR) );
  NAND2X0 U10 ( .IN1(in2[17]), .IN2(in1[17]), .QN(cout_17__BAR) );
  NAND2X0 U11 ( .IN1(in2[18]), .IN2(in1[18]), .QN(cout_18__BAR) );
  NAND2X0 U12 ( .IN1(in2[19]), .IN2(in1[19]), .QN(cout_19__BAR) );
  NAND2X0 U13 ( .IN1(in2[20]), .IN2(in1[20]), .QN(cout_20__BAR) );
  NAND2X0 U14 ( .IN1(in2[21]), .IN2(in1[21]), .QN(cout_21__BAR) );
  NAND2X0 U15 ( .IN1(in2[22]), .IN2(in1[22]), .QN(cout_22__BAR) );
  NAND2X0 U16 ( .IN1(in2[23]), .IN2(in1[23]), .QN(cout_23__BAR) );
  NAND2X0 U17 ( .IN1(in2[24]), .IN2(in1[24]), .QN(cout_24__BAR) );
  NAND2X0 U18 ( .IN1(in2[25]), .IN2(in1[25]), .QN(cout_25__BAR) );
  NAND2X0 U19 ( .IN1(in2[26]), .IN2(in1[26]), .QN(cout_26__BAR) );
  NAND2X0 U20 ( .IN1(in2[29]), .IN2(in1[29]), .QN(cout_29__BAR) );
  NAND2X0 U21 ( .IN1(in2[31]), .IN2(in1[31]), .QN(cout_31__BAR) );
  NAND2X0 U22 ( .IN1(in2[33]), .IN2(in1[33]), .QN(cout_33__BAR) );
  NAND2X0 U23 ( .IN1(in2[35]), .IN2(in1[35]), .QN(cout_35__BAR) );
  NAND2X0 U24 ( .IN1(in2[37]), .IN2(in1[37]), .QN(cout_37__BAR) );
  NAND2X0 U25 ( .IN1(in2[39]), .IN2(in1[39]), .QN(cout_39__BAR) );
  NAND2X0 U26 ( .IN1(in2[41]), .IN2(in1[41]), .QN(cout_41__BAR) );
  NAND2X0 U27 ( .IN1(in2[43]), .IN2(in1[43]), .QN(cout_43__BAR) );
  NAND2X0 U28 ( .IN1(in2[45]), .IN2(in1[45]), .QN(cout_45__BAR) );
  NAND2X0 U29 ( .IN1(in2[7]), .IN2(in1[7]), .QN(cout_7__BAR) );
  NAND2X0 U30 ( .IN1(n1), .IN2(cout_27_), .QN(sumout[27]) );
  NAND2X0 U31 ( .IN1(in1[27]), .IN2(in2[27]), .QN(n1) );
  NAND2X0 U32 ( .IN1(n2), .IN2(cout_28_), .QN(sumout[28]) );
  NAND2X0 U33 ( .IN1(in1[28]), .IN2(in2[28]), .QN(n2) );
  NAND2X0 U34 ( .IN1(n3), .IN2(cout_30_), .QN(sumout[30]) );
  NAND2X0 U35 ( .IN1(in1[30]), .IN2(in2[30]), .QN(n3) );
  NAND2X0 U36 ( .IN1(n4), .IN2(cout_32_), .QN(sumout[32]) );
  NAND2X0 U37 ( .IN1(in1[32]), .IN2(in2[32]), .QN(n4) );
  NAND2X0 U38 ( .IN1(n5), .IN2(cout_34_), .QN(sumout[34]) );
  NAND2X0 U39 ( .IN1(in1[34]), .IN2(in2[34]), .QN(n5) );
  NAND2X0 U40 ( .IN1(n6), .IN2(cout_36_), .QN(sumout[36]) );
  NAND2X0 U41 ( .IN1(in1[36]), .IN2(in2[36]), .QN(n6) );
  NAND2X0 U42 ( .IN1(n7), .IN2(cout_38_), .QN(sumout[38]) );
  NAND2X0 U43 ( .IN1(in1[38]), .IN2(in2[38]), .QN(n7) );
  NAND2X0 U44 ( .IN1(n8), .IN2(cout_40_), .QN(sumout[40]) );
  NAND2X0 U45 ( .IN1(in1[40]), .IN2(in2[40]), .QN(n8) );
  NAND2X0 U46 ( .IN1(n9), .IN2(cout_42_), .QN(sumout[42]) );
  NAND2X0 U47 ( .IN1(in1[42]), .IN2(in2[42]), .QN(n9) );
  NAND2X0 U48 ( .IN1(n10), .IN2(cout_44_), .QN(sumout[44]) );
  NAND2X0 U49 ( .IN1(in1[44]), .IN2(in2[44]), .QN(n10) );
  NAND2X0 U50 ( .IN1(n11), .IN2(cout_46_), .QN(sumout[46]) );
  NAND2X0 U51 ( .IN1(in1[46]), .IN2(in2[46]), .QN(n11) );
  OR2X1 U52 ( .IN1(in2[27]), .IN2(in1[27]), .Q(cout_27_) );
  OR2X1 U53 ( .IN1(in2[28]), .IN2(in1[28]), .Q(cout_28_) );
  OR2X1 U54 ( .IN1(in2[30]), .IN2(in1[30]), .Q(cout_30_) );
  OR2X1 U55 ( .IN1(in2[32]), .IN2(in1[32]), .Q(cout_32_) );
  OR2X1 U56 ( .IN1(in2[34]), .IN2(in1[34]), .Q(cout_34_) );
  OR2X1 U57 ( .IN1(in2[36]), .IN2(in1[36]), .Q(cout_36_) );
  OR2X1 U58 ( .IN1(in2[38]), .IN2(in1[38]), .Q(cout_38_) );
  OR2X1 U59 ( .IN1(in2[40]), .IN2(in1[40]), .Q(cout_40_) );
  OR2X1 U60 ( .IN1(in2[42]), .IN2(in1[42]), .Q(cout_42_) );
  OR2X1 U61 ( .IN1(in2[44]), .IN2(in1[44]), .Q(cout_44_) );
  OR2X1 U62 ( .IN1(in2[46]), .IN2(in1[46]), .Q(cout_46_) );
  OA21X1 U63 ( .IN1(in2[8]), .IN2(in1[8]), .IN3(cout_8__BAR), .Q(sumout[8]) );
  OA21X1 U64 ( .IN1(in2[9]), .IN2(in1[9]), .IN3(cout_9__BAR), .Q(sumout[9]) );
  OA21X1 U65 ( .IN1(in2[10]), .IN2(in1[10]), .IN3(cout_10__BAR), .Q(sumout[10]) );
  OA21X1 U66 ( .IN1(in2[11]), .IN2(in1[11]), .IN3(cout_11__BAR), .Q(sumout[11]) );
  OA21X1 U67 ( .IN1(in2[12]), .IN2(in1[12]), .IN3(cout_12__BAR), .Q(sumout[12]) );
  OA21X1 U68 ( .IN1(in2[13]), .IN2(in1[13]), .IN3(cout_13__BAR), .Q(sumout[13]) );
  OA21X1 U69 ( .IN1(in2[14]), .IN2(in1[14]), .IN3(cout_14__BAR), .Q(sumout[14]) );
  OA21X1 U70 ( .IN1(in2[15]), .IN2(in1[15]), .IN3(cout_15__BAR), .Q(sumout[15]) );
  OA21X1 U71 ( .IN1(in2[16]), .IN2(in1[16]), .IN3(cout_16__BAR), .Q(sumout[16]) );
  OA21X1 U72 ( .IN1(in2[17]), .IN2(in1[17]), .IN3(cout_17__BAR), .Q(sumout[17]) );
  OA21X1 U73 ( .IN1(in2[18]), .IN2(in1[18]), .IN3(cout_18__BAR), .Q(sumout[18]) );
  OA21X1 U74 ( .IN1(in2[19]), .IN2(in1[19]), .IN3(cout_19__BAR), .Q(sumout[19]) );
  OA21X1 U75 ( .IN1(in2[20]), .IN2(in1[20]), .IN3(cout_20__BAR), .Q(sumout[20]) );
  OA21X1 U76 ( .IN1(in2[21]), .IN2(in1[21]), .IN3(cout_21__BAR), .Q(sumout[21]) );
  OA21X1 U77 ( .IN1(in2[22]), .IN2(in1[22]), .IN3(cout_22__BAR), .Q(sumout[22]) );
  OA21X1 U78 ( .IN1(in2[23]), .IN2(in1[23]), .IN3(cout_23__BAR), .Q(sumout[23]) );
  OA21X1 U79 ( .IN1(in2[24]), .IN2(in1[24]), .IN3(cout_24__BAR), .Q(sumout[24]) );
  OA21X1 U80 ( .IN1(in2[25]), .IN2(in1[25]), .IN3(cout_25__BAR), .Q(sumout[25]) );
  OA21X1 U81 ( .IN1(in2[26]), .IN2(in1[26]), .IN3(cout_26__BAR), .Q(sumout[26]) );
  OA21X1 U82 ( .IN1(in2[29]), .IN2(in1[29]), .IN3(cout_29__BAR), .Q(sumout[29]) );
  OA21X1 U83 ( .IN1(in2[31]), .IN2(in1[31]), .IN3(cout_31__BAR), .Q(sumout[31]) );
  OA21X1 U84 ( .IN1(in2[33]), .IN2(in1[33]), .IN3(cout_33__BAR), .Q(sumout[33]) );
  OA21X1 U85 ( .IN1(in2[35]), .IN2(in1[35]), .IN3(cout_35__BAR), .Q(sumout[35]) );
  OA21X1 U86 ( .IN1(in2[37]), .IN2(in1[37]), .IN3(cout_37__BAR), .Q(sumout[37]) );
  OA21X1 U87 ( .IN1(in2[39]), .IN2(in1[39]), .IN3(cout_39__BAR), .Q(sumout[39]) );
  OA21X1 U88 ( .IN1(in2[41]), .IN2(in1[41]), .IN3(cout_41__BAR), .Q(sumout[41]) );
  OA21X1 U89 ( .IN1(in2[43]), .IN2(in1[43]), .IN3(cout_43__BAR), .Q(sumout[43]) );
  OA21X1 U90 ( .IN1(in2[45]), .IN2(in1[45]), .IN3(cout_45__BAR), .Q(sumout[45]) );
  XOR2X1 U91 ( .IN1(in1[47]), .IN2(in2[47]), .Q(sumout[47]) );
endmodule


module csa51squ_2 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;


  AO222X1 U1 ( .IN1(in2[6]), .IN2(in3[6]), .IN3(in2[6]), .IN4(in1[6]), .IN5(
        in3[6]), .IN6(in1[6]), .Q(cout[6]) );
  FADDX1 U2 ( .A(in1[10]), .B(in2[10]), .CI(in3[10]), .CO(cout[10]), .S(
        sumout[10]) );
  FADDX1 U3 ( .A(in1[11]), .B(in2[11]), .CI(in3[11]), .CO(cout[11]), .S(
        sumout[11]) );
  FADDX1 U4 ( .A(in1[12]), .B(in2[12]), .CI(in3[12]), .CO(cout[12]), .S(
        sumout[12]) );
  FADDX1 U5 ( .A(in1[13]), .B(in2[13]), .CI(in3[13]), .CO(cout[13]), .S(
        sumout[13]) );
  FADDX1 U6 ( .A(in1[14]), .B(in2[14]), .CI(in3[14]), .CO(cout[14]), .S(
        sumout[14]) );
  FADDX1 U7 ( .A(in1[15]), .B(in2[15]), .CI(in3[15]), .CO(cout[15]), .S(
        sumout[15]) );
  FADDX1 U8 ( .A(in1[16]), .B(in2[16]), .CI(in3[16]), .CO(cout[16]), .S(
        sumout[16]) );
  FADDX1 U9 ( .A(in1[17]), .B(in2[17]), .CI(in3[17]), .CO(cout[17]), .S(
        sumout[17]) );
  FADDX1 U10 ( .A(in1[18]), .B(in2[18]), .CI(in3[18]), .CO(cout[18]), .S(
        sumout[18]) );
  FADDX1 U11 ( .A(in1[19]), .B(in2[19]), .CI(in3[19]), .CO(cout[19]), .S(
        sumout[19]) );
  FADDX1 U12 ( .A(in1[20]), .B(in2[20]), .CI(in3[20]), .CO(cout[20]), .S(
        sumout[20]) );
  FADDX1 U13 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U14 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U15 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U16 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U17 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U18 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U19 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U20 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U21 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U22 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U23 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U24 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
  FADDX1 U25 ( .A(in1[33]), .B(in2[33]), .CI(in3[33]), .CO(cout[33]), .S(
        sumout[33]) );
  FADDX1 U26 ( .A(in1[34]), .B(in2[34]), .CI(in3[34]), .CO(cout[34]), .S(
        sumout[34]) );
  FADDX1 U27 ( .A(in1[35]), .B(in2[35]), .CI(in3[35]), .CO(cout[35]), .S(
        sumout[35]) );
  FADDX1 U28 ( .A(in1[36]), .B(in2[36]), .CI(in3[36]), .CO(cout[36]), .S(
        sumout[36]) );
  FADDX1 U29 ( .A(in1[37]), .B(in2[37]), .CI(in3[37]), .CO(cout[37]), .S(
        sumout[37]) );
  FADDX1 U30 ( .A(in1[38]), .B(in2[38]), .CI(in3[38]), .CO(cout[38]), .S(
        sumout[38]) );
  FADDX1 U31 ( .A(in1[39]), .B(in2[39]), .CI(in3[39]), .CO(cout[39]), .S(
        sumout[39]) );
  FADDX1 U32 ( .A(in1[40]), .B(in2[40]), .CI(in3[40]), .CO(cout[40]), .S(
        sumout[40]) );
  FADDX1 U33 ( .A(in1[41]), .B(in2[41]), .CI(in3[41]), .CO(cout[41]), .S(
        sumout[41]) );
  FADDX1 U34 ( .A(in1[42]), .B(in2[42]), .CI(in3[42]), .CO(cout[42]), .S(
        sumout[42]) );
  FADDX1 U35 ( .A(in1[43]), .B(in2[43]), .CI(in3[43]), .CO(cout[43]), .S(
        sumout[43]) );
  FADDX1 U36 ( .A(in1[44]), .B(in2[44]), .CI(in3[44]), .CO(cout[44]), .S(
        sumout[44]) );
  FADDX1 U37 ( .A(in1[45]), .B(in2[45]), .CI(in3[45]), .CO(cout[45]), .S(
        sumout[45]) );
  FADDX1 U38 ( .A(in1[46]), .B(in2[46]), .CI(in3[46]), .CO(cout[46]), .S(
        sumout[46]) );
  XOR3X1 U39 ( .IN1(in2[47]), .IN2(in3[47]), .IN3(in1[47]), .Q(sumout[47]) );
  FADDX1 U40 ( .A(in1[7]), .B(in2[7]), .CI(in3[7]), .CO(cout[7]), .S(sumout[7]) );
  FADDX1 U41 ( .A(in1[8]), .B(in2[8]), .CI(in3[8]), .CO(cout[8]), .S(sumout[8]) );
  FADDX1 U42 ( .A(in1[9]), .B(in2[9]), .CI(in3[9]), .CO(cout[9]), .S(sumout[9]) );
endmodule


module csa51squ_3 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14;

  AND2X1 U1 ( .IN1(in2[7]), .IN2(in1[7]), .Q(cout[7]) );
  NOR2X0 U2 ( .IN1(in2[7]), .IN2(in1[7]), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(cout[7]), .QN(sumout[7]) );
  AND2X1 U4 ( .IN1(in2[8]), .IN2(in1[8]), .Q(cout[8]) );
  NOR2X0 U5 ( .IN1(in2[8]), .IN2(in1[8]), .QN(n2) );
  NOR2X0 U6 ( .IN1(n2), .IN2(cout[8]), .QN(sumout[8]) );
  AND2X1 U7 ( .IN1(in2[9]), .IN2(in1[9]), .Q(cout[9]) );
  NOR2X0 U8 ( .IN1(in2[9]), .IN2(in1[9]), .QN(n3) );
  NOR2X0 U9 ( .IN1(n3), .IN2(cout[9]), .QN(sumout[9]) );
  AND2X1 U10 ( .IN1(in2[10]), .IN2(in1[10]), .Q(cout[10]) );
  NOR2X0 U11 ( .IN1(in2[10]), .IN2(in1[10]), .QN(n4) );
  NOR2X0 U12 ( .IN1(n4), .IN2(cout[10]), .QN(sumout[10]) );
  AND2X1 U13 ( .IN1(in2[11]), .IN2(in1[11]), .Q(cout[11]) );
  NOR2X0 U14 ( .IN1(in2[11]), .IN2(in1[11]), .QN(n5) );
  NOR2X0 U15 ( .IN1(n5), .IN2(cout[11]), .QN(sumout[11]) );
  AND2X1 U16 ( .IN1(in2[12]), .IN2(in1[12]), .Q(cout[12]) );
  NOR2X0 U17 ( .IN1(in2[12]), .IN2(in1[12]), .QN(n6) );
  NOR2X0 U18 ( .IN1(n6), .IN2(cout[12]), .QN(sumout[12]) );
  AND2X1 U19 ( .IN1(in3[40]), .IN2(in2[40]), .Q(cout[40]) );
  NOR2X0 U20 ( .IN1(in3[40]), .IN2(in2[40]), .QN(n7) );
  NOR2X0 U21 ( .IN1(n7), .IN2(cout[40]), .QN(sumout[40]) );
  AND2X1 U22 ( .IN1(in3[41]), .IN2(in2[41]), .Q(cout[41]) );
  NOR2X0 U23 ( .IN1(in3[41]), .IN2(in2[41]), .QN(n8) );
  NOR2X0 U24 ( .IN1(n8), .IN2(cout[41]), .QN(sumout[41]) );
  AND2X1 U25 ( .IN1(in3[42]), .IN2(in2[42]), .Q(cout[42]) );
  NOR2X0 U26 ( .IN1(in3[42]), .IN2(in2[42]), .QN(n9) );
  NOR2X0 U27 ( .IN1(n9), .IN2(cout[42]), .QN(sumout[42]) );
  AND2X1 U28 ( .IN1(in3[43]), .IN2(in2[43]), .Q(cout[43]) );
  NOR2X0 U29 ( .IN1(in3[43]), .IN2(in2[43]), .QN(n10) );
  NOR2X0 U30 ( .IN1(n10), .IN2(cout[43]), .QN(sumout[43]) );
  AND2X1 U31 ( .IN1(in3[44]), .IN2(in2[44]), .Q(cout[44]) );
  NOR2X0 U32 ( .IN1(in3[44]), .IN2(in2[44]), .QN(n11) );
  NOR2X0 U33 ( .IN1(n11), .IN2(cout[44]), .QN(sumout[44]) );
  AND2X1 U34 ( .IN1(in3[45]), .IN2(in2[45]), .Q(cout[45]) );
  NOR2X0 U35 ( .IN1(in3[45]), .IN2(in2[45]), .QN(n12) );
  NOR2X0 U36 ( .IN1(n12), .IN2(cout[45]), .QN(sumout[45]) );
  AND2X1 U37 ( .IN1(in3[46]), .IN2(in2[46]), .Q(cout[46]) );
  NOR2X0 U38 ( .IN1(in3[46]), .IN2(in2[46]), .QN(n13) );
  NOR2X0 U39 ( .IN1(n13), .IN2(cout[46]), .QN(sumout[46]) );
  INVX0 U40 ( .INP(in3[47]), .ZN(sumout[47]) );
  AND2X1 U41 ( .IN1(in2[5]), .IN2(in1[5]), .Q(cout[5]) );
  AND2X1 U42 ( .IN1(in2[6]), .IN2(in1[6]), .Q(cout[6]) );
  NOR2X0 U43 ( .IN1(in2[6]), .IN2(in1[6]), .QN(n14) );
  NOR2X0 U44 ( .IN1(n14), .IN2(cout[6]), .QN(sumout[6]) );
  FADDX1 U45 ( .A(in1[13]), .B(in2[13]), .CI(in3[13]), .CO(cout[13]), .S(
        sumout[13]) );
  FADDX1 U46 ( .A(in1[14]), .B(in2[14]), .CI(in3[14]), .CO(cout[14]), .S(
        sumout[14]) );
  FADDX1 U47 ( .A(in1[15]), .B(in2[15]), .CI(in3[15]), .CO(cout[15]), .S(
        sumout[15]) );
  FADDX1 U48 ( .A(in1[16]), .B(in2[16]), .CI(in3[16]), .CO(cout[16]), .S(
        sumout[16]) );
  FADDX1 U49 ( .A(in1[17]), .B(in2[17]), .CI(in3[17]), .CO(cout[17]), .S(
        sumout[17]) );
  FADDX1 U50 ( .A(in1[18]), .B(in2[18]), .CI(in3[18]), .CO(cout[18]), .S(
        sumout[18]) );
  FADDX1 U51 ( .A(in1[19]), .B(in2[19]), .CI(in3[19]), .CO(cout[19]), .S(
        sumout[19]) );
  FADDX1 U52 ( .A(in1[20]), .B(in2[20]), .CI(in3[20]), .CO(cout[20]), .S(
        sumout[20]) );
  FADDX1 U53 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U54 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U55 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U56 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U57 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U58 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U59 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U60 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U61 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U62 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U63 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U64 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
  FADDX1 U65 ( .A(in1[33]), .B(in2[33]), .CI(in3[33]), .CO(cout[33]), .S(
        sumout[33]) );
  FADDX1 U66 ( .A(in1[34]), .B(in2[34]), .CI(in3[34]), .CO(cout[34]), .S(
        sumout[34]) );
  FADDX1 U67 ( .A(in1[35]), .B(in2[35]), .CI(in3[35]), .CO(cout[35]), .S(
        sumout[35]) );
  FADDX1 U68 ( .A(in1[36]), .B(in2[36]), .CI(in3[36]), .CO(cout[36]), .S(
        sumout[36]) );
  FADDX1 U69 ( .A(in1[37]), .B(in2[37]), .CI(in3[37]), .CO(cout[37]), .S(
        sumout[37]) );
  FADDX1 U70 ( .A(in1[38]), .B(in2[38]), .CI(in3[38]), .CO(cout[38]), .S(
        sumout[38]) );
  FADDX1 U71 ( .A(in1[39]), .B(in2[39]), .CI(in3[39]), .CO(cout[39]), .S(
        sumout[39]) );
endmodule


module csa51squ_4 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17;

  NBUFFX2 U1 ( .INP(in1[6]), .Z(sumout[6]) );
  NBUFFX2 U2 ( .INP(in1[7]), .Z(sumout[7]) );
  NBUFFX2 U3 ( .INP(in1[8]), .Z(sumout[8]) );
  NBUFFX2 U4 ( .INP(in1[9]), .Z(sumout[9]) );
  NBUFFX2 U5 ( .INP(in1[10]), .Z(sumout[10]) );
  NBUFFX2 U6 ( .INP(in1[11]), .Z(sumout[11]) );
  AND2X1 U7 ( .IN1(in3[13]), .IN2(in1[13]), .Q(cout[13]) );
  NOR2X0 U8 ( .IN1(in3[13]), .IN2(in1[13]), .QN(n7) );
  NOR2X0 U9 ( .IN1(n7), .IN2(cout[13]), .QN(sumout[13]) );
  AND2X1 U10 ( .IN1(in3[15]), .IN2(in1[15]), .Q(cout[15]) );
  NOR2X0 U11 ( .IN1(in3[15]), .IN2(in1[15]), .QN(n8) );
  NOR2X0 U12 ( .IN1(n8), .IN2(cout[15]), .QN(sumout[15]) );
  AND2X1 U13 ( .IN1(in3[17]), .IN2(in1[17]), .Q(cout[17]) );
  NOR2X0 U14 ( .IN1(in3[17]), .IN2(in1[17]), .QN(n9) );
  NOR2X0 U15 ( .IN1(n9), .IN2(cout[17]), .QN(sumout[17]) );
  AND2X1 U16 ( .IN1(in3[43]), .IN2(in2[43]), .Q(cout[43]) );
  NOR2X0 U17 ( .IN1(in3[43]), .IN2(in2[43]), .QN(n10) );
  NOR2X0 U18 ( .IN1(n10), .IN2(cout[43]), .QN(sumout[43]) );
  AND2X1 U19 ( .IN1(in3[44]), .IN2(in2[44]), .Q(cout[44]) );
  NOR2X0 U20 ( .IN1(in3[44]), .IN2(in2[44]), .QN(n11) );
  NOR2X0 U21 ( .IN1(n11), .IN2(cout[44]), .QN(sumout[44]) );
  AND2X1 U22 ( .IN1(in3[45]), .IN2(in2[45]), .Q(cout[45]) );
  NOR2X0 U23 ( .IN1(in3[45]), .IN2(in2[45]), .QN(n12) );
  NOR2X0 U24 ( .IN1(n12), .IN2(cout[45]), .QN(sumout[45]) );
  AND2X1 U25 ( .IN1(in3[46]), .IN2(in2[46]), .Q(cout[46]) );
  NOR2X0 U26 ( .IN1(in3[46]), .IN2(in2[46]), .QN(n13) );
  NOR2X0 U27 ( .IN1(n13), .IN2(cout[46]), .QN(sumout[46]) );
  XOR2X1 U28 ( .IN1(in3[47]), .IN2(in2[47]), .Q(sumout[47]) );
  AND2X1 U29 ( .IN1(in3[12]), .IN2(in1[12]), .Q(cout[12]) );
  NOR2X0 U30 ( .IN1(in3[12]), .IN2(in1[12]), .QN(n14) );
  NOR2X0 U31 ( .IN1(n14), .IN2(cout[12]), .QN(sumout[12]) );
  AND2X1 U32 ( .IN1(in3[14]), .IN2(in1[14]), .Q(cout[14]) );
  NOR2X0 U33 ( .IN1(in3[14]), .IN2(in1[14]), .QN(n15) );
  NOR2X0 U34 ( .IN1(n15), .IN2(cout[14]), .QN(sumout[14]) );
  AND2X1 U35 ( .IN1(in3[16]), .IN2(in1[16]), .Q(cout[16]) );
  NOR2X0 U36 ( .IN1(in3[16]), .IN2(in1[16]), .QN(n16) );
  NOR2X0 U37 ( .IN1(n16), .IN2(cout[16]), .QN(sumout[16]) );
  AND2X1 U38 ( .IN1(in3[18]), .IN2(in1[18]), .Q(cout[18]) );
  NOR2X0 U39 ( .IN1(in3[18]), .IN2(in1[18]), .QN(n17) );
  NOR2X0 U40 ( .IN1(n17), .IN2(cout[18]), .QN(sumout[18]) );
  FADDX1 U41 ( .A(in1[19]), .B(in2[19]), .CI(in3[19]), .CO(cout[19]), .S(
        sumout[19]) );
  FADDX1 U42 ( .A(in1[20]), .B(in2[20]), .CI(in3[20]), .CO(cout[20]), .S(
        sumout[20]) );
  FADDX1 U43 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U44 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U45 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U46 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U47 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U48 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U49 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U50 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U51 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U52 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U53 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U54 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
  FADDX1 U55 ( .A(in1[33]), .B(in2[33]), .CI(in3[33]), .CO(cout[33]), .S(
        sumout[33]) );
  FADDX1 U56 ( .A(in1[34]), .B(in2[34]), .CI(in3[34]), .CO(cout[34]), .S(
        sumout[34]) );
  FADDX1 U57 ( .A(in1[35]), .B(in2[35]), .CI(in3[35]), .CO(cout[35]), .S(
        sumout[35]) );
  FADDX1 U58 ( .A(in1[36]), .B(in2[36]), .CI(in3[36]), .CO(cout[36]), .S(
        sumout[36]) );
  FADDX1 U59 ( .A(in1[37]), .B(in2[37]), .CI(in3[37]), .CO(cout[37]), .S(
        sumout[37]) );
  FADDX1 U60 ( .A(in1[38]), .B(in2[38]), .CI(in3[38]), .CO(cout[38]), .S(
        sumout[38]) );
  FADDX1 U61 ( .A(in1[39]), .B(in2[39]), .CI(in3[39]), .CO(cout[39]), .S(
        sumout[39]) );
  FADDX1 U62 ( .A(in1[40]), .B(in2[40]), .CI(in3[40]), .CO(cout[40]), .S(
        sumout[40]) );
  FADDX1 U63 ( .A(in1[41]), .B(in2[41]), .CI(in3[41]), .CO(cout[41]), .S(
        sumout[41]) );
  FADDX1 U64 ( .A(in1[42]), .B(in2[42]), .CI(in3[42]), .CO(cout[42]), .S(
        sumout[42]) );
endmodule


module csa51squ_5 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19;

  NBUFFX2 U1 ( .INP(in2[46]), .Z(sumout[46]) );
  NBUFFX2 U2 ( .INP(in2[45]), .Z(sumout[45]) );
  NBUFFX2 U3 ( .INP(in2[44]), .Z(sumout[44]) );
  NBUFFX2 U4 ( .INP(in2[43]), .Z(sumout[43]) );
  NBUFFX2 U5 ( .INP(in2[42]), .Z(sumout[42]) );
  NBUFFX2 U6 ( .INP(in2[41]), .Z(sumout[41]) );
  NBUFFX2 U7 ( .INP(in2[40]), .Z(sumout[40]) );
  NBUFFX2 U8 ( .INP(in2[39]), .Z(sumout[39]) );
  AND2X1 U9 ( .IN1(in2[7]), .IN2(in1[7]), .Q(cout[7]) );
  NOR2X0 U10 ( .IN1(in2[7]), .IN2(in1[7]), .QN(n9) );
  NOR2X0 U11 ( .IN1(n9), .IN2(cout[7]), .QN(sumout[7]) );
  AND2X1 U12 ( .IN1(in2[8]), .IN2(in1[8]), .Q(cout[8]) );
  NOR2X0 U13 ( .IN1(in2[8]), .IN2(in1[8]), .QN(n10) );
  NOR2X0 U14 ( .IN1(n10), .IN2(cout[8]), .QN(sumout[8]) );
  AND2X1 U15 ( .IN1(in2[9]), .IN2(in1[9]), .Q(cout[9]) );
  NOR2X0 U16 ( .IN1(in2[9]), .IN2(in1[9]), .QN(n11) );
  NOR2X0 U17 ( .IN1(n11), .IN2(cout[9]), .QN(sumout[9]) );
  AND2X1 U18 ( .IN1(in3[33]), .IN2(in2[33]), .Q(cout[33]) );
  NOR2X0 U19 ( .IN1(in3[33]), .IN2(in2[33]), .QN(n12) );
  NOR2X0 U20 ( .IN1(n12), .IN2(cout[33]), .QN(sumout[33]) );
  AND2X1 U21 ( .IN1(in3[34]), .IN2(in2[34]), .Q(cout[34]) );
  NOR2X0 U22 ( .IN1(in3[34]), .IN2(in2[34]), .QN(n13) );
  NOR2X0 U23 ( .IN1(n13), .IN2(cout[34]), .QN(sumout[34]) );
  AND2X1 U24 ( .IN1(in3[35]), .IN2(in2[35]), .Q(cout[35]) );
  NOR2X0 U25 ( .IN1(in3[35]), .IN2(in2[35]), .QN(n14) );
  NOR2X0 U26 ( .IN1(n14), .IN2(cout[35]), .QN(sumout[35]) );
  AND2X1 U27 ( .IN1(in3[36]), .IN2(in2[36]), .Q(cout[36]) );
  NOR2X0 U28 ( .IN1(in3[36]), .IN2(in2[36]), .QN(n15) );
  NOR2X0 U29 ( .IN1(n15), .IN2(cout[36]), .QN(sumout[36]) );
  AND2X1 U30 ( .IN1(in3[37]), .IN2(in2[37]), .Q(cout[37]) );
  NOR2X0 U31 ( .IN1(in3[37]), .IN2(in2[37]), .QN(n16) );
  NOR2X0 U32 ( .IN1(n16), .IN2(cout[37]), .QN(sumout[37]) );
  AND2X1 U33 ( .IN1(in3[38]), .IN2(in2[38]), .Q(cout[38]) );
  NOR2X0 U34 ( .IN1(in3[38]), .IN2(in2[38]), .QN(n17) );
  NOR2X0 U35 ( .IN1(n17), .IN2(cout[38]), .QN(sumout[38]) );
  AND2X1 U36 ( .IN1(in2[4]), .IN2(in1[4]), .Q(cout[4]) );
  AND2X1 U37 ( .IN1(in2[5]), .IN2(in1[5]), .Q(cout[5]) );
  NOR2X0 U38 ( .IN1(in2[5]), .IN2(in1[5]), .QN(n18) );
  NOR2X0 U39 ( .IN1(n18), .IN2(cout[5]), .QN(sumout[5]) );
  AND2X1 U40 ( .IN1(in2[6]), .IN2(in1[6]), .Q(cout[6]) );
  NOR2X0 U41 ( .IN1(in2[6]), .IN2(in1[6]), .QN(n19) );
  NOR2X0 U42 ( .IN1(n19), .IN2(cout[6]), .QN(sumout[6]) );
  FADDX1 U43 ( .A(in1[10]), .B(in2[10]), .CI(in3[10]), .CO(cout[10]), .S(
        sumout[10]) );
  FADDX1 U44 ( .A(in1[11]), .B(in2[11]), .CI(in3[11]), .CO(cout[11]), .S(
        sumout[11]) );
  FADDX1 U45 ( .A(in1[12]), .B(in2[12]), .CI(in3[12]), .CO(cout[12]), .S(
        sumout[12]) );
  FADDX1 U46 ( .A(in1[13]), .B(in2[13]), .CI(in3[13]), .CO(cout[13]), .S(
        sumout[13]) );
  FADDX1 U47 ( .A(in1[14]), .B(in2[14]), .CI(in3[14]), .CO(cout[14]), .S(
        sumout[14]) );
  FADDX1 U48 ( .A(in1[15]), .B(in2[15]), .CI(in3[15]), .CO(cout[15]), .S(
        sumout[15]) );
  FADDX1 U49 ( .A(in1[16]), .B(in2[16]), .CI(in3[16]), .CO(cout[16]), .S(
        sumout[16]) );
  FADDX1 U50 ( .A(in1[17]), .B(in2[17]), .CI(in3[17]), .CO(cout[17]), .S(
        sumout[17]) );
  FADDX1 U51 ( .A(in1[18]), .B(in2[18]), .CI(in3[18]), .CO(cout[18]), .S(
        sumout[18]) );
  FADDX1 U52 ( .A(in1[19]), .B(in2[19]), .CI(in3[19]), .CO(cout[19]), .S(
        sumout[19]) );
  FADDX1 U53 ( .A(in1[20]), .B(in2[20]), .CI(in3[20]), .CO(cout[20]), .S(
        sumout[20]) );
  FADDX1 U54 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U55 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U56 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U57 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U58 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U59 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U60 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U61 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U62 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U63 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U64 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U65 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
endmodule


module csa51squ_6 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n7, n8, n9, n10, n11, n12, n13;

  NBUFFX2 U1 ( .INP(in1[12]), .Z(sumout[12]) );
  NBUFFX2 U2 ( .INP(in1[13]), .Z(sumout[13]) );
  NBUFFX2 U3 ( .INP(in1[14]), .Z(sumout[14]) );
  NBUFFX2 U4 ( .INP(in1[15]), .Z(sumout[15]) );
  NBUFFX2 U5 ( .INP(in1[16]), .Z(sumout[16]) );
  NBUFFX2 U6 ( .INP(in1[17]), .Z(sumout[17]) );
  AND2X1 U7 ( .IN1(in3[19]), .IN2(in1[19]), .Q(cout[19]) );
  NOR2X0 U8 ( .IN1(in3[19]), .IN2(in1[19]), .QN(n7) );
  NOR2X0 U9 ( .IN1(n7), .IN2(cout[19]), .QN(sumout[19]) );
  AND2X1 U10 ( .IN1(in3[44]), .IN2(in2[44]), .Q(cout[44]) );
  NOR2X0 U11 ( .IN1(in3[44]), .IN2(in2[44]), .QN(n8) );
  NOR2X0 U12 ( .IN1(n8), .IN2(cout[44]), .QN(sumout[44]) );
  AND2X1 U13 ( .IN1(in3[45]), .IN2(in2[45]), .Q(cout[45]) );
  NOR2X0 U14 ( .IN1(in3[45]), .IN2(in2[45]), .QN(n9) );
  NOR2X0 U15 ( .IN1(n9), .IN2(cout[45]), .QN(sumout[45]) );
  AND2X1 U16 ( .IN1(in3[46]), .IN2(in2[46]), .Q(cout[46]) );
  NOR2X0 U17 ( .IN1(in3[46]), .IN2(in2[46]), .QN(n10) );
  NOR2X0 U18 ( .IN1(n10), .IN2(cout[46]), .QN(sumout[46]) );
  XOR2X1 U19 ( .IN1(in3[47]), .IN2(in2[47]), .Q(sumout[47]) );
  AND2X1 U20 ( .IN1(in3[18]), .IN2(in1[18]), .Q(cout[18]) );
  NOR2X0 U21 ( .IN1(in3[18]), .IN2(in1[18]), .QN(n11) );
  NOR2X0 U22 ( .IN1(n11), .IN2(cout[18]), .QN(sumout[18]) );
  AND2X1 U23 ( .IN1(in3[20]), .IN2(in1[20]), .Q(cout[20]) );
  NOR2X0 U24 ( .IN1(in3[20]), .IN2(in1[20]), .QN(n12) );
  NOR2X0 U25 ( .IN1(n12), .IN2(cout[20]), .QN(sumout[20]) );
  INVX0 U26 ( .INP(in1[42]), .ZN(n13) );
  FADDX1 U27 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U28 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U29 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U30 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U31 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U32 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U33 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U34 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U35 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U36 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U37 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U38 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
  FADDX1 U39 ( .A(in1[33]), .B(in2[33]), .CI(in3[33]), .CO(cout[33]), .S(
        sumout[33]) );
  FADDX1 U40 ( .A(in1[34]), .B(in2[34]), .CI(in3[34]), .CO(cout[34]), .S(
        sumout[34]) );
  FADDX1 U41 ( .A(in1[35]), .B(in2[35]), .CI(in3[35]), .CO(cout[35]), .S(
        sumout[35]) );
  FADDX1 U42 ( .A(in1[36]), .B(in2[36]), .CI(in3[36]), .CO(cout[36]), .S(
        sumout[36]) );
  FADDX1 U43 ( .A(in1[37]), .B(in2[37]), .CI(in3[37]), .CO(cout[37]), .S(
        sumout[37]) );
  FADDX1 U44 ( .A(in1[38]), .B(in2[38]), .CI(in3[38]), .CO(cout[38]), .S(
        sumout[38]) );
  FADDX1 U45 ( .A(in1[39]), .B(in2[39]), .CI(in3[39]), .CO(cout[39]), .S(
        sumout[39]) );
  FADDX1 U46 ( .A(in1[40]), .B(in2[40]), .CI(in3[40]), .CO(cout[40]), .S(
        sumout[40]) );
  FADDX1 U47 ( .A(in1[41]), .B(in2[41]), .CI(in3[41]), .CO(cout[41]), .S(
        sumout[41]) );
  FADDX1 U48 ( .A(in1[42]), .B(in2[42]), .CI(in3[42]), .CO(cout[42]), .S(
        sumout[42]) );
  FADDX1 U49 ( .A(in2[43]), .B(in3[43]), .CI(n13), .CO(cout[43]), .S(
        sumout[43]) );
endmodule


module csa51squ_7 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n9, n10, n11, n12, n13, n14, n15;

  NBUFFX2 U1 ( .INP(in2[6]), .Z(sumout[6]) );
  NBUFFX2 U2 ( .INP(in2[7]), .Z(sumout[7]) );
  NBUFFX2 U3 ( .INP(in2[8]), .Z(sumout[8]) );
  NBUFFX2 U4 ( .INP(in3[42]), .Z(sumout[42]) );
  NBUFFX2 U5 ( .INP(in3[41]), .Z(sumout[41]) );
  NBUFFX2 U6 ( .INP(in3[39]), .Z(sumout[39]) );
  NBUFFX2 U7 ( .INP(in3[38]), .Z(sumout[38]) );
  NBUFFX2 U8 ( .INP(in3[40]), .Z(sumout[40]) );
  AND2X1 U9 ( .IN1(in2[13]), .IN2(in1[13]), .Q(cout[13]) );
  NOR2X0 U10 ( .IN1(in2[13]), .IN2(in1[13]), .QN(n9) );
  NOR2X0 U11 ( .IN1(n9), .IN2(cout[13]), .QN(sumout[13]) );
  AND2X1 U12 ( .IN1(in2[37]), .IN2(in3[37]), .Q(cout[37]) );
  INVX0 U13 ( .INP(in2[37]), .ZN(n15) );
  MUX21X1 U14 ( .IN1(in2[37]), .IN2(n15), .S(in3[37]), .Q(sumout[37]) );
  AND2X1 U15 ( .IN1(in2[9]), .IN2(in1[9]), .Q(cout[9]) );
  NOR2X0 U16 ( .IN1(in2[9]), .IN2(in1[9]), .QN(n10) );
  NOR2X0 U17 ( .IN1(n10), .IN2(cout[9]), .QN(sumout[9]) );
  AND2X1 U18 ( .IN1(in2[10]), .IN2(in1[10]), .Q(cout[10]) );
  NOR2X0 U19 ( .IN1(in2[10]), .IN2(in1[10]), .QN(n11) );
  NOR2X0 U20 ( .IN1(n11), .IN2(cout[10]), .QN(sumout[10]) );
  AND2X1 U21 ( .IN1(in2[11]), .IN2(in1[11]), .Q(cout[11]) );
  NOR2X0 U22 ( .IN1(in2[11]), .IN2(in1[11]), .QN(n12) );
  NOR2X0 U23 ( .IN1(n12), .IN2(cout[11]), .QN(sumout[11]) );
  AND2X1 U24 ( .IN1(in2[12]), .IN2(in1[12]), .Q(cout[12]) );
  NOR2X0 U25 ( .IN1(in2[12]), .IN2(in1[12]), .QN(n13) );
  NOR2X0 U26 ( .IN1(n13), .IN2(cout[12]), .QN(sumout[12]) );
  AND2X1 U27 ( .IN1(in2[14]), .IN2(in1[14]), .Q(cout[14]) );
  NOR2X0 U28 ( .IN1(in2[14]), .IN2(in1[14]), .QN(n14) );
  NOR2X0 U29 ( .IN1(n14), .IN2(cout[14]), .QN(sumout[14]) );
  FADDX1 U30 ( .A(in1[15]), .B(in2[15]), .CI(in3[15]), .CO(cout[15]), .S(
        sumout[15]) );
  FADDX1 U31 ( .A(in1[16]), .B(in2[16]), .CI(in3[16]), .CO(cout[16]), .S(
        sumout[16]) );
  FADDX1 U32 ( .A(in1[17]), .B(in2[17]), .CI(in3[17]), .CO(cout[17]), .S(
        sumout[17]) );
  FADDX1 U33 ( .A(in1[18]), .B(in2[18]), .CI(in3[18]), .CO(cout[18]), .S(
        sumout[18]) );
  FADDX1 U34 ( .A(in1[19]), .B(in2[19]), .CI(in3[19]), .CO(cout[19]), .S(
        sumout[19]) );
  FADDX1 U35 ( .A(in1[20]), .B(in2[20]), .CI(in3[20]), .CO(cout[20]), .S(
        sumout[20]) );
  FADDX1 U36 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U37 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U38 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U39 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U40 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U41 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U42 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U43 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U44 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U45 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U46 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U47 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
  FADDX1 U48 ( .A(in1[33]), .B(in2[33]), .CI(in3[33]), .CO(cout[33]), .S(
        sumout[33]) );
  FADDX1 U49 ( .A(in1[34]), .B(in2[34]), .CI(in3[34]), .CO(cout[34]), .S(
        sumout[34]) );
  FADDX1 U50 ( .A(in1[35]), .B(in2[35]), .CI(in3[35]), .CO(cout[35]), .S(
        sumout[35]) );
  FADDX1 U51 ( .A(in1[36]), .B(in3[36]), .CI(n15), .CO(cout[36]), .S(
        sumout[36]) );
endmodule


module csa51squ_8 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36;

  NBUFFX2 U1 ( .INP(in3[46]), .Z(sumout[46]) );
  NBUFFX2 U2 ( .INP(in3[45]), .Z(sumout[45]) );
  NBUFFX2 U3 ( .INP(in3[44]), .Z(sumout[44]) );
  NBUFFX2 U4 ( .INP(in3[43]), .Z(sumout[43]) );
  NBUFFX2 U5 ( .INP(in3[42]), .Z(sumout[42]) );
  NBUFFX2 U6 ( .INP(in3[33]), .Z(sumout[33]) );
  NBUFFX2 U7 ( .INP(in3[32]), .Z(sumout[32]) );
  NBUFFX2 U8 ( .INP(in3[35]), .Z(sumout[35]) );
  NBUFFX2 U9 ( .INP(in3[34]), .Z(sumout[34]) );
  NBUFFX2 U10 ( .INP(in3[37]), .Z(sumout[37]) );
  NBUFFX2 U11 ( .INP(in3[36]), .Z(sumout[36]) );
  NBUFFX2 U12 ( .INP(in3[41]), .Z(sumout[41]) );
  NBUFFX2 U13 ( .INP(in3[40]), .Z(sumout[40]) );
  NBUFFX2 U14 ( .INP(in3[39]), .Z(sumout[39]) );
  NBUFFX2 U15 ( .INP(in3[38]), .Z(sumout[38]) );
  AND2X1 U16 ( .IN1(in2[31]), .IN2(in3[31]), .Q(cout[31]) );
  INVX0 U17 ( .INP(in2[31]), .ZN(n36) );
  MUX21X1 U18 ( .IN1(in2[31]), .IN2(n36), .S(in3[31]), .Q(sumout[31]) );
  AND2X1 U19 ( .IN1(in2[3]), .IN2(in1[3]), .Q(cout[3]) );
  AND2X1 U20 ( .IN1(in2[4]), .IN2(in1[4]), .Q(cout[4]) );
  NOR2X0 U21 ( .IN1(in2[4]), .IN2(in1[4]), .QN(n16) );
  NOR2X0 U22 ( .IN1(n16), .IN2(cout[4]), .QN(sumout[4]) );
  AND2X1 U23 ( .IN1(in2[5]), .IN2(in1[5]), .Q(cout[5]) );
  NOR2X0 U24 ( .IN1(in2[5]), .IN2(in1[5]), .QN(n17) );
  NOR2X0 U25 ( .IN1(n17), .IN2(cout[5]), .QN(sumout[5]) );
  AND2X1 U26 ( .IN1(in2[6]), .IN2(in1[6]), .Q(cout[6]) );
  NOR2X0 U27 ( .IN1(in2[6]), .IN2(in1[6]), .QN(n18) );
  NOR2X0 U28 ( .IN1(n18), .IN2(cout[6]), .QN(sumout[6]) );
  AND2X1 U29 ( .IN1(in2[7]), .IN2(in1[7]), .Q(cout[7]) );
  NOR2X0 U30 ( .IN1(in2[7]), .IN2(in1[7]), .QN(n19) );
  NOR2X0 U31 ( .IN1(n19), .IN2(cout[7]), .QN(sumout[7]) );
  AND2X1 U32 ( .IN1(in2[8]), .IN2(in1[8]), .Q(cout[8]) );
  NOR2X0 U33 ( .IN1(in2[8]), .IN2(in1[8]), .QN(n20) );
  NOR2X0 U34 ( .IN1(n20), .IN2(cout[8]), .QN(sumout[8]) );
  AND2X1 U35 ( .IN1(in2[9]), .IN2(in1[9]), .Q(cout[9]) );
  NOR2X0 U36 ( .IN1(in2[9]), .IN2(in1[9]), .QN(n21) );
  NOR2X0 U37 ( .IN1(n21), .IN2(cout[9]), .QN(sumout[9]) );
  AND2X1 U38 ( .IN1(in2[10]), .IN2(in1[10]), .Q(cout[10]) );
  NOR2X0 U39 ( .IN1(in2[10]), .IN2(in1[10]), .QN(n22) );
  NOR2X0 U40 ( .IN1(n22), .IN2(cout[10]), .QN(sumout[10]) );
  AND2X1 U41 ( .IN1(in2[11]), .IN2(in1[11]), .Q(cout[11]) );
  NOR2X0 U42 ( .IN1(in2[11]), .IN2(in1[11]), .QN(n23) );
  NOR2X0 U43 ( .IN1(n23), .IN2(cout[11]), .QN(sumout[11]) );
  AND2X1 U44 ( .IN1(in2[12]), .IN2(in1[12]), .Q(cout[12]) );
  NOR2X0 U45 ( .IN1(in2[12]), .IN2(in1[12]), .QN(n24) );
  NOR2X0 U46 ( .IN1(n24), .IN2(cout[12]), .QN(sumout[12]) );
  AND2X1 U47 ( .IN1(in2[13]), .IN2(in1[13]), .Q(cout[13]) );
  NOR2X0 U48 ( .IN1(in2[13]), .IN2(in1[13]), .QN(n25) );
  NOR2X0 U49 ( .IN1(n25), .IN2(cout[13]), .QN(sumout[13]) );
  AND2X1 U50 ( .IN1(in2[14]), .IN2(in1[14]), .Q(cout[14]) );
  NOR2X0 U51 ( .IN1(in2[14]), .IN2(in1[14]), .QN(n26) );
  NOR2X0 U52 ( .IN1(n26), .IN2(cout[14]), .QN(sumout[14]) );
  AND2X1 U53 ( .IN1(in2[15]), .IN2(in1[15]), .Q(cout[15]) );
  NOR2X0 U54 ( .IN1(in2[15]), .IN2(in1[15]), .QN(n27) );
  NOR2X0 U55 ( .IN1(n27), .IN2(cout[15]), .QN(sumout[15]) );
  AND2X1 U56 ( .IN1(in2[16]), .IN2(in1[16]), .Q(cout[16]) );
  NOR2X0 U57 ( .IN1(in2[16]), .IN2(in1[16]), .QN(n28) );
  NOR2X0 U58 ( .IN1(n28), .IN2(cout[16]), .QN(sumout[16]) );
  AND2X1 U59 ( .IN1(in2[17]), .IN2(in1[17]), .Q(cout[17]) );
  NOR2X0 U60 ( .IN1(in2[17]), .IN2(in1[17]), .QN(n29) );
  NOR2X0 U61 ( .IN1(n29), .IN2(cout[17]), .QN(sumout[17]) );
  AND2X1 U62 ( .IN1(in2[18]), .IN2(in1[18]), .Q(cout[18]) );
  NOR2X0 U63 ( .IN1(in2[18]), .IN2(in1[18]), .QN(n30) );
  NOR2X0 U64 ( .IN1(n30), .IN2(cout[18]), .QN(sumout[18]) );
  AND2X1 U65 ( .IN1(in2[19]), .IN2(in1[19]), .Q(cout[19]) );
  NOR2X0 U66 ( .IN1(in2[19]), .IN2(in1[19]), .QN(n31) );
  NOR2X0 U67 ( .IN1(n31), .IN2(cout[19]), .QN(sumout[19]) );
  AND2X1 U68 ( .IN1(in2[20]), .IN2(in1[20]), .Q(cout[20]) );
  NOR2X0 U69 ( .IN1(in2[20]), .IN2(in1[20]), .QN(n32) );
  NOR2X0 U70 ( .IN1(n32), .IN2(cout[20]), .QN(sumout[20]) );
  AND2X1 U71 ( .IN1(in2[21]), .IN2(in1[21]), .Q(cout[21]) );
  NOR2X0 U72 ( .IN1(in2[21]), .IN2(in1[21]), .QN(n33) );
  NOR2X0 U73 ( .IN1(n33), .IN2(cout[21]), .QN(sumout[21]) );
  AND2X1 U74 ( .IN1(in2[22]), .IN2(in1[22]), .Q(cout[22]) );
  NOR2X0 U75 ( .IN1(in2[22]), .IN2(in1[22]), .QN(n34) );
  NOR2X0 U76 ( .IN1(n34), .IN2(cout[22]), .QN(sumout[22]) );
  AND2X1 U77 ( .IN1(in2[23]), .IN2(in1[23]), .Q(cout[23]) );
  NOR2X0 U78 ( .IN1(in2[23]), .IN2(in1[23]), .QN(n35) );
  NOR2X0 U79 ( .IN1(n35), .IN2(cout[23]), .QN(sumout[23]) );
  FADDX1 U80 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U81 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U82 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U83 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U84 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U85 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U86 ( .A(in1[30]), .B(in3[30]), .CI(n36), .CO(cout[30]), .S(
        sumout[30]) );
endmodule


module csa51squ_9 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n3, n4, n5, n6, n7;

  NBUFFX2 U1 ( .INP(in1[18]), .Z(sumout[18]) );
  NBUFFX2 U2 ( .INP(in1[19]), .Z(sumout[19]) );
  AND2X1 U3 ( .IN1(in2[20]), .IN2(in1[20]), .Q(cout[20]) );
  NOR2X0 U4 ( .IN1(in2[20]), .IN2(in1[20]), .QN(n3) );
  NOR2X0 U5 ( .IN1(n3), .IN2(cout[20]), .QN(sumout[20]) );
  AND2X1 U6 ( .IN1(in2[21]), .IN2(in1[21]), .Q(cout[21]) );
  NOR2X0 U7 ( .IN1(in2[21]), .IN2(in1[21]), .QN(n4) );
  NOR2X0 U8 ( .IN1(n4), .IN2(cout[21]), .QN(sumout[21]) );
  AND2X1 U9 ( .IN1(in2[46]), .IN2(in3[46]), .Q(cout[46]) );
  NOR2X0 U10 ( .IN1(in2[46]), .IN2(in3[46]), .QN(n5) );
  NOR2X0 U11 ( .IN1(n5), .IN2(cout[46]), .QN(sumout[46]) );
  INVX0 U12 ( .INP(in2[46]), .ZN(n6) );
  MUX21X1 U13 ( .IN1(n6), .IN2(in2[46]), .S(in3[47]), .Q(sumout[47]) );
  INVX0 U14 ( .INP(in1[44]), .ZN(n7) );
  FADDX1 U15 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U16 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U17 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U18 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U19 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U20 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U21 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U22 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U23 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U24 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U25 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
  FADDX1 U26 ( .A(in1[33]), .B(in2[33]), .CI(in3[33]), .CO(cout[33]), .S(
        sumout[33]) );
  FADDX1 U27 ( .A(in1[34]), .B(in2[34]), .CI(in3[34]), .CO(cout[34]), .S(
        sumout[34]) );
  FADDX1 U28 ( .A(in1[35]), .B(in2[35]), .CI(in3[35]), .CO(cout[35]), .S(
        sumout[35]) );
  FADDX1 U29 ( .A(in1[36]), .B(in2[36]), .CI(in3[36]), .CO(cout[36]), .S(
        sumout[36]) );
  FADDX1 U30 ( .A(in1[37]), .B(in2[37]), .CI(in3[37]), .CO(cout[37]), .S(
        sumout[37]) );
  FADDX1 U31 ( .A(in1[38]), .B(in2[38]), .CI(in3[38]), .CO(cout[38]), .S(
        sumout[38]) );
  FADDX1 U32 ( .A(in1[39]), .B(in2[39]), .CI(in3[39]), .CO(cout[39]), .S(
        sumout[39]) );
  FADDX1 U33 ( .A(in1[40]), .B(in2[40]), .CI(in3[40]), .CO(cout[40]), .S(
        sumout[40]) );
  FADDX1 U34 ( .A(in1[41]), .B(in2[41]), .CI(in3[41]), .CO(cout[41]), .S(
        sumout[41]) );
  FADDX1 U35 ( .A(in1[42]), .B(in2[42]), .CI(in3[42]), .CO(cout[42]), .S(
        sumout[42]) );
  FADDX1 U36 ( .A(in1[43]), .B(in2[43]), .CI(in3[43]), .CO(cout[43]), .S(
        sumout[43]) );
  FADDX1 U37 ( .A(in1[44]), .B(in2[44]), .CI(in3[44]), .CO(cout[44]), .S(
        sumout[44]) );
  FADDX1 U38 ( .A(in2[45]), .B(in3[45]), .CI(n7), .CO(cout[45]), .S(sumout[45]) );
endmodule


module csa51squ_10 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n4, n5, n6, n7, n8;

  NBUFFX2 U1 ( .INP(in1[12]), .Z(sumout[12]) );
  NBUFFX2 U2 ( .INP(in1[13]), .Z(sumout[13]) );
  NBUFFX2 U3 ( .INP(in3[42]), .Z(sumout[42]) );
  AND2X1 U4 ( .IN1(in2[14]), .IN2(in1[14]), .Q(cout[14]) );
  NOR2X0 U5 ( .IN1(in2[14]), .IN2(in1[14]), .QN(n4) );
  NOR2X0 U6 ( .IN1(n4), .IN2(cout[14]), .QN(sumout[14]) );
  AND2X1 U7 ( .IN1(in2[15]), .IN2(in1[15]), .Q(cout[15]) );
  NOR2X0 U8 ( .IN1(in2[15]), .IN2(in1[15]), .QN(n5) );
  NOR2X0 U9 ( .IN1(n5), .IN2(cout[15]), .QN(sumout[15]) );
  AND2X1 U10 ( .IN1(in2[40]), .IN2(in3[40]), .Q(cout[40]) );
  NOR2X0 U11 ( .IN1(in2[40]), .IN2(in3[40]), .QN(n6) );
  NOR2X0 U12 ( .IN1(n6), .IN2(cout[40]), .QN(sumout[40]) );
  INVX0 U13 ( .INP(in3[41]), .ZN(n7) );
  NOR2X0 U14 ( .IN1(in2[40]), .IN2(n7), .QN(cout[41]) );
  MUX21X1 U15 ( .IN1(n7), .IN2(in3[41]), .S(in2[40]), .Q(sumout[41]) );
  INVX0 U16 ( .INP(in1[38]), .ZN(n8) );
  FADDX1 U17 ( .A(in1[16]), .B(in2[16]), .CI(in3[16]), .CO(cout[16]), .S(
        sumout[16]) );
  FADDX1 U18 ( .A(in1[17]), .B(in2[17]), .CI(in3[17]), .CO(cout[17]), .S(
        sumout[17]) );
  FADDX1 U19 ( .A(in1[18]), .B(in2[18]), .CI(in3[18]), .CO(cout[18]), .S(
        sumout[18]) );
  FADDX1 U20 ( .A(in1[19]), .B(in2[19]), .CI(in3[19]), .CO(cout[19]), .S(
        sumout[19]) );
  FADDX1 U21 ( .A(in1[20]), .B(in2[20]), .CI(in3[20]), .CO(cout[20]), .S(
        sumout[20]) );
  FADDX1 U22 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U23 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U24 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U25 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U26 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U27 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U28 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U29 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U30 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U31 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U32 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U33 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
  FADDX1 U34 ( .A(in1[33]), .B(in2[33]), .CI(in3[33]), .CO(cout[33]), .S(
        sumout[33]) );
  FADDX1 U35 ( .A(in1[34]), .B(in2[34]), .CI(in3[34]), .CO(cout[34]), .S(
        sumout[34]) );
  FADDX1 U36 ( .A(in1[35]), .B(in2[35]), .CI(in3[35]), .CO(cout[35]), .S(
        sumout[35]) );
  FADDX1 U37 ( .A(in1[36]), .B(in2[36]), .CI(in3[36]), .CO(cout[36]), .S(
        sumout[36]) );
  FADDX1 U38 ( .A(in1[37]), .B(in2[37]), .CI(in3[37]), .CO(cout[37]), .S(
        sumout[37]) );
  FADDX1 U39 ( .A(in1[38]), .B(in2[38]), .CI(in3[38]), .CO(cout[38]), .S(
        sumout[38]) );
  FADDX1 U40 ( .A(in2[39]), .B(in3[39]), .CI(n8), .CO(cout[39]), .S(sumout[39]) );
endmodule


module csa51squ_11 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n4, n5, n6, n7, n8;

  NBUFFX2 U1 ( .INP(in1[6]), .Z(sumout[6]) );
  NBUFFX2 U2 ( .INP(in1[7]), .Z(sumout[7]) );
  NBUFFX2 U3 ( .INP(in3[37]), .Z(sumout[37]) );
  AND2X1 U4 ( .IN1(in2[8]), .IN2(in1[8]), .Q(cout[8]) );
  NOR2X0 U5 ( .IN1(in2[8]), .IN2(in1[8]), .QN(n4) );
  NOR2X0 U6 ( .IN1(n4), .IN2(cout[8]), .QN(sumout[8]) );
  AND2X1 U7 ( .IN1(in2[9]), .IN2(in1[9]), .Q(cout[9]) );
  NOR2X0 U8 ( .IN1(in2[9]), .IN2(in1[9]), .QN(n5) );
  NOR2X0 U9 ( .IN1(n5), .IN2(cout[9]), .QN(sumout[9]) );
  AND2X1 U10 ( .IN1(in2[34]), .IN2(in3[34]), .Q(cout[34]) );
  NOR2X0 U11 ( .IN1(in2[34]), .IN2(in3[34]), .QN(n6) );
  NOR2X0 U12 ( .IN1(n6), .IN2(cout[34]), .QN(sumout[34]) );
  INVX0 U13 ( .INP(in3[35]), .ZN(n7) );
  NOR2X0 U14 ( .IN1(in2[34]), .IN2(n7), .QN(cout[35]) );
  MUX21X1 U15 ( .IN1(n7), .IN2(in3[35]), .S(in2[34]), .Q(sumout[35]) );
  INVX0 U16 ( .INP(in1[32]), .ZN(n8) );
  FADDX1 U17 ( .A(in1[10]), .B(in2[10]), .CI(in3[10]), .CO(cout[10]), .S(
        sumout[10]) );
  FADDX1 U18 ( .A(in1[11]), .B(in2[11]), .CI(in3[11]), .CO(cout[11]), .S(
        sumout[11]) );
  FADDX1 U19 ( .A(in1[12]), .B(in2[12]), .CI(in3[12]), .CO(cout[12]), .S(
        sumout[12]) );
  FADDX1 U20 ( .A(in1[13]), .B(in2[13]), .CI(in3[13]), .CO(cout[13]), .S(
        sumout[13]) );
  FADDX1 U21 ( .A(in1[14]), .B(in2[14]), .CI(in3[14]), .CO(cout[14]), .S(
        sumout[14]) );
  FADDX1 U22 ( .A(in1[15]), .B(in2[15]), .CI(in3[15]), .CO(cout[15]), .S(
        sumout[15]) );
  FADDX1 U23 ( .A(in1[16]), .B(in2[16]), .CI(in3[16]), .CO(cout[16]), .S(
        sumout[16]) );
  FADDX1 U24 ( .A(in1[17]), .B(in2[17]), .CI(in3[17]), .CO(cout[17]), .S(
        sumout[17]) );
  FADDX1 U25 ( .A(in1[18]), .B(in2[18]), .CI(in3[18]), .CO(cout[18]), .S(
        sumout[18]) );
  FADDX1 U26 ( .A(in1[19]), .B(in2[19]), .CI(in3[19]), .CO(cout[19]), .S(
        sumout[19]) );
  FADDX1 U27 ( .A(in1[20]), .B(in2[20]), .CI(in3[20]), .CO(cout[20]), .S(
        sumout[20]) );
  FADDX1 U28 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U29 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U30 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U31 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U32 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U33 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U34 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U35 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U36 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U37 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U38 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U39 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
  FADDX1 U40 ( .A(in2[33]), .B(in3[33]), .CI(n8), .CO(cout[33]), .S(sumout[33]) );
endmodule


module csa51squ_12 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n2, n3, n4, n5;

  NBUFFX2 U1 ( .INP(in3[31]), .Z(sumout[31]) );
  AND2X1 U2 ( .IN1(in2[2]), .IN2(in1[2]), .Q(cout[2]) );
  AND2X1 U3 ( .IN1(in2[3]), .IN2(in1[3]), .Q(cout[3]) );
  NOR2X0 U4 ( .IN1(in2[3]), .IN2(in1[3]), .QN(n2) );
  NOR2X0 U5 ( .IN1(n2), .IN2(cout[3]), .QN(sumout[3]) );
  AND2X1 U6 ( .IN1(in2[28]), .IN2(in3[28]), .Q(cout[28]) );
  NOR2X0 U7 ( .IN1(in2[28]), .IN2(in3[28]), .QN(n3) );
  NOR2X0 U8 ( .IN1(n3), .IN2(cout[28]), .QN(sumout[28]) );
  INVX0 U9 ( .INP(in3[29]), .ZN(n4) );
  NOR2X0 U10 ( .IN1(in2[28]), .IN2(n4), .QN(cout[29]) );
  MUX21X1 U11 ( .IN1(n4), .IN2(in3[29]), .S(in2[28]), .Q(sumout[29]) );
  INVX0 U12 ( .INP(in1[26]), .ZN(n5) );
  FADDX1 U13 ( .A(in1[10]), .B(in2[10]), .CI(in3[10]), .CO(cout[10]), .S(
        sumout[10]) );
  FADDX1 U14 ( .A(in1[11]), .B(in2[11]), .CI(in3[11]), .CO(cout[11]), .S(
        sumout[11]) );
  FADDX1 U15 ( .A(in1[12]), .B(in2[12]), .CI(in3[12]), .CO(cout[12]), .S(
        sumout[12]) );
  FADDX1 U16 ( .A(in1[13]), .B(in2[13]), .CI(in3[13]), .CO(cout[13]), .S(
        sumout[13]) );
  FADDX1 U17 ( .A(in1[14]), .B(in2[14]), .CI(in3[14]), .CO(cout[14]), .S(
        sumout[14]) );
  FADDX1 U18 ( .A(in1[15]), .B(in2[15]), .CI(in3[15]), .CO(cout[15]), .S(
        sumout[15]) );
  FADDX1 U19 ( .A(in1[16]), .B(in2[16]), .CI(in3[16]), .CO(cout[16]), .S(
        sumout[16]) );
  FADDX1 U20 ( .A(in1[17]), .B(in2[17]), .CI(in3[17]), .CO(cout[17]), .S(
        sumout[17]) );
  FADDX1 U21 ( .A(in1[18]), .B(in2[18]), .CI(in3[18]), .CO(cout[18]), .S(
        sumout[18]) );
  FADDX1 U22 ( .A(in1[19]), .B(in2[19]), .CI(in3[19]), .CO(cout[19]), .S(
        sumout[19]) );
  FADDX1 U23 ( .A(in1[20]), .B(in2[20]), .CI(in3[20]), .CO(cout[20]), .S(
        sumout[20]) );
  FADDX1 U24 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U25 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U26 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U27 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U28 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U29 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U30 ( .A(in2[27]), .B(in3[27]), .CI(n5), .CO(cout[27]), .S(sumout[27]) );
  FADDX1 U31 ( .A(in1[4]), .B(in2[4]), .CI(in3[4]), .CO(cout[4]), .S(sumout[4]) );
  FADDX1 U32 ( .A(in1[5]), .B(in2[5]), .CI(in3[5]), .CO(cout[5]), .S(sumout[5]) );
  FADDX1 U33 ( .A(in1[6]), .B(in2[6]), .CI(in3[6]), .CO(cout[6]), .S(sumout[6]) );
  FADDX1 U34 ( .A(in1[7]), .B(in2[7]), .CI(in3[7]), .CO(cout[7]), .S(sumout[7]) );
  FADDX1 U35 ( .A(in1[8]), .B(in2[8]), .CI(in3[8]), .CO(cout[8]), .S(sumout[8]) );
  FADDX1 U36 ( .A(in1[9]), .B(in2[9]), .CI(in3[9]), .CO(cout[9]), .S(sumout[9]) );
endmodule


module booth27_1 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;


  NBUFFX2 U3 ( .INP(in2[22]), .Z(out1[22]) );
  NBUFFX2 U4 ( .INP(in2[21]), .Z(out1[21]) );
  NBUFFX2 U5 ( .INP(in2[20]), .Z(out1[20]) );
  NBUFFX2 U6 ( .INP(in2[0]), .Z(out1[0]) );
  NBUFFX2 U7 ( .INP(in2[2]), .Z(out1[2]) );
  NBUFFX2 U8 ( .INP(in2[1]), .Z(out1[1]) );
  NBUFFX2 U9 ( .INP(in2[19]), .Z(out1[19]) );
  NBUFFX2 U10 ( .INP(in2[18]), .Z(out1[18]) );
  NBUFFX2 U11 ( .INP(in2[6]), .Z(out1[6]) );
  NBUFFX2 U12 ( .INP(in2[5]), .Z(out1[5]) );
  NBUFFX2 U13 ( .INP(in2[4]), .Z(out1[4]) );
  NBUFFX2 U14 ( .INP(in2[3]), .Z(out1[3]) );
  NBUFFX2 U15 ( .INP(in2[9]), .Z(out1[9]) );
  NBUFFX2 U16 ( .INP(in2[8]), .Z(out1[8]) );
  NBUFFX2 U17 ( .INP(in2[7]), .Z(out1[7]) );
  NBUFFX2 U18 ( .INP(in2[11]), .Z(out1[11]) );
  NBUFFX2 U19 ( .INP(in2[10]), .Z(out1[10]) );
  NBUFFX2 U20 ( .INP(in2[13]), .Z(out1[13]) );
  NBUFFX2 U21 ( .INP(in2[12]), .Z(out1[12]) );
  NBUFFX2 U22 ( .INP(in2[17]), .Z(out1[17]) );
  NBUFFX2 U23 ( .INP(in2[16]), .Z(out1[16]) );
  NBUFFX2 U24 ( .INP(in2[15]), .Z(out1[15]) );
  NBUFFX2 U25 ( .INP(in2[14]), .Z(out1[14]) );
endmodule


module booth27_2 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76;

  NAND2X0 U3 ( .IN1(n1), .IN2(n2), .QN(n8) );
  NAND2X0 U4 ( .IN1(n71), .IN2(in2[0]), .QN(n15) );
  NAND2X0 U5 ( .IN1(n16), .IN2(in2[4]), .QN(n17) );
  NAND2X0 U6 ( .IN1(n19), .IN2(in2[5]), .QN(n20) );
  NAND2X0 U7 ( .IN1(n25), .IN2(in2[7]), .QN(n26) );
  NAND2X0 U8 ( .IN1(n28), .IN2(in2[8]), .QN(n29) );
  NAND2X0 U9 ( .IN1(n34), .IN2(in2[10]), .QN(n35) );
  NAND2X0 U10 ( .IN1(n40), .IN2(in2[12]), .QN(n41) );
  NAND2X0 U11 ( .IN1(n43), .IN2(in2[13]), .QN(n44) );
  NAND2X0 U12 ( .IN1(n46), .IN2(in2[14]), .QN(n47) );
  NAND2X0 U13 ( .IN1(n52), .IN2(in2[16]), .QN(n53) );
  NAND2X0 U14 ( .IN1(n55), .IN2(in2[17]), .QN(n56) );
  NAND2X0 U15 ( .IN1(n7), .IN2(n15), .QN(out1[1]) );
  NAND2X0 U16 ( .IN1(n10), .IN2(n9), .QN(out1[2]) );
  NAND2X0 U17 ( .IN1(n61), .IN2(in2[19]), .QN(n62) );
  NAND2X0 U18 ( .IN1(in1[1]), .IN2(in1[0]), .QN(out1[25]) );
  NOR2X0 U19 ( .IN1(in1[1]), .IN2(in1[0]), .QN(n71) );
  INVX0 U20 ( .INP(in2[0]), .ZN(n1) );
  INVX0 U21 ( .INP(in2[1]), .ZN(n2) );
  INVX0 U22 ( .INP(in2[3]), .ZN(n3) );
  INVX0 U23 ( .INP(in2[21]), .ZN(n4) );
  INVX0 U24 ( .INP(in2[22]), .ZN(n5) );
  INVX0 U25 ( .INP(in1[1]), .ZN(n6) );
  MUX21X1 U26 ( .IN1(in1[1]), .IN2(n6), .S(in1[0]), .Q(n74) );
  INVX0 U27 ( .INP(n74), .ZN(n76) );
  AO221X1 U28 ( .IN1(in2[0]), .IN2(in2[1]), .IN3(n1), .IN4(n2), .IN5(n76), .Q(
        n7) );
  MUX21X1 U29 ( .IN1(n2), .IN2(n8), .S(in2[2]), .Q(n12) );
  AO221X1 U30 ( .IN1(n12), .IN2(in2[2]), .IN3(n12), .IN4(n1), .IN5(n76), .Q(
        n10) );
  INVX0 U31 ( .INP(n71), .ZN(n13) );
  AO221X1 U32 ( .IN1(in2[0]), .IN2(in2[1]), .IN3(n1), .IN4(n2), .IN5(n13), .Q(
        n9) );
  NOR3X0 U33 ( .IN1(in2[0]), .IN2(in2[2]), .IN3(in2[1]), .QN(n11) );
  OR4X1 U34 ( .IN1(in2[3]), .IN2(in2[0]), .IN3(in2[2]), .IN4(in2[1]), .Q(n16)
         );
  OA21X1 U35 ( .IN1(n11), .IN2(n3), .IN3(n16), .Q(n18) );
  INVX0 U36 ( .INP(n18), .ZN(n14) );
  OAI222X1 U37 ( .IN1(n15), .IN2(in2[2]), .IN3(n14), .IN4(n76), .IN5(n13), 
        .IN6(n12), .QN(out1[3]) );
  OR2X1 U38 ( .IN1(in2[4]), .IN2(n16), .Q(n19) );
  AND2X1 U39 ( .IN1(n19), .IN2(n17), .Q(n21) );
  AO22X1 U40 ( .IN1(n71), .IN2(n18), .IN3(n21), .IN4(n74), .Q(out1[4]) );
  OR2X1 U41 ( .IN1(in2[5]), .IN2(n19), .Q(n22) );
  AND2X1 U42 ( .IN1(n22), .IN2(n20), .Q(n24) );
  AO22X1 U43 ( .IN1(n71), .IN2(n21), .IN3(n24), .IN4(n74), .Q(out1[5]) );
  OR2X1 U44 ( .IN1(in2[6]), .IN2(n22), .Q(n25) );
  NAND2X0 U45 ( .IN1(n22), .IN2(in2[6]), .QN(n23) );
  AND2X1 U46 ( .IN1(n25), .IN2(n23), .Q(n27) );
  AO22X1 U47 ( .IN1(n71), .IN2(n24), .IN3(n27), .IN4(n74), .Q(out1[6]) );
  OR2X1 U48 ( .IN1(in2[7]), .IN2(n25), .Q(n28) );
  AND2X1 U49 ( .IN1(n28), .IN2(n26), .Q(n30) );
  AO22X1 U50 ( .IN1(n71), .IN2(n27), .IN3(n30), .IN4(n74), .Q(out1[7]) );
  OR2X1 U51 ( .IN1(in2[8]), .IN2(n28), .Q(n31) );
  AND2X1 U52 ( .IN1(n31), .IN2(n29), .Q(n33) );
  AO22X1 U53 ( .IN1(n71), .IN2(n30), .IN3(n33), .IN4(n74), .Q(out1[8]) );
  OR2X1 U54 ( .IN1(in2[9]), .IN2(n31), .Q(n34) );
  NAND2X0 U55 ( .IN1(n31), .IN2(in2[9]), .QN(n32) );
  AND2X1 U56 ( .IN1(n34), .IN2(n32), .Q(n36) );
  AO22X1 U57 ( .IN1(n71), .IN2(n33), .IN3(n36), .IN4(n74), .Q(out1[9]) );
  OR2X1 U58 ( .IN1(in2[10]), .IN2(n34), .Q(n37) );
  AND2X1 U59 ( .IN1(n37), .IN2(n35), .Q(n39) );
  AO22X1 U60 ( .IN1(n71), .IN2(n36), .IN3(n39), .IN4(n74), .Q(out1[10]) );
  OR2X1 U61 ( .IN1(in2[11]), .IN2(n37), .Q(n40) );
  NAND2X0 U62 ( .IN1(n37), .IN2(in2[11]), .QN(n38) );
  AND2X1 U63 ( .IN1(n40), .IN2(n38), .Q(n42) );
  AO22X1 U64 ( .IN1(n71), .IN2(n39), .IN3(n42), .IN4(n74), .Q(out1[11]) );
  OR2X1 U65 ( .IN1(in2[12]), .IN2(n40), .Q(n43) );
  AND2X1 U66 ( .IN1(n43), .IN2(n41), .Q(n45) );
  AO22X1 U67 ( .IN1(n71), .IN2(n42), .IN3(n45), .IN4(n74), .Q(out1[12]) );
  OR2X1 U68 ( .IN1(in2[13]), .IN2(n43), .Q(n46) );
  AND2X1 U69 ( .IN1(n46), .IN2(n44), .Q(n48) );
  AO22X1 U70 ( .IN1(n71), .IN2(n45), .IN3(n48), .IN4(n74), .Q(out1[13]) );
  OR2X1 U71 ( .IN1(in2[14]), .IN2(n46), .Q(n49) );
  AND2X1 U72 ( .IN1(n49), .IN2(n47), .Q(n51) );
  AO22X1 U73 ( .IN1(n71), .IN2(n48), .IN3(n51), .IN4(n74), .Q(out1[14]) );
  OR2X1 U74 ( .IN1(in2[15]), .IN2(n49), .Q(n52) );
  NAND2X0 U75 ( .IN1(n49), .IN2(in2[15]), .QN(n50) );
  AND2X1 U76 ( .IN1(n52), .IN2(n50), .Q(n54) );
  AO22X1 U77 ( .IN1(n71), .IN2(n51), .IN3(n54), .IN4(n74), .Q(out1[15]) );
  OR2X1 U78 ( .IN1(in2[16]), .IN2(n52), .Q(n55) );
  AND2X1 U79 ( .IN1(n55), .IN2(n53), .Q(n57) );
  AO22X1 U80 ( .IN1(n71), .IN2(n54), .IN3(n57), .IN4(n74), .Q(out1[16]) );
  OR2X1 U81 ( .IN1(in2[17]), .IN2(n55), .Q(n58) );
  AND2X1 U82 ( .IN1(n58), .IN2(n56), .Q(n60) );
  AO22X1 U83 ( .IN1(n71), .IN2(n57), .IN3(n60), .IN4(n74), .Q(out1[17]) );
  OR2X1 U84 ( .IN1(in2[18]), .IN2(n58), .Q(n61) );
  NAND2X0 U85 ( .IN1(n58), .IN2(in2[18]), .QN(n59) );
  AND2X1 U86 ( .IN1(n61), .IN2(n59), .Q(n63) );
  AO22X1 U87 ( .IN1(n71), .IN2(n60), .IN3(n63), .IN4(n74), .Q(out1[18]) );
  OR2X1 U88 ( .IN1(in2[19]), .IN2(n61), .Q(n64) );
  AND2X1 U89 ( .IN1(n64), .IN2(n62), .Q(n65) );
  AO22X1 U90 ( .IN1(n71), .IN2(n63), .IN3(n65), .IN4(n74), .Q(out1[19]) );
  NOR2X0 U91 ( .IN1(in2[20]), .IN2(n64), .QN(n72) );
  AOI21X1 U92 ( .IN1(in2[20]), .IN2(n64), .IN3(n72), .QN(n66) );
  AO22X1 U93 ( .IN1(n71), .IN2(n65), .IN3(n66), .IN4(n74), .Q(out1[20]) );
  MUX21X1 U94 ( .IN1(n4), .IN2(in2[21]), .S(n72), .Q(n69) );
  AO22X1 U95 ( .IN1(n71), .IN2(n66), .IN3(n69), .IN4(n74), .Q(out1[21]) );
  INVX0 U96 ( .INP(n72), .ZN(n67) );
  NOR2X0 U97 ( .IN1(in2[21]), .IN2(n67), .QN(n70) );
  MUX21X1 U98 ( .IN1(n5), .IN2(in2[22]), .S(n70), .Q(n68) );
  AO22X1 U99 ( .IN1(n71), .IN2(n69), .IN3(n68), .IN4(n74), .Q(out1[22]) );
  MUX21X1 U100 ( .IN1(n71), .IN2(n74), .S(n70), .Q(n73) );
  AND3X1 U101 ( .IN1(n72), .IN2(n71), .IN3(n4), .Q(n75) );
  MUX21X1 U102 ( .IN1(n73), .IN2(n75), .S(in2[22]), .Q(out1[23]) );
  AO21X1 U103 ( .IN1(n75), .IN2(n5), .IN3(n74), .Q(out1[24]) );
  NOR2X0 U104 ( .IN1(n76), .IN2(n1), .QN(out1[0]) );
endmodule


module booth27_3 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n25), .IN2(n6), .QN(n30) );
  NAND2X0 U4 ( .IN1(n33), .IN2(n7), .QN(n37) );
  NAND2X0 U5 ( .IN1(n41), .IN2(n8), .QN(n45) );
  NAND2X0 U6 ( .IN1(n49), .IN2(n9), .QN(n53) );
  NAND2X0 U7 ( .IN1(n57), .IN2(n10), .QN(n61) );
  NAND2X0 U8 ( .IN1(n65), .IN2(n11), .QN(n77) );
  NAND2X0 U9 ( .IN1(n81), .IN2(n13), .QN(n89) );
  NAND2X0 U10 ( .IN1(n93), .IN2(n15), .QN(n101) );
  NAND2X0 U11 ( .IN1(n105), .IN2(n17), .QN(n114) );
  NAND2X0 U12 ( .IN1(n27), .IN2(n132), .QN(n4) );
  NAND2X0 U13 ( .IN1(in1[2]), .IN2(n77), .QN(n71) );
  NAND2X0 U14 ( .IN1(n70), .IN2(n132), .QN(n74) );
  NAND2X0 U15 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U16 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U17 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U18 ( .IN1(n118), .IN2(n19), .QN(n125) );
  NAND2X0 U19 ( .IN1(n141), .IN2(n130), .QN(n24) );
  NAND2X0 U20 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NAND2X0 U21 ( .IN1(n32), .IN2(n31), .QN(out1[3]) );
  NAND2X0 U22 ( .IN1(n36), .IN2(n35), .QN(out1[4]) );
  NAND2X0 U23 ( .IN1(n40), .IN2(n39), .QN(out1[5]) );
  NAND2X0 U24 ( .IN1(n44), .IN2(n43), .QN(out1[6]) );
  NAND2X0 U25 ( .IN1(n48), .IN2(n47), .QN(out1[7]) );
  NAND2X0 U26 ( .IN1(n52), .IN2(n51), .QN(out1[8]) );
  NAND2X0 U27 ( .IN1(n56), .IN2(n55), .QN(out1[9]) );
  NAND2X0 U28 ( .IN1(n60), .IN2(n59), .QN(out1[10]) );
  NAND2X0 U29 ( .IN1(n64), .IN2(n63), .QN(out1[11]) );
  NAND2X0 U30 ( .IN1(n69), .IN2(n68), .QN(out1[12]) );
  NAND2X0 U31 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U32 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U33 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U34 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U35 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U36 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U37 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U38 ( .IN1(n23), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U39 ( .IN1(in1[2]), .IN2(n22), .QN(n23) );
  NOR2X0 U40 ( .IN1(n28), .IN2(n26), .QN(n3) );
  NOR2X0 U41 ( .IN1(n142), .IN2(n21), .QN(n1) );
  NOR2X0 U42 ( .IN1(n142), .IN2(n111), .QN(n138) );
  INVX0 U43 ( .INP(n130), .ZN(n137) );
  INVX0 U44 ( .INP(n132), .ZN(n141) );
  NOR3X0 U45 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  NAND3X0 U46 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  MUX21X1 U47 ( .IN1(n22), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  INVX0 U48 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U49 ( .INP(in2[2]), .ZN(n6) );
  INVX0 U50 ( .INP(in2[4]), .ZN(n7) );
  INVX0 U51 ( .INP(in2[6]), .ZN(n8) );
  INVX0 U52 ( .INP(in2[8]), .ZN(n9) );
  INVX0 U53 ( .INP(in2[10]), .ZN(n10) );
  INVX0 U54 ( .INP(in2[12]), .ZN(n11) );
  INVX0 U55 ( .INP(in2[13]), .ZN(n12) );
  INVX0 U56 ( .INP(in2[14]), .ZN(n13) );
  INVX0 U57 ( .INP(in2[15]), .ZN(n14) );
  INVX0 U58 ( .INP(in2[16]), .ZN(n15) );
  INVX0 U59 ( .INP(in2[17]), .ZN(n16) );
  INVX0 U60 ( .INP(in2[18]), .ZN(n17) );
  INVX0 U61 ( .INP(in2[19]), .ZN(n18) );
  INVX0 U62 ( .INP(in2[20]), .ZN(n19) );
  INVX0 U63 ( .INP(in2[21]), .ZN(n20) );
  INVX0 U64 ( .INP(in2[22]), .ZN(n21) );
  INVX0 U65 ( .INP(in1[1]), .ZN(n22) );
  INVX0 U66 ( .INP(in1[2]), .ZN(n111) );
  INVX0 U67 ( .INP(n138), .ZN(n140) );
  NOR2X0 U68 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n25) );
  AOI21X1 U69 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n25), .QN(n27) );
  NOR2X0 U70 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U71 ( .IN1(n24), .IN2(in2[0]), .IN3(n138), .IN4(n27), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U72 ( .INP(n133), .ZN(n67) );
  NOR2X0 U73 ( .IN1(n67), .IN2(n6), .QN(n28) );
  OA21X1 U74 ( .IN1(n25), .IN2(n6), .IN3(n30), .Q(n29) );
  AO22X1 U75 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n29), .Q(n26) );
  AOI22X1 U76 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n29), .QN(n32) );
  NOR2X0 U77 ( .IN1(in2[3]), .IN2(n30), .QN(n33) );
  AO21X1 U78 ( .IN1(in2[3]), .IN2(n30), .IN3(n33), .Q(n34) );
  OA22X1 U79 ( .IN1(n6), .IN2(n130), .IN3(n140), .IN4(n34), .Q(n31) );
  OA21X1 U80 ( .IN1(n33), .IN2(n7), .IN3(n37), .Q(n38) );
  AOI22X1 U81 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n38), .QN(n36) );
  OA22X1 U82 ( .IN1(n67), .IN2(n7), .IN3(n141), .IN4(n34), .Q(n35) );
  NOR2X0 U83 ( .IN1(in2[5]), .IN2(n37), .QN(n41) );
  AO21X1 U84 ( .IN1(in2[5]), .IN2(n37), .IN3(n41), .Q(n42) );
  OA22X1 U85 ( .IN1(n7), .IN2(n130), .IN3(n140), .IN4(n42), .Q(n40) );
  AOI22X1 U86 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n38), .QN(n39) );
  OA21X1 U87 ( .IN1(n41), .IN2(n8), .IN3(n45), .Q(n46) );
  AOI22X1 U88 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n46), .QN(n44) );
  OA22X1 U89 ( .IN1(n67), .IN2(n8), .IN3(n141), .IN4(n42), .Q(n43) );
  NOR2X0 U90 ( .IN1(in2[7]), .IN2(n45), .QN(n49) );
  AO21X1 U91 ( .IN1(in2[7]), .IN2(n45), .IN3(n49), .Q(n50) );
  OA22X1 U92 ( .IN1(n8), .IN2(n130), .IN3(n140), .IN4(n50), .Q(n48) );
  AOI22X1 U93 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n46), .QN(n47) );
  OA21X1 U94 ( .IN1(n49), .IN2(n9), .IN3(n53), .Q(n54) );
  AOI22X1 U95 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n54), .QN(n52) );
  OA22X1 U96 ( .IN1(n67), .IN2(n9), .IN3(n141), .IN4(n50), .Q(n51) );
  NOR2X0 U97 ( .IN1(in2[9]), .IN2(n53), .QN(n57) );
  AO21X1 U98 ( .IN1(in2[9]), .IN2(n53), .IN3(n57), .Q(n58) );
  OA22X1 U99 ( .IN1(n9), .IN2(n130), .IN3(n140), .IN4(n58), .Q(n56) );
  AOI22X1 U100 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n54), .QN(n55) );
  OA21X1 U101 ( .IN1(n57), .IN2(n10), .IN3(n61), .Q(n62) );
  AOI22X1 U102 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n62), .QN(n60) );
  OA22X1 U103 ( .IN1(n67), .IN2(n10), .IN3(n141), .IN4(n58), .Q(n59) );
  NOR2X0 U104 ( .IN1(in2[11]), .IN2(n61), .QN(n65) );
  AO21X1 U105 ( .IN1(in2[11]), .IN2(n61), .IN3(n65), .Q(n66) );
  OA22X1 U106 ( .IN1(n10), .IN2(n130), .IN3(n140), .IN4(n66), .Q(n64) );
  AOI22X1 U107 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n62), .QN(n63) );
  OA21X1 U108 ( .IN1(n65), .IN2(n11), .IN3(n77), .Q(n70) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n70), .QN(n69) );
  OA22X1 U110 ( .IN1(n67), .IN2(n11), .IN3(n141), .IN4(n66), .Q(n68) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n12), .S(n71), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n11), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n13), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n12), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n12), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n14), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n13), .IN4(n85), .IN5(n84), 
        .Q(out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n15), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n14), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n14), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n16), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n15), .IN4(n97), .IN5(n96), 
        .Q(out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n17), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n16), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n16), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n18), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n17), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n19), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n18), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n18), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n20), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n19), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n21), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n20), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n20), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n21), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_4 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n33), .IN2(n7), .QN(n37) );
  NAND2X0 U4 ( .IN1(n41), .IN2(n8), .QN(n45) );
  NAND2X0 U5 ( .IN1(n49), .IN2(n9), .QN(n53) );
  NAND2X0 U6 ( .IN1(n57), .IN2(n10), .QN(n61) );
  NAND2X0 U7 ( .IN1(n25), .IN2(n6), .QN(n30) );
  NAND2X0 U8 ( .IN1(n65), .IN2(n11), .QN(n77) );
  NAND2X0 U9 ( .IN1(n81), .IN2(n13), .QN(n89) );
  NAND2X0 U10 ( .IN1(n93), .IN2(n15), .QN(n101) );
  NAND2X0 U11 ( .IN1(n105), .IN2(n17), .QN(n114) );
  NAND2X0 U12 ( .IN1(n118), .IN2(n19), .QN(n125) );
  NAND2X0 U13 ( .IN1(in1[2]), .IN2(n77), .QN(n71) );
  NAND2X0 U14 ( .IN1(n70), .IN2(n132), .QN(n74) );
  NAND2X0 U15 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U16 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U17 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U18 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U19 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U20 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U21 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U22 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NAND2X0 U23 ( .IN1(n27), .IN2(n132), .QN(n4) );
  NAND2X0 U24 ( .IN1(n32), .IN2(n31), .QN(out1[3]) );
  NAND2X0 U25 ( .IN1(n36), .IN2(n35), .QN(out1[4]) );
  NAND2X0 U26 ( .IN1(n40), .IN2(n39), .QN(out1[5]) );
  NAND2X0 U27 ( .IN1(n44), .IN2(n43), .QN(out1[6]) );
  NAND2X0 U28 ( .IN1(n48), .IN2(n47), .QN(out1[7]) );
  NAND2X0 U29 ( .IN1(n52), .IN2(n51), .QN(out1[8]) );
  NAND2X0 U30 ( .IN1(n56), .IN2(n55), .QN(out1[9]) );
  NAND2X0 U31 ( .IN1(n60), .IN2(n59), .QN(out1[10]) );
  NAND2X0 U32 ( .IN1(n64), .IN2(n63), .QN(out1[11]) );
  NAND2X0 U33 ( .IN1(n69), .IN2(n68), .QN(out1[12]) );
  NAND2X0 U34 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U35 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U36 ( .IN1(n141), .IN2(n130), .QN(n24) );
  NAND2X0 U37 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U38 ( .IN1(n23), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U39 ( .IN1(in1[2]), .IN2(n22), .QN(n23) );
  NOR2X0 U40 ( .IN1(n28), .IN2(n26), .QN(n3) );
  NOR2X0 U41 ( .IN1(n142), .IN2(n111), .QN(n138) );
  NOR2X0 U42 ( .IN1(n142), .IN2(n21), .QN(n1) );
  INVX0 U43 ( .INP(n130), .ZN(n137) );
  INVX0 U44 ( .INP(n132), .ZN(n141) );
  NOR3X0 U45 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  NAND3X0 U46 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  MUX21X1 U47 ( .IN1(n22), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  INVX0 U48 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U49 ( .INP(in2[2]), .ZN(n6) );
  INVX0 U50 ( .INP(in2[4]), .ZN(n7) );
  INVX0 U51 ( .INP(in2[6]), .ZN(n8) );
  INVX0 U52 ( .INP(in2[8]), .ZN(n9) );
  INVX0 U53 ( .INP(in2[10]), .ZN(n10) );
  INVX0 U54 ( .INP(in2[12]), .ZN(n11) );
  INVX0 U55 ( .INP(in2[13]), .ZN(n12) );
  INVX0 U56 ( .INP(in2[14]), .ZN(n13) );
  INVX0 U57 ( .INP(in2[15]), .ZN(n14) );
  INVX0 U58 ( .INP(in2[16]), .ZN(n15) );
  INVX0 U59 ( .INP(in2[17]), .ZN(n16) );
  INVX0 U60 ( .INP(in2[18]), .ZN(n17) );
  INVX0 U61 ( .INP(in2[19]), .ZN(n18) );
  INVX0 U62 ( .INP(in2[20]), .ZN(n19) );
  INVX0 U63 ( .INP(in2[21]), .ZN(n20) );
  INVX0 U64 ( .INP(in2[22]), .ZN(n21) );
  INVX0 U65 ( .INP(in1[1]), .ZN(n22) );
  INVX0 U66 ( .INP(in1[2]), .ZN(n111) );
  INVX0 U67 ( .INP(n138), .ZN(n140) );
  NOR2X0 U68 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n25) );
  AOI21X1 U69 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n25), .QN(n27) );
  NOR2X0 U70 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U71 ( .IN1(n24), .IN2(in2[0]), .IN3(n138), .IN4(n27), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U72 ( .INP(n133), .ZN(n67) );
  NOR2X0 U73 ( .IN1(n67), .IN2(n6), .QN(n28) );
  OA21X1 U74 ( .IN1(n25), .IN2(n6), .IN3(n30), .Q(n29) );
  AO22X1 U75 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n29), .Q(n26) );
  AOI22X1 U76 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n29), .QN(n32) );
  NOR2X0 U77 ( .IN1(in2[3]), .IN2(n30), .QN(n33) );
  AO21X1 U78 ( .IN1(in2[3]), .IN2(n30), .IN3(n33), .Q(n34) );
  OA22X1 U79 ( .IN1(n6), .IN2(n130), .IN3(n140), .IN4(n34), .Q(n31) );
  OA21X1 U80 ( .IN1(n33), .IN2(n7), .IN3(n37), .Q(n38) );
  AOI22X1 U81 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n38), .QN(n36) );
  OA22X1 U82 ( .IN1(n67), .IN2(n7), .IN3(n141), .IN4(n34), .Q(n35) );
  NOR2X0 U83 ( .IN1(in2[5]), .IN2(n37), .QN(n41) );
  AO21X1 U84 ( .IN1(in2[5]), .IN2(n37), .IN3(n41), .Q(n42) );
  OA22X1 U85 ( .IN1(n7), .IN2(n130), .IN3(n140), .IN4(n42), .Q(n40) );
  AOI22X1 U86 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n38), .QN(n39) );
  OA21X1 U87 ( .IN1(n41), .IN2(n8), .IN3(n45), .Q(n46) );
  AOI22X1 U88 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n46), .QN(n44) );
  OA22X1 U89 ( .IN1(n67), .IN2(n8), .IN3(n141), .IN4(n42), .Q(n43) );
  NOR2X0 U90 ( .IN1(in2[7]), .IN2(n45), .QN(n49) );
  AO21X1 U91 ( .IN1(in2[7]), .IN2(n45), .IN3(n49), .Q(n50) );
  OA22X1 U92 ( .IN1(n8), .IN2(n130), .IN3(n140), .IN4(n50), .Q(n48) );
  AOI22X1 U93 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n46), .QN(n47) );
  OA21X1 U94 ( .IN1(n49), .IN2(n9), .IN3(n53), .Q(n54) );
  AOI22X1 U95 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n54), .QN(n52) );
  OA22X1 U96 ( .IN1(n67), .IN2(n9), .IN3(n141), .IN4(n50), .Q(n51) );
  NOR2X0 U97 ( .IN1(in2[9]), .IN2(n53), .QN(n57) );
  AO21X1 U98 ( .IN1(in2[9]), .IN2(n53), .IN3(n57), .Q(n58) );
  OA22X1 U99 ( .IN1(n9), .IN2(n130), .IN3(n140), .IN4(n58), .Q(n56) );
  AOI22X1 U100 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n54), .QN(n55) );
  OA21X1 U101 ( .IN1(n57), .IN2(n10), .IN3(n61), .Q(n62) );
  AOI22X1 U102 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n62), .QN(n60) );
  OA22X1 U103 ( .IN1(n67), .IN2(n10), .IN3(n141), .IN4(n58), .Q(n59) );
  NOR2X0 U104 ( .IN1(in2[11]), .IN2(n61), .QN(n65) );
  AO21X1 U105 ( .IN1(in2[11]), .IN2(n61), .IN3(n65), .Q(n66) );
  OA22X1 U106 ( .IN1(n10), .IN2(n130), .IN3(n140), .IN4(n66), .Q(n64) );
  AOI22X1 U107 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n62), .QN(n63) );
  OA21X1 U108 ( .IN1(n65), .IN2(n11), .IN3(n77), .Q(n70) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n70), .QN(n69) );
  OA22X1 U110 ( .IN1(n67), .IN2(n11), .IN3(n141), .IN4(n66), .Q(n68) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n12), .S(n71), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n11), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n13), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n12), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n12), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n14), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n13), .IN4(n85), .IN5(n84), 
        .Q(out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n15), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n14), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n14), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n16), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n15), .IN4(n97), .IN5(n96), 
        .Q(out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n17), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n16), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n16), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n18), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n17), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n19), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n18), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n18), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n20), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n19), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n21), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n20), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n20), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n21), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_5 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n41), .IN2(n8), .QN(n45) );
  NAND2X0 U4 ( .IN1(n49), .IN2(n9), .QN(n53) );
  NAND2X0 U5 ( .IN1(n57), .IN2(n10), .QN(n61) );
  NAND2X0 U6 ( .IN1(n33), .IN2(n7), .QN(n37) );
  NAND2X0 U7 ( .IN1(n25), .IN2(n6), .QN(n30) );
  NAND2X0 U8 ( .IN1(n65), .IN2(n11), .QN(n77) );
  NAND2X0 U9 ( .IN1(n81), .IN2(n13), .QN(n89) );
  NAND2X0 U10 ( .IN1(n93), .IN2(n15), .QN(n101) );
  NAND2X0 U11 ( .IN1(in1[2]), .IN2(n77), .QN(n71) );
  NAND2X0 U12 ( .IN1(n70), .IN2(n132), .QN(n74) );
  NAND2X0 U13 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U14 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U15 ( .IN1(n105), .IN2(n17), .QN(n114) );
  NAND2X0 U16 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U17 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U18 ( .IN1(n27), .IN2(n132), .QN(n4) );
  NAND2X0 U19 ( .IN1(n141), .IN2(n130), .QN(n24) );
  NAND2X0 U20 ( .IN1(n40), .IN2(n39), .QN(out1[5]) );
  NAND2X0 U21 ( .IN1(n44), .IN2(n43), .QN(out1[6]) );
  NAND2X0 U22 ( .IN1(n48), .IN2(n47), .QN(out1[7]) );
  NAND2X0 U23 ( .IN1(n52), .IN2(n51), .QN(out1[8]) );
  NAND2X0 U24 ( .IN1(n56), .IN2(n55), .QN(out1[9]) );
  NAND2X0 U25 ( .IN1(n60), .IN2(n59), .QN(out1[10]) );
  NAND2X0 U26 ( .IN1(n64), .IN2(n63), .QN(out1[11]) );
  NAND2X0 U27 ( .IN1(n69), .IN2(n68), .QN(out1[12]) );
  NAND2X0 U28 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U29 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U30 ( .IN1(n118), .IN2(n19), .QN(n125) );
  NAND2X0 U31 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U32 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U33 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U34 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U35 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NAND2X0 U36 ( .IN1(n32), .IN2(n31), .QN(out1[3]) );
  NAND2X0 U37 ( .IN1(n36), .IN2(n35), .QN(out1[4]) );
  NAND2X0 U38 ( .IN1(n23), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U39 ( .IN1(in1[2]), .IN2(n22), .QN(n23) );
  INVX0 U40 ( .INP(in1[2]), .ZN(n111) );
  NOR2X0 U41 ( .IN1(n28), .IN2(n26), .QN(n3) );
  NOR2X0 U42 ( .IN1(n142), .IN2(n21), .QN(n1) );
  INVX0 U43 ( .INP(n132), .ZN(n141) );
  INVX0 U44 ( .INP(n130), .ZN(n137) );
  NOR2X0 U45 ( .IN1(n142), .IN2(n111), .QN(n138) );
  MUX21X1 U46 ( .IN1(n22), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  NAND3X0 U47 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  NOR3X0 U48 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  INVX0 U49 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U50 ( .INP(in2[2]), .ZN(n6) );
  INVX0 U51 ( .INP(in2[4]), .ZN(n7) );
  INVX0 U52 ( .INP(in2[6]), .ZN(n8) );
  INVX0 U53 ( .INP(in2[8]), .ZN(n9) );
  INVX0 U54 ( .INP(in2[10]), .ZN(n10) );
  INVX0 U55 ( .INP(in2[12]), .ZN(n11) );
  INVX0 U56 ( .INP(in2[13]), .ZN(n12) );
  INVX0 U57 ( .INP(in2[14]), .ZN(n13) );
  INVX0 U58 ( .INP(in2[15]), .ZN(n14) );
  INVX0 U59 ( .INP(in2[16]), .ZN(n15) );
  INVX0 U60 ( .INP(in2[17]), .ZN(n16) );
  INVX0 U61 ( .INP(in2[18]), .ZN(n17) );
  INVX0 U62 ( .INP(in2[19]), .ZN(n18) );
  INVX0 U63 ( .INP(in2[20]), .ZN(n19) );
  INVX0 U64 ( .INP(in2[21]), .ZN(n20) );
  INVX0 U65 ( .INP(in2[22]), .ZN(n21) );
  INVX0 U66 ( .INP(in1[1]), .ZN(n22) );
  INVX0 U67 ( .INP(n138), .ZN(n140) );
  NOR2X0 U68 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n25) );
  AOI21X1 U69 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n25), .QN(n27) );
  NOR2X0 U70 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U71 ( .IN1(n24), .IN2(in2[0]), .IN3(n138), .IN4(n27), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U72 ( .INP(n133), .ZN(n67) );
  NOR2X0 U73 ( .IN1(n67), .IN2(n6), .QN(n28) );
  OA21X1 U74 ( .IN1(n25), .IN2(n6), .IN3(n30), .Q(n29) );
  AO22X1 U75 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n29), .Q(n26) );
  AOI22X1 U76 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n29), .QN(n32) );
  NOR2X0 U77 ( .IN1(in2[3]), .IN2(n30), .QN(n33) );
  AO21X1 U78 ( .IN1(in2[3]), .IN2(n30), .IN3(n33), .Q(n34) );
  OA22X1 U79 ( .IN1(n6), .IN2(n130), .IN3(n140), .IN4(n34), .Q(n31) );
  OA21X1 U80 ( .IN1(n33), .IN2(n7), .IN3(n37), .Q(n38) );
  AOI22X1 U81 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n38), .QN(n36) );
  OA22X1 U82 ( .IN1(n67), .IN2(n7), .IN3(n141), .IN4(n34), .Q(n35) );
  NOR2X0 U83 ( .IN1(in2[5]), .IN2(n37), .QN(n41) );
  AO21X1 U84 ( .IN1(in2[5]), .IN2(n37), .IN3(n41), .Q(n42) );
  OA22X1 U85 ( .IN1(n7), .IN2(n130), .IN3(n140), .IN4(n42), .Q(n40) );
  AOI22X1 U86 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n38), .QN(n39) );
  OA21X1 U87 ( .IN1(n41), .IN2(n8), .IN3(n45), .Q(n46) );
  AOI22X1 U88 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n46), .QN(n44) );
  OA22X1 U89 ( .IN1(n67), .IN2(n8), .IN3(n141), .IN4(n42), .Q(n43) );
  NOR2X0 U90 ( .IN1(in2[7]), .IN2(n45), .QN(n49) );
  AO21X1 U91 ( .IN1(in2[7]), .IN2(n45), .IN3(n49), .Q(n50) );
  OA22X1 U92 ( .IN1(n8), .IN2(n130), .IN3(n140), .IN4(n50), .Q(n48) );
  AOI22X1 U93 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n46), .QN(n47) );
  OA21X1 U94 ( .IN1(n49), .IN2(n9), .IN3(n53), .Q(n54) );
  AOI22X1 U95 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n54), .QN(n52) );
  OA22X1 U96 ( .IN1(n67), .IN2(n9), .IN3(n141), .IN4(n50), .Q(n51) );
  NOR2X0 U97 ( .IN1(in2[9]), .IN2(n53), .QN(n57) );
  AO21X1 U98 ( .IN1(in2[9]), .IN2(n53), .IN3(n57), .Q(n58) );
  OA22X1 U99 ( .IN1(n9), .IN2(n130), .IN3(n140), .IN4(n58), .Q(n56) );
  AOI22X1 U100 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n54), .QN(n55) );
  OA21X1 U101 ( .IN1(n57), .IN2(n10), .IN3(n61), .Q(n62) );
  AOI22X1 U102 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n62), .QN(n60) );
  OA22X1 U103 ( .IN1(n67), .IN2(n10), .IN3(n141), .IN4(n58), .Q(n59) );
  NOR2X0 U104 ( .IN1(in2[11]), .IN2(n61), .QN(n65) );
  AO21X1 U105 ( .IN1(in2[11]), .IN2(n61), .IN3(n65), .Q(n66) );
  OA22X1 U106 ( .IN1(n10), .IN2(n130), .IN3(n140), .IN4(n66), .Q(n64) );
  AOI22X1 U107 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n62), .QN(n63) );
  OA21X1 U108 ( .IN1(n65), .IN2(n11), .IN3(n77), .Q(n70) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n70), .QN(n69) );
  OA22X1 U110 ( .IN1(n67), .IN2(n11), .IN3(n141), .IN4(n66), .Q(n68) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n12), .S(n71), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n11), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n13), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n12), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n12), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n14), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n13), .IN4(n85), .IN5(n84), 
        .Q(out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n15), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n14), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n14), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n16), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n15), .IN4(n97), .IN5(n96), 
        .Q(out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n17), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n16), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n16), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n18), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n17), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n19), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n18), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n18), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n20), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n19), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n21), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n20), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n20), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n21), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_6 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n49), .IN2(n9), .QN(n53) );
  NAND2X0 U4 ( .IN1(n57), .IN2(n10), .QN(n61) );
  NAND2X0 U5 ( .IN1(n25), .IN2(n6), .QN(n30) );
  NAND2X0 U6 ( .IN1(n41), .IN2(n8), .QN(n45) );
  NAND2X0 U7 ( .IN1(n33), .IN2(n7), .QN(n37) );
  NAND2X0 U8 ( .IN1(n65), .IN2(n11), .QN(n77) );
  NAND2X0 U9 ( .IN1(n81), .IN2(n13), .QN(n89) );
  NAND2X0 U10 ( .IN1(n93), .IN2(n15), .QN(n101) );
  NAND2X0 U11 ( .IN1(n105), .IN2(n17), .QN(n114) );
  NAND2X0 U12 ( .IN1(in1[2]), .IN2(n77), .QN(n71) );
  NAND2X0 U13 ( .IN1(n70), .IN2(n132), .QN(n74) );
  NAND2X0 U14 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U15 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U16 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U17 ( .IN1(n118), .IN2(n19), .QN(n125) );
  NAND2X0 U18 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U19 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U20 ( .IN1(n27), .IN2(n132), .QN(n4) );
  NAND2X0 U21 ( .IN1(n48), .IN2(n47), .QN(out1[7]) );
  NAND2X0 U22 ( .IN1(n52), .IN2(n51), .QN(out1[8]) );
  NAND2X0 U23 ( .IN1(n56), .IN2(n55), .QN(out1[9]) );
  NAND2X0 U24 ( .IN1(n60), .IN2(n59), .QN(out1[10]) );
  NAND2X0 U25 ( .IN1(n64), .IN2(n63), .QN(out1[11]) );
  NAND2X0 U26 ( .IN1(n69), .IN2(n68), .QN(out1[12]) );
  NAND2X0 U27 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U28 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U29 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U30 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U31 ( .IN1(n141), .IN2(n130), .QN(n24) );
  NAND2X0 U32 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NAND2X0 U33 ( .IN1(n36), .IN2(n35), .QN(out1[4]) );
  NAND2X0 U34 ( .IN1(n32), .IN2(n31), .QN(out1[3]) );
  NAND2X0 U35 ( .IN1(n40), .IN2(n39), .QN(out1[5]) );
  NAND2X0 U36 ( .IN1(n44), .IN2(n43), .QN(out1[6]) );
  NAND2X0 U37 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U38 ( .IN1(n23), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U39 ( .IN1(in1[2]), .IN2(n22), .QN(n23) );
  NOR2X0 U40 ( .IN1(n28), .IN2(n26), .QN(n3) );
  INVX0 U41 ( .INP(n130), .ZN(n137) );
  NAND3X0 U42 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  NOR2X0 U43 ( .IN1(n142), .IN2(n21), .QN(n1) );
  NOR2X0 U44 ( .IN1(n142), .IN2(n111), .QN(n138) );
  MUX21X1 U45 ( .IN1(n22), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  INVX0 U46 ( .INP(n132), .ZN(n141) );
  NOR3X0 U47 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  INVX0 U48 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U49 ( .INP(in2[2]), .ZN(n6) );
  INVX0 U50 ( .INP(in2[4]), .ZN(n7) );
  INVX0 U51 ( .INP(in2[6]), .ZN(n8) );
  INVX0 U52 ( .INP(in2[8]), .ZN(n9) );
  INVX0 U53 ( .INP(in2[10]), .ZN(n10) );
  INVX0 U54 ( .INP(in2[12]), .ZN(n11) );
  INVX0 U55 ( .INP(in2[13]), .ZN(n12) );
  INVX0 U56 ( .INP(in2[14]), .ZN(n13) );
  INVX0 U57 ( .INP(in2[15]), .ZN(n14) );
  INVX0 U58 ( .INP(in2[16]), .ZN(n15) );
  INVX0 U59 ( .INP(in2[17]), .ZN(n16) );
  INVX0 U60 ( .INP(in2[18]), .ZN(n17) );
  INVX0 U61 ( .INP(in2[19]), .ZN(n18) );
  INVX0 U62 ( .INP(in2[20]), .ZN(n19) );
  INVX0 U63 ( .INP(in2[21]), .ZN(n20) );
  INVX0 U64 ( .INP(in2[22]), .ZN(n21) );
  INVX0 U65 ( .INP(in1[1]), .ZN(n22) );
  INVX0 U66 ( .INP(in1[2]), .ZN(n111) );
  INVX0 U67 ( .INP(n138), .ZN(n140) );
  NOR2X0 U68 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n25) );
  AOI21X1 U69 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n25), .QN(n27) );
  NOR2X0 U70 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U71 ( .IN1(n24), .IN2(in2[0]), .IN3(n138), .IN4(n27), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U72 ( .INP(n133), .ZN(n67) );
  NOR2X0 U73 ( .IN1(n67), .IN2(n6), .QN(n28) );
  OA21X1 U74 ( .IN1(n25), .IN2(n6), .IN3(n30), .Q(n29) );
  AO22X1 U75 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n29), .Q(n26) );
  AOI22X1 U76 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n29), .QN(n32) );
  NOR2X0 U77 ( .IN1(in2[3]), .IN2(n30), .QN(n33) );
  AO21X1 U78 ( .IN1(in2[3]), .IN2(n30), .IN3(n33), .Q(n34) );
  OA22X1 U79 ( .IN1(n6), .IN2(n130), .IN3(n140), .IN4(n34), .Q(n31) );
  OA21X1 U80 ( .IN1(n33), .IN2(n7), .IN3(n37), .Q(n38) );
  AOI22X1 U81 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n38), .QN(n36) );
  OA22X1 U82 ( .IN1(n67), .IN2(n7), .IN3(n141), .IN4(n34), .Q(n35) );
  NOR2X0 U83 ( .IN1(in2[5]), .IN2(n37), .QN(n41) );
  AO21X1 U84 ( .IN1(in2[5]), .IN2(n37), .IN3(n41), .Q(n42) );
  OA22X1 U85 ( .IN1(n7), .IN2(n130), .IN3(n140), .IN4(n42), .Q(n40) );
  AOI22X1 U86 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n38), .QN(n39) );
  OA21X1 U87 ( .IN1(n41), .IN2(n8), .IN3(n45), .Q(n46) );
  AOI22X1 U88 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n46), .QN(n44) );
  OA22X1 U89 ( .IN1(n67), .IN2(n8), .IN3(n141), .IN4(n42), .Q(n43) );
  NOR2X0 U90 ( .IN1(in2[7]), .IN2(n45), .QN(n49) );
  AO21X1 U91 ( .IN1(in2[7]), .IN2(n45), .IN3(n49), .Q(n50) );
  OA22X1 U92 ( .IN1(n8), .IN2(n130), .IN3(n140), .IN4(n50), .Q(n48) );
  AOI22X1 U93 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n46), .QN(n47) );
  OA21X1 U94 ( .IN1(n49), .IN2(n9), .IN3(n53), .Q(n54) );
  AOI22X1 U95 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n54), .QN(n52) );
  OA22X1 U96 ( .IN1(n67), .IN2(n9), .IN3(n141), .IN4(n50), .Q(n51) );
  NOR2X0 U97 ( .IN1(in2[9]), .IN2(n53), .QN(n57) );
  AO21X1 U98 ( .IN1(in2[9]), .IN2(n53), .IN3(n57), .Q(n58) );
  OA22X1 U99 ( .IN1(n9), .IN2(n130), .IN3(n140), .IN4(n58), .Q(n56) );
  AOI22X1 U100 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n54), .QN(n55) );
  OA21X1 U101 ( .IN1(n57), .IN2(n10), .IN3(n61), .Q(n62) );
  AOI22X1 U102 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n62), .QN(n60) );
  OA22X1 U103 ( .IN1(n67), .IN2(n10), .IN3(n141), .IN4(n58), .Q(n59) );
  NOR2X0 U104 ( .IN1(in2[11]), .IN2(n61), .QN(n65) );
  AO21X1 U105 ( .IN1(in2[11]), .IN2(n61), .IN3(n65), .Q(n66) );
  OA22X1 U106 ( .IN1(n10), .IN2(n130), .IN3(n140), .IN4(n66), .Q(n64) );
  AOI22X1 U107 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n62), .QN(n63) );
  OA21X1 U108 ( .IN1(n65), .IN2(n11), .IN3(n77), .Q(n70) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n70), .QN(n69) );
  OA22X1 U110 ( .IN1(n67), .IN2(n11), .IN3(n141), .IN4(n66), .Q(n68) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n12), .S(n71), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n11), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n13), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n12), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n12), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n14), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n13), .IN4(n85), .IN5(n84), 
        .Q(out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n15), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n14), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n14), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n16), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n15), .IN4(n97), .IN5(n96), 
        .Q(out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n17), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n16), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n16), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n18), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n17), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n19), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n18), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n18), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n20), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n19), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n21), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n20), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n20), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n21), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_7 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n57), .IN2(n10), .QN(n61) );
  NAND2X0 U4 ( .IN1(n33), .IN2(n7), .QN(n37) );
  NAND2X0 U5 ( .IN1(n49), .IN2(n9), .QN(n53) );
  NAND2X0 U6 ( .IN1(n41), .IN2(n8), .QN(n45) );
  NAND2X0 U7 ( .IN1(n65), .IN2(n11), .QN(n77) );
  NAND2X0 U8 ( .IN1(n81), .IN2(n13), .QN(n89) );
  NAND2X0 U9 ( .IN1(n93), .IN2(n15), .QN(n101) );
  NAND2X0 U10 ( .IN1(n105), .IN2(n17), .QN(n114) );
  NAND2X0 U11 ( .IN1(n118), .IN2(n19), .QN(n125) );
  NAND2X0 U12 ( .IN1(n25), .IN2(n6), .QN(n30) );
  NAND2X0 U13 ( .IN1(in1[2]), .IN2(n77), .QN(n71) );
  NAND2X0 U14 ( .IN1(n70), .IN2(n132), .QN(n74) );
  NAND2X0 U15 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U16 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U17 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U18 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U19 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U20 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U21 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U22 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U23 ( .IN1(n56), .IN2(n55), .QN(out1[9]) );
  NAND2X0 U24 ( .IN1(n60), .IN2(n59), .QN(out1[10]) );
  NAND2X0 U25 ( .IN1(n64), .IN2(n63), .QN(out1[11]) );
  NAND2X0 U26 ( .IN1(n69), .IN2(n68), .QN(out1[12]) );
  NAND2X0 U27 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U28 ( .IN1(n23), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U29 ( .IN1(in1[2]), .IN2(n22), .QN(n23) );
  NAND2X0 U30 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NAND2X0 U31 ( .IN1(n27), .IN2(n132), .QN(n4) );
  NAND2X0 U32 ( .IN1(n32), .IN2(n31), .QN(out1[3]) );
  NAND2X0 U33 ( .IN1(n36), .IN2(n35), .QN(out1[4]) );
  NAND2X0 U34 ( .IN1(n44), .IN2(n43), .QN(out1[6]) );
  NAND2X0 U35 ( .IN1(n40), .IN2(n39), .QN(out1[5]) );
  NAND2X0 U36 ( .IN1(n48), .IN2(n47), .QN(out1[7]) );
  NAND2X0 U37 ( .IN1(n52), .IN2(n51), .QN(out1[8]) );
  NAND2X0 U38 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U39 ( .IN1(n141), .IN2(n130), .QN(n24) );
  NOR2X0 U40 ( .IN1(n28), .IN2(n26), .QN(n3) );
  NOR2X0 U41 ( .IN1(n142), .IN2(n21), .QN(n1) );
  INVX0 U42 ( .INP(n132), .ZN(n141) );
  INVX0 U43 ( .INP(n130), .ZN(n137) );
  NAND3X0 U44 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  NOR3X0 U45 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  NOR2X0 U46 ( .IN1(n142), .IN2(n111), .QN(n138) );
  MUX21X1 U47 ( .IN1(n22), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  INVX0 U48 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U49 ( .INP(in2[2]), .ZN(n6) );
  INVX0 U50 ( .INP(in2[4]), .ZN(n7) );
  INVX0 U51 ( .INP(in2[6]), .ZN(n8) );
  INVX0 U52 ( .INP(in2[8]), .ZN(n9) );
  INVX0 U53 ( .INP(in2[10]), .ZN(n10) );
  INVX0 U54 ( .INP(in2[12]), .ZN(n11) );
  INVX0 U55 ( .INP(in2[13]), .ZN(n12) );
  INVX0 U56 ( .INP(in2[14]), .ZN(n13) );
  INVX0 U57 ( .INP(in2[15]), .ZN(n14) );
  INVX0 U58 ( .INP(in2[16]), .ZN(n15) );
  INVX0 U59 ( .INP(in2[17]), .ZN(n16) );
  INVX0 U60 ( .INP(in2[18]), .ZN(n17) );
  INVX0 U61 ( .INP(in2[19]), .ZN(n18) );
  INVX0 U62 ( .INP(in2[20]), .ZN(n19) );
  INVX0 U63 ( .INP(in2[21]), .ZN(n20) );
  INVX0 U64 ( .INP(in2[22]), .ZN(n21) );
  INVX0 U65 ( .INP(in1[1]), .ZN(n22) );
  INVX0 U66 ( .INP(in1[2]), .ZN(n111) );
  INVX0 U67 ( .INP(n138), .ZN(n140) );
  NOR2X0 U68 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n25) );
  AOI21X1 U69 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n25), .QN(n27) );
  NOR2X0 U70 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U71 ( .IN1(n24), .IN2(in2[0]), .IN3(n138), .IN4(n27), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U72 ( .INP(n133), .ZN(n67) );
  NOR2X0 U73 ( .IN1(n67), .IN2(n6), .QN(n28) );
  OA21X1 U74 ( .IN1(n25), .IN2(n6), .IN3(n30), .Q(n29) );
  AO22X1 U75 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n29), .Q(n26) );
  AOI22X1 U76 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n29), .QN(n32) );
  NOR2X0 U77 ( .IN1(in2[3]), .IN2(n30), .QN(n33) );
  AO21X1 U78 ( .IN1(in2[3]), .IN2(n30), .IN3(n33), .Q(n34) );
  OA22X1 U79 ( .IN1(n6), .IN2(n130), .IN3(n140), .IN4(n34), .Q(n31) );
  OA21X1 U80 ( .IN1(n33), .IN2(n7), .IN3(n37), .Q(n38) );
  AOI22X1 U81 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n38), .QN(n36) );
  OA22X1 U82 ( .IN1(n67), .IN2(n7), .IN3(n141), .IN4(n34), .Q(n35) );
  NOR2X0 U83 ( .IN1(in2[5]), .IN2(n37), .QN(n41) );
  AO21X1 U84 ( .IN1(in2[5]), .IN2(n37), .IN3(n41), .Q(n42) );
  OA22X1 U85 ( .IN1(n7), .IN2(n130), .IN3(n140), .IN4(n42), .Q(n40) );
  AOI22X1 U86 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n38), .QN(n39) );
  OA21X1 U87 ( .IN1(n41), .IN2(n8), .IN3(n45), .Q(n46) );
  AOI22X1 U88 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n46), .QN(n44) );
  OA22X1 U89 ( .IN1(n67), .IN2(n8), .IN3(n141), .IN4(n42), .Q(n43) );
  NOR2X0 U90 ( .IN1(in2[7]), .IN2(n45), .QN(n49) );
  AO21X1 U91 ( .IN1(in2[7]), .IN2(n45), .IN3(n49), .Q(n50) );
  OA22X1 U92 ( .IN1(n8), .IN2(n130), .IN3(n140), .IN4(n50), .Q(n48) );
  AOI22X1 U93 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n46), .QN(n47) );
  OA21X1 U94 ( .IN1(n49), .IN2(n9), .IN3(n53), .Q(n54) );
  AOI22X1 U95 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n54), .QN(n52) );
  OA22X1 U96 ( .IN1(n67), .IN2(n9), .IN3(n141), .IN4(n50), .Q(n51) );
  NOR2X0 U97 ( .IN1(in2[9]), .IN2(n53), .QN(n57) );
  AO21X1 U98 ( .IN1(in2[9]), .IN2(n53), .IN3(n57), .Q(n58) );
  OA22X1 U99 ( .IN1(n9), .IN2(n130), .IN3(n140), .IN4(n58), .Q(n56) );
  AOI22X1 U100 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n54), .QN(n55) );
  OA21X1 U101 ( .IN1(n57), .IN2(n10), .IN3(n61), .Q(n62) );
  AOI22X1 U102 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n62), .QN(n60) );
  OA22X1 U103 ( .IN1(n67), .IN2(n10), .IN3(n141), .IN4(n58), .Q(n59) );
  NOR2X0 U104 ( .IN1(in2[11]), .IN2(n61), .QN(n65) );
  AO21X1 U105 ( .IN1(in2[11]), .IN2(n61), .IN3(n65), .Q(n66) );
  OA22X1 U106 ( .IN1(n10), .IN2(n130), .IN3(n140), .IN4(n66), .Q(n64) );
  AOI22X1 U107 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n62), .QN(n63) );
  OA21X1 U108 ( .IN1(n65), .IN2(n11), .IN3(n77), .Q(n70) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n70), .QN(n69) );
  OA22X1 U110 ( .IN1(n67), .IN2(n11), .IN3(n141), .IN4(n66), .Q(n68) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n12), .S(n71), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n11), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n13), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n12), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n12), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n14), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n13), .IN4(n85), .IN5(n84), 
        .Q(out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n15), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n14), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n14), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n16), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n15), .IN4(n97), .IN5(n96), 
        .Q(out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n17), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n16), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n16), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n18), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n17), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n19), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n18), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n18), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n20), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n19), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n21), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n20), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n20), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n21), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_8 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n57), .IN2(n10), .QN(n61) );
  NAND2X0 U4 ( .IN1(n25), .IN2(n6), .QN(n30) );
  NAND2X0 U5 ( .IN1(n33), .IN2(n7), .QN(n37) );
  NAND2X0 U6 ( .IN1(n49), .IN2(n9), .QN(n53) );
  NAND2X0 U7 ( .IN1(n41), .IN2(n8), .QN(n45) );
  NAND2X0 U8 ( .IN1(n65), .IN2(n11), .QN(n77) );
  NAND2X0 U9 ( .IN1(n81), .IN2(n13), .QN(n89) );
  NAND2X0 U10 ( .IN1(n93), .IN2(n15), .QN(n101) );
  NAND2X0 U11 ( .IN1(n105), .IN2(n17), .QN(n114) );
  NAND2X0 U12 ( .IN1(in1[2]), .IN2(n77), .QN(n71) );
  NAND2X0 U13 ( .IN1(n70), .IN2(n132), .QN(n74) );
  NAND2X0 U14 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U15 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U16 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U17 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U18 ( .IN1(n118), .IN2(n19), .QN(n125) );
  NAND2X0 U19 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U20 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U21 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U22 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U23 ( .IN1(n141), .IN2(n130), .QN(n24) );
  NAND2X0 U24 ( .IN1(n27), .IN2(n132), .QN(n4) );
  NAND2X0 U25 ( .IN1(n56), .IN2(n55), .QN(out1[9]) );
  NAND2X0 U26 ( .IN1(n60), .IN2(n59), .QN(out1[10]) );
  NAND2X0 U27 ( .IN1(n64), .IN2(n63), .QN(out1[11]) );
  NAND2X0 U28 ( .IN1(n69), .IN2(n68), .QN(out1[12]) );
  NAND2X0 U29 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U30 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U31 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NAND2X0 U32 ( .IN1(n32), .IN2(n31), .QN(out1[3]) );
  NAND2X0 U33 ( .IN1(n36), .IN2(n35), .QN(out1[4]) );
  NAND2X0 U34 ( .IN1(n40), .IN2(n39), .QN(out1[5]) );
  NAND2X0 U35 ( .IN1(n44), .IN2(n43), .QN(out1[6]) );
  NAND2X0 U36 ( .IN1(n48), .IN2(n47), .QN(out1[7]) );
  NAND2X0 U37 ( .IN1(n52), .IN2(n51), .QN(out1[8]) );
  NAND2X0 U38 ( .IN1(n23), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U39 ( .IN1(in1[2]), .IN2(n22), .QN(n23) );
  NOR2X0 U40 ( .IN1(n28), .IN2(n26), .QN(n3) );
  NOR2X0 U41 ( .IN1(n142), .IN2(n21), .QN(n1) );
  INVX0 U42 ( .INP(n132), .ZN(n141) );
  INVX0 U43 ( .INP(n130), .ZN(n137) );
  NAND3X0 U44 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  NOR3X0 U45 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  NOR2X0 U46 ( .IN1(n142), .IN2(n111), .QN(n138) );
  MUX21X1 U47 ( .IN1(n22), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  INVX0 U48 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U49 ( .INP(in2[2]), .ZN(n6) );
  INVX0 U50 ( .INP(in2[4]), .ZN(n7) );
  INVX0 U51 ( .INP(in2[6]), .ZN(n8) );
  INVX0 U52 ( .INP(in2[8]), .ZN(n9) );
  INVX0 U53 ( .INP(in2[10]), .ZN(n10) );
  INVX0 U54 ( .INP(in2[12]), .ZN(n11) );
  INVX0 U55 ( .INP(in2[13]), .ZN(n12) );
  INVX0 U56 ( .INP(in2[14]), .ZN(n13) );
  INVX0 U57 ( .INP(in2[15]), .ZN(n14) );
  INVX0 U58 ( .INP(in2[16]), .ZN(n15) );
  INVX0 U59 ( .INP(in2[17]), .ZN(n16) );
  INVX0 U60 ( .INP(in2[18]), .ZN(n17) );
  INVX0 U61 ( .INP(in2[19]), .ZN(n18) );
  INVX0 U62 ( .INP(in2[20]), .ZN(n19) );
  INVX0 U63 ( .INP(in2[21]), .ZN(n20) );
  INVX0 U64 ( .INP(in2[22]), .ZN(n21) );
  INVX0 U65 ( .INP(in1[1]), .ZN(n22) );
  INVX0 U66 ( .INP(in1[2]), .ZN(n111) );
  INVX0 U67 ( .INP(n138), .ZN(n140) );
  NOR2X0 U68 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n25) );
  AOI21X1 U69 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n25), .QN(n27) );
  NOR2X0 U70 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U71 ( .IN1(n24), .IN2(in2[0]), .IN3(n138), .IN4(n27), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U72 ( .INP(n133), .ZN(n67) );
  NOR2X0 U73 ( .IN1(n67), .IN2(n6), .QN(n28) );
  OA21X1 U74 ( .IN1(n25), .IN2(n6), .IN3(n30), .Q(n29) );
  AO22X1 U75 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n29), .Q(n26) );
  AOI22X1 U76 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n29), .QN(n32) );
  NOR2X0 U77 ( .IN1(in2[3]), .IN2(n30), .QN(n33) );
  AO21X1 U78 ( .IN1(in2[3]), .IN2(n30), .IN3(n33), .Q(n34) );
  OA22X1 U79 ( .IN1(n6), .IN2(n130), .IN3(n140), .IN4(n34), .Q(n31) );
  OA21X1 U80 ( .IN1(n33), .IN2(n7), .IN3(n37), .Q(n38) );
  AOI22X1 U81 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n38), .QN(n36) );
  OA22X1 U82 ( .IN1(n67), .IN2(n7), .IN3(n141), .IN4(n34), .Q(n35) );
  NOR2X0 U83 ( .IN1(in2[5]), .IN2(n37), .QN(n41) );
  AO21X1 U84 ( .IN1(in2[5]), .IN2(n37), .IN3(n41), .Q(n42) );
  OA22X1 U85 ( .IN1(n7), .IN2(n130), .IN3(n140), .IN4(n42), .Q(n40) );
  AOI22X1 U86 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n38), .QN(n39) );
  OA21X1 U87 ( .IN1(n41), .IN2(n8), .IN3(n45), .Q(n46) );
  AOI22X1 U88 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n46), .QN(n44) );
  OA22X1 U89 ( .IN1(n67), .IN2(n8), .IN3(n141), .IN4(n42), .Q(n43) );
  NOR2X0 U90 ( .IN1(in2[7]), .IN2(n45), .QN(n49) );
  AO21X1 U91 ( .IN1(in2[7]), .IN2(n45), .IN3(n49), .Q(n50) );
  OA22X1 U92 ( .IN1(n8), .IN2(n130), .IN3(n140), .IN4(n50), .Q(n48) );
  AOI22X1 U93 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n46), .QN(n47) );
  OA21X1 U94 ( .IN1(n49), .IN2(n9), .IN3(n53), .Q(n54) );
  AOI22X1 U95 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n54), .QN(n52) );
  OA22X1 U96 ( .IN1(n67), .IN2(n9), .IN3(n141), .IN4(n50), .Q(n51) );
  NOR2X0 U97 ( .IN1(in2[9]), .IN2(n53), .QN(n57) );
  AO21X1 U98 ( .IN1(in2[9]), .IN2(n53), .IN3(n57), .Q(n58) );
  OA22X1 U99 ( .IN1(n9), .IN2(n130), .IN3(n140), .IN4(n58), .Q(n56) );
  AOI22X1 U100 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n54), .QN(n55) );
  OA21X1 U101 ( .IN1(n57), .IN2(n10), .IN3(n61), .Q(n62) );
  AOI22X1 U102 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n62), .QN(n60) );
  OA22X1 U103 ( .IN1(n67), .IN2(n10), .IN3(n141), .IN4(n58), .Q(n59) );
  NOR2X0 U104 ( .IN1(in2[11]), .IN2(n61), .QN(n65) );
  AO21X1 U105 ( .IN1(in2[11]), .IN2(n61), .IN3(n65), .Q(n66) );
  OA22X1 U106 ( .IN1(n10), .IN2(n130), .IN3(n140), .IN4(n66), .Q(n64) );
  AOI22X1 U107 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n62), .QN(n63) );
  OA21X1 U108 ( .IN1(n65), .IN2(n11), .IN3(n77), .Q(n70) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n70), .QN(n69) );
  OA22X1 U110 ( .IN1(n67), .IN2(n11), .IN3(n141), .IN4(n66), .Q(n68) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n12), .S(n71), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n11), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n13), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n12), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n12), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n14), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n13), .IN4(n85), .IN5(n84), 
        .Q(out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n15), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n14), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n14), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n16), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n15), .IN4(n97), .IN5(n96), 
        .Q(out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n17), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n16), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n16), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n18), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n17), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n19), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n18), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n18), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n20), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n19), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n21), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n20), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n20), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n21), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_9 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n25), .IN2(n6), .QN(n30) );
  NAND2X0 U4 ( .IN1(n33), .IN2(n7), .QN(n37) );
  NAND2X0 U5 ( .IN1(n41), .IN2(n8), .QN(n45) );
  NAND2X0 U6 ( .IN1(n57), .IN2(n10), .QN(n61) );
  NAND2X0 U7 ( .IN1(n49), .IN2(n9), .QN(n53) );
  NAND2X0 U8 ( .IN1(n65), .IN2(n11), .QN(n77) );
  NAND2X0 U9 ( .IN1(n81), .IN2(n13), .QN(n89) );
  NAND2X0 U10 ( .IN1(n93), .IN2(n15), .QN(n101) );
  NAND2X0 U11 ( .IN1(n105), .IN2(n17), .QN(n114) );
  NAND2X0 U12 ( .IN1(n118), .IN2(n19), .QN(n125) );
  NAND2X0 U13 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U14 ( .IN1(in1[2]), .IN2(n77), .QN(n71) );
  NAND2X0 U15 ( .IN1(n70), .IN2(n132), .QN(n74) );
  NAND2X0 U16 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U17 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U18 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U19 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U20 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U21 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U22 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U23 ( .IN1(n141), .IN2(n130), .QN(n24) );
  NAND2X0 U24 ( .IN1(n27), .IN2(n132), .QN(n4) );
  NAND2X0 U25 ( .IN1(n64), .IN2(n63), .QN(out1[11]) );
  NAND2X0 U26 ( .IN1(n69), .IN2(n68), .QN(out1[12]) );
  NAND2X0 U27 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U28 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U29 ( .IN1(n23), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U30 ( .IN1(in1[2]), .IN2(n22), .QN(n23) );
  NAND2X0 U31 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NAND2X0 U32 ( .IN1(n32), .IN2(n31), .QN(out1[3]) );
  NAND2X0 U33 ( .IN1(n36), .IN2(n35), .QN(out1[4]) );
  NAND2X0 U34 ( .IN1(n40), .IN2(n39), .QN(out1[5]) );
  NAND2X0 U35 ( .IN1(n44), .IN2(n43), .QN(out1[6]) );
  NAND2X0 U36 ( .IN1(n48), .IN2(n47), .QN(out1[7]) );
  NAND2X0 U37 ( .IN1(n52), .IN2(n51), .QN(out1[8]) );
  NAND2X0 U38 ( .IN1(n56), .IN2(n55), .QN(out1[9]) );
  NAND2X0 U39 ( .IN1(n60), .IN2(n59), .QN(out1[10]) );
  NOR2X0 U40 ( .IN1(n28), .IN2(n26), .QN(n3) );
  NOR2X0 U41 ( .IN1(n142), .IN2(n21), .QN(n1) );
  INVX0 U42 ( .INP(n132), .ZN(n141) );
  INVX0 U43 ( .INP(n130), .ZN(n137) );
  NAND3X0 U44 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  NOR3X0 U45 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  NOR2X0 U46 ( .IN1(n142), .IN2(n111), .QN(n138) );
  MUX21X1 U47 ( .IN1(n22), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  INVX0 U48 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U49 ( .INP(in2[2]), .ZN(n6) );
  INVX0 U50 ( .INP(in2[4]), .ZN(n7) );
  INVX0 U51 ( .INP(in2[6]), .ZN(n8) );
  INVX0 U52 ( .INP(in2[8]), .ZN(n9) );
  INVX0 U53 ( .INP(in2[10]), .ZN(n10) );
  INVX0 U54 ( .INP(in2[12]), .ZN(n11) );
  INVX0 U55 ( .INP(in2[13]), .ZN(n12) );
  INVX0 U56 ( .INP(in2[14]), .ZN(n13) );
  INVX0 U57 ( .INP(in2[15]), .ZN(n14) );
  INVX0 U58 ( .INP(in2[16]), .ZN(n15) );
  INVX0 U59 ( .INP(in2[17]), .ZN(n16) );
  INVX0 U60 ( .INP(in2[18]), .ZN(n17) );
  INVX0 U61 ( .INP(in2[19]), .ZN(n18) );
  INVX0 U62 ( .INP(in2[20]), .ZN(n19) );
  INVX0 U63 ( .INP(in2[21]), .ZN(n20) );
  INVX0 U64 ( .INP(in2[22]), .ZN(n21) );
  INVX0 U65 ( .INP(in1[1]), .ZN(n22) );
  INVX0 U66 ( .INP(in1[2]), .ZN(n111) );
  INVX0 U67 ( .INP(n138), .ZN(n140) );
  NOR2X0 U68 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n25) );
  AOI21X1 U69 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n25), .QN(n27) );
  NOR2X0 U70 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U71 ( .IN1(n24), .IN2(in2[0]), .IN3(n138), .IN4(n27), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U72 ( .INP(n133), .ZN(n67) );
  NOR2X0 U73 ( .IN1(n67), .IN2(n6), .QN(n28) );
  OA21X1 U74 ( .IN1(n25), .IN2(n6), .IN3(n30), .Q(n29) );
  AO22X1 U75 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n29), .Q(n26) );
  AOI22X1 U76 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n29), .QN(n32) );
  NOR2X0 U77 ( .IN1(in2[3]), .IN2(n30), .QN(n33) );
  AO21X1 U78 ( .IN1(in2[3]), .IN2(n30), .IN3(n33), .Q(n34) );
  OA22X1 U79 ( .IN1(n6), .IN2(n130), .IN3(n140), .IN4(n34), .Q(n31) );
  OA21X1 U80 ( .IN1(n33), .IN2(n7), .IN3(n37), .Q(n38) );
  AOI22X1 U81 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n38), .QN(n36) );
  OA22X1 U82 ( .IN1(n67), .IN2(n7), .IN3(n141), .IN4(n34), .Q(n35) );
  NOR2X0 U83 ( .IN1(in2[5]), .IN2(n37), .QN(n41) );
  AO21X1 U84 ( .IN1(in2[5]), .IN2(n37), .IN3(n41), .Q(n42) );
  OA22X1 U85 ( .IN1(n7), .IN2(n130), .IN3(n140), .IN4(n42), .Q(n40) );
  AOI22X1 U86 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n38), .QN(n39) );
  OA21X1 U87 ( .IN1(n41), .IN2(n8), .IN3(n45), .Q(n46) );
  AOI22X1 U88 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n46), .QN(n44) );
  OA22X1 U89 ( .IN1(n67), .IN2(n8), .IN3(n141), .IN4(n42), .Q(n43) );
  NOR2X0 U90 ( .IN1(in2[7]), .IN2(n45), .QN(n49) );
  AO21X1 U91 ( .IN1(in2[7]), .IN2(n45), .IN3(n49), .Q(n50) );
  OA22X1 U92 ( .IN1(n8), .IN2(n130), .IN3(n140), .IN4(n50), .Q(n48) );
  AOI22X1 U93 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n46), .QN(n47) );
  OA21X1 U94 ( .IN1(n49), .IN2(n9), .IN3(n53), .Q(n54) );
  AOI22X1 U95 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n54), .QN(n52) );
  OA22X1 U96 ( .IN1(n67), .IN2(n9), .IN3(n141), .IN4(n50), .Q(n51) );
  NOR2X0 U97 ( .IN1(in2[9]), .IN2(n53), .QN(n57) );
  AO21X1 U98 ( .IN1(in2[9]), .IN2(n53), .IN3(n57), .Q(n58) );
  OA22X1 U99 ( .IN1(n9), .IN2(n130), .IN3(n140), .IN4(n58), .Q(n56) );
  AOI22X1 U100 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n54), .QN(n55) );
  OA21X1 U101 ( .IN1(n57), .IN2(n10), .IN3(n61), .Q(n62) );
  AOI22X1 U102 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n62), .QN(n60) );
  OA22X1 U103 ( .IN1(n67), .IN2(n10), .IN3(n141), .IN4(n58), .Q(n59) );
  NOR2X0 U104 ( .IN1(in2[11]), .IN2(n61), .QN(n65) );
  AO21X1 U105 ( .IN1(in2[11]), .IN2(n61), .IN3(n65), .Q(n66) );
  OA22X1 U106 ( .IN1(n10), .IN2(n130), .IN3(n140), .IN4(n66), .Q(n64) );
  AOI22X1 U107 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n62), .QN(n63) );
  OA21X1 U108 ( .IN1(n65), .IN2(n11), .IN3(n77), .Q(n70) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n70), .QN(n69) );
  OA22X1 U110 ( .IN1(n67), .IN2(n11), .IN3(n141), .IN4(n66), .Q(n68) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n12), .S(n71), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n11), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n13), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n12), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n12), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n14), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n13), .IN4(n85), .IN5(n84), 
        .Q(out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n15), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n14), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n14), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n16), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n15), .IN4(n97), .IN5(n96), 
        .Q(out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n17), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n16), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n16), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n18), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n17), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n19), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n18), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n18), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n20), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n19), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n21), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n20), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n20), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n21), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_10 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n25), .IN2(n6), .QN(n30) );
  NAND2X0 U4 ( .IN1(n33), .IN2(n7), .QN(n37) );
  NAND2X0 U5 ( .IN1(n41), .IN2(n8), .QN(n45) );
  NAND2X0 U6 ( .IN1(n49), .IN2(n9), .QN(n53) );
  NAND2X0 U7 ( .IN1(n57), .IN2(n10), .QN(n61) );
  NAND2X0 U8 ( .IN1(n65), .IN2(n11), .QN(n77) );
  NAND2X0 U9 ( .IN1(n81), .IN2(n13), .QN(n89) );
  NAND2X0 U10 ( .IN1(n93), .IN2(n15), .QN(n101) );
  NAND2X0 U11 ( .IN1(n105), .IN2(n17), .QN(n114) );
  NAND2X0 U12 ( .IN1(n118), .IN2(n19), .QN(n125) );
  NAND2X0 U13 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U14 ( .IN1(in1[2]), .IN2(n77), .QN(n71) );
  NAND2X0 U15 ( .IN1(n70), .IN2(n132), .QN(n74) );
  NAND2X0 U16 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U17 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U18 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U19 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U20 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U21 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U22 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U23 ( .IN1(n23), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U24 ( .IN1(in1[2]), .IN2(n22), .QN(n23) );
  NAND2X0 U25 ( .IN1(n32), .IN2(n31), .QN(out1[3]) );
  NAND2X0 U26 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U27 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U28 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NAND2X0 U29 ( .IN1(n27), .IN2(n132), .QN(n4) );
  NAND2X0 U30 ( .IN1(n36), .IN2(n35), .QN(out1[4]) );
  NAND2X0 U31 ( .IN1(n40), .IN2(n39), .QN(out1[5]) );
  NAND2X0 U32 ( .IN1(n44), .IN2(n43), .QN(out1[6]) );
  NAND2X0 U33 ( .IN1(n48), .IN2(n47), .QN(out1[7]) );
  NAND2X0 U34 ( .IN1(n52), .IN2(n51), .QN(out1[8]) );
  NAND2X0 U35 ( .IN1(n56), .IN2(n55), .QN(out1[9]) );
  NAND2X0 U36 ( .IN1(n60), .IN2(n59), .QN(out1[10]) );
  NAND2X0 U37 ( .IN1(n64), .IN2(n63), .QN(out1[11]) );
  NAND2X0 U38 ( .IN1(n69), .IN2(n68), .QN(out1[12]) );
  NAND2X0 U39 ( .IN1(n141), .IN2(n130), .QN(n24) );
  NOR2X0 U40 ( .IN1(n28), .IN2(n26), .QN(n3) );
  NOR2X0 U41 ( .IN1(n142), .IN2(n21), .QN(n1) );
  INVX0 U42 ( .INP(n132), .ZN(n141) );
  INVX0 U43 ( .INP(n130), .ZN(n137) );
  NAND3X0 U44 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  NOR3X0 U45 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  NOR2X0 U46 ( .IN1(n142), .IN2(n111), .QN(n138) );
  MUX21X1 U47 ( .IN1(n22), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  INVX0 U48 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U49 ( .INP(in2[2]), .ZN(n6) );
  INVX0 U50 ( .INP(in2[4]), .ZN(n7) );
  INVX0 U51 ( .INP(in2[6]), .ZN(n8) );
  INVX0 U52 ( .INP(in2[8]), .ZN(n9) );
  INVX0 U53 ( .INP(in2[10]), .ZN(n10) );
  INVX0 U54 ( .INP(in2[12]), .ZN(n11) );
  INVX0 U55 ( .INP(in2[13]), .ZN(n12) );
  INVX0 U56 ( .INP(in2[14]), .ZN(n13) );
  INVX0 U57 ( .INP(in2[15]), .ZN(n14) );
  INVX0 U58 ( .INP(in2[16]), .ZN(n15) );
  INVX0 U59 ( .INP(in2[17]), .ZN(n16) );
  INVX0 U60 ( .INP(in2[18]), .ZN(n17) );
  INVX0 U61 ( .INP(in2[19]), .ZN(n18) );
  INVX0 U62 ( .INP(in2[20]), .ZN(n19) );
  INVX0 U63 ( .INP(in2[21]), .ZN(n20) );
  INVX0 U64 ( .INP(in2[22]), .ZN(n21) );
  INVX0 U65 ( .INP(in1[1]), .ZN(n22) );
  INVX0 U66 ( .INP(in1[2]), .ZN(n111) );
  INVX0 U67 ( .INP(n138), .ZN(n140) );
  NOR2X0 U68 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n25) );
  AOI21X1 U69 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n25), .QN(n27) );
  NOR2X0 U70 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U71 ( .IN1(n24), .IN2(in2[0]), .IN3(n138), .IN4(n27), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U72 ( .INP(n133), .ZN(n67) );
  NOR2X0 U73 ( .IN1(n67), .IN2(n6), .QN(n28) );
  OA21X1 U74 ( .IN1(n25), .IN2(n6), .IN3(n30), .Q(n29) );
  AO22X1 U75 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n29), .Q(n26) );
  AOI22X1 U76 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n29), .QN(n32) );
  NOR2X0 U77 ( .IN1(in2[3]), .IN2(n30), .QN(n33) );
  AO21X1 U78 ( .IN1(in2[3]), .IN2(n30), .IN3(n33), .Q(n34) );
  OA22X1 U79 ( .IN1(n6), .IN2(n130), .IN3(n140), .IN4(n34), .Q(n31) );
  OA21X1 U80 ( .IN1(n33), .IN2(n7), .IN3(n37), .Q(n38) );
  AOI22X1 U81 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n38), .QN(n36) );
  OA22X1 U82 ( .IN1(n67), .IN2(n7), .IN3(n141), .IN4(n34), .Q(n35) );
  NOR2X0 U83 ( .IN1(in2[5]), .IN2(n37), .QN(n41) );
  AO21X1 U84 ( .IN1(in2[5]), .IN2(n37), .IN3(n41), .Q(n42) );
  OA22X1 U85 ( .IN1(n7), .IN2(n130), .IN3(n140), .IN4(n42), .Q(n40) );
  AOI22X1 U86 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n38), .QN(n39) );
  OA21X1 U87 ( .IN1(n41), .IN2(n8), .IN3(n45), .Q(n46) );
  AOI22X1 U88 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n46), .QN(n44) );
  OA22X1 U89 ( .IN1(n67), .IN2(n8), .IN3(n141), .IN4(n42), .Q(n43) );
  NOR2X0 U90 ( .IN1(in2[7]), .IN2(n45), .QN(n49) );
  AO21X1 U91 ( .IN1(in2[7]), .IN2(n45), .IN3(n49), .Q(n50) );
  OA22X1 U92 ( .IN1(n8), .IN2(n130), .IN3(n140), .IN4(n50), .Q(n48) );
  AOI22X1 U93 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n46), .QN(n47) );
  OA21X1 U94 ( .IN1(n49), .IN2(n9), .IN3(n53), .Q(n54) );
  AOI22X1 U95 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n54), .QN(n52) );
  OA22X1 U96 ( .IN1(n67), .IN2(n9), .IN3(n141), .IN4(n50), .Q(n51) );
  NOR2X0 U97 ( .IN1(in2[9]), .IN2(n53), .QN(n57) );
  AO21X1 U98 ( .IN1(in2[9]), .IN2(n53), .IN3(n57), .Q(n58) );
  OA22X1 U99 ( .IN1(n9), .IN2(n130), .IN3(n140), .IN4(n58), .Q(n56) );
  AOI22X1 U100 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n54), .QN(n55) );
  OA21X1 U101 ( .IN1(n57), .IN2(n10), .IN3(n61), .Q(n62) );
  AOI22X1 U102 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n62), .QN(n60) );
  OA22X1 U103 ( .IN1(n67), .IN2(n10), .IN3(n141), .IN4(n58), .Q(n59) );
  NOR2X0 U104 ( .IN1(in2[11]), .IN2(n61), .QN(n65) );
  AO21X1 U105 ( .IN1(in2[11]), .IN2(n61), .IN3(n65), .Q(n66) );
  OA22X1 U106 ( .IN1(n10), .IN2(n130), .IN3(n140), .IN4(n66), .Q(n64) );
  AOI22X1 U107 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n62), .QN(n63) );
  OA21X1 U108 ( .IN1(n65), .IN2(n11), .IN3(n77), .Q(n70) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n70), .QN(n69) );
  OA22X1 U110 ( .IN1(n67), .IN2(n11), .IN3(n141), .IN4(n66), .Q(n68) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n12), .S(n71), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n11), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n13), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n12), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n12), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n14), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n13), .IN4(n85), .IN5(n84), 
        .Q(out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n15), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n14), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n14), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n16), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n15), .IN4(n97), .IN5(n96), 
        .Q(out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n17), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n16), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n16), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n18), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n17), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n19), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n18), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n18), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n20), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n19), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n21), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n20), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n20), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n21), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_11 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n25), .IN2(n6), .QN(n30) );
  NAND2X0 U4 ( .IN1(n33), .IN2(n7), .QN(n37) );
  NAND2X0 U5 ( .IN1(n41), .IN2(n8), .QN(n45) );
  NAND2X0 U6 ( .IN1(n49), .IN2(n9), .QN(n53) );
  NAND2X0 U7 ( .IN1(n57), .IN2(n10), .QN(n61) );
  NAND2X0 U8 ( .IN1(n118), .IN2(n19), .QN(n125) );
  NAND2X0 U9 ( .IN1(n65), .IN2(n11), .QN(n77) );
  NAND2X0 U10 ( .IN1(n81), .IN2(n13), .QN(n89) );
  NAND2X0 U11 ( .IN1(n105), .IN2(n17), .QN(n114) );
  NAND2X0 U12 ( .IN1(n93), .IN2(n15), .QN(n101) );
  NAND2X0 U13 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U14 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U15 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U16 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U17 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U18 ( .IN1(n27), .IN2(n132), .QN(n4) );
  NAND2X0 U19 ( .IN1(n141), .IN2(n130), .QN(n24) );
  NAND2X0 U20 ( .IN1(n32), .IN2(n31), .QN(out1[3]) );
  NAND2X0 U21 ( .IN1(n36), .IN2(n35), .QN(out1[4]) );
  NAND2X0 U22 ( .IN1(in1[2]), .IN2(n77), .QN(n71) );
  NAND2X0 U23 ( .IN1(n70), .IN2(n132), .QN(n74) );
  NAND2X0 U24 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U25 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U26 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U27 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U28 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NAND2X0 U29 ( .IN1(n40), .IN2(n39), .QN(out1[5]) );
  NAND2X0 U30 ( .IN1(n44), .IN2(n43), .QN(out1[6]) );
  NAND2X0 U31 ( .IN1(n48), .IN2(n47), .QN(out1[7]) );
  NAND2X0 U32 ( .IN1(n52), .IN2(n51), .QN(out1[8]) );
  NAND2X0 U33 ( .IN1(n56), .IN2(n55), .QN(out1[9]) );
  NAND2X0 U34 ( .IN1(n60), .IN2(n59), .QN(out1[10]) );
  NAND2X0 U35 ( .IN1(n64), .IN2(n63), .QN(out1[11]) );
  NAND2X0 U36 ( .IN1(n69), .IN2(n68), .QN(out1[12]) );
  NAND2X0 U37 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U38 ( .IN1(n23), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U39 ( .IN1(in1[2]), .IN2(n22), .QN(n23) );
  INVX0 U40 ( .INP(in1[2]), .ZN(n111) );
  NOR2X0 U41 ( .IN1(n28), .IN2(n26), .QN(n3) );
  INVX0 U42 ( .INP(n130), .ZN(n137) );
  INVX0 U43 ( .INP(n132), .ZN(n141) );
  NOR3X0 U44 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  NAND3X0 U45 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  NOR2X0 U46 ( .IN1(n142), .IN2(n21), .QN(n1) );
  NOR2X0 U47 ( .IN1(n142), .IN2(n111), .QN(n138) );
  MUX21X1 U48 ( .IN1(n22), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  INVX0 U49 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U50 ( .INP(in2[2]), .ZN(n6) );
  INVX0 U51 ( .INP(in2[4]), .ZN(n7) );
  INVX0 U52 ( .INP(in2[6]), .ZN(n8) );
  INVX0 U53 ( .INP(in2[8]), .ZN(n9) );
  INVX0 U54 ( .INP(in2[10]), .ZN(n10) );
  INVX0 U55 ( .INP(in2[12]), .ZN(n11) );
  INVX0 U56 ( .INP(in2[13]), .ZN(n12) );
  INVX0 U57 ( .INP(in2[14]), .ZN(n13) );
  INVX0 U58 ( .INP(in2[15]), .ZN(n14) );
  INVX0 U59 ( .INP(in2[16]), .ZN(n15) );
  INVX0 U60 ( .INP(in2[17]), .ZN(n16) );
  INVX0 U61 ( .INP(in2[18]), .ZN(n17) );
  INVX0 U62 ( .INP(in2[19]), .ZN(n18) );
  INVX0 U63 ( .INP(in2[20]), .ZN(n19) );
  INVX0 U64 ( .INP(in2[21]), .ZN(n20) );
  INVX0 U65 ( .INP(in2[22]), .ZN(n21) );
  INVX0 U66 ( .INP(in1[1]), .ZN(n22) );
  INVX0 U67 ( .INP(n138), .ZN(n140) );
  NOR2X0 U68 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n25) );
  AOI21X1 U69 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n25), .QN(n27) );
  NOR2X0 U70 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U71 ( .IN1(n24), .IN2(in2[0]), .IN3(n138), .IN4(n27), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U72 ( .INP(n133), .ZN(n67) );
  NOR2X0 U73 ( .IN1(n67), .IN2(n6), .QN(n28) );
  OA21X1 U74 ( .IN1(n25), .IN2(n6), .IN3(n30), .Q(n29) );
  AO22X1 U75 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n29), .Q(n26) );
  AOI22X1 U76 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n29), .QN(n32) );
  NOR2X0 U77 ( .IN1(in2[3]), .IN2(n30), .QN(n33) );
  AO21X1 U78 ( .IN1(in2[3]), .IN2(n30), .IN3(n33), .Q(n34) );
  OA22X1 U79 ( .IN1(n6), .IN2(n130), .IN3(n140), .IN4(n34), .Q(n31) );
  OA21X1 U80 ( .IN1(n33), .IN2(n7), .IN3(n37), .Q(n38) );
  AOI22X1 U81 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n38), .QN(n36) );
  OA22X1 U82 ( .IN1(n67), .IN2(n7), .IN3(n141), .IN4(n34), .Q(n35) );
  NOR2X0 U83 ( .IN1(in2[5]), .IN2(n37), .QN(n41) );
  AO21X1 U84 ( .IN1(in2[5]), .IN2(n37), .IN3(n41), .Q(n42) );
  OA22X1 U85 ( .IN1(n7), .IN2(n130), .IN3(n140), .IN4(n42), .Q(n40) );
  AOI22X1 U86 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n38), .QN(n39) );
  OA21X1 U87 ( .IN1(n41), .IN2(n8), .IN3(n45), .Q(n46) );
  AOI22X1 U88 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n46), .QN(n44) );
  OA22X1 U89 ( .IN1(n67), .IN2(n8), .IN3(n141), .IN4(n42), .Q(n43) );
  NOR2X0 U90 ( .IN1(in2[7]), .IN2(n45), .QN(n49) );
  AO21X1 U91 ( .IN1(in2[7]), .IN2(n45), .IN3(n49), .Q(n50) );
  OA22X1 U92 ( .IN1(n8), .IN2(n130), .IN3(n140), .IN4(n50), .Q(n48) );
  AOI22X1 U93 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n46), .QN(n47) );
  OA21X1 U94 ( .IN1(n49), .IN2(n9), .IN3(n53), .Q(n54) );
  AOI22X1 U95 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n54), .QN(n52) );
  OA22X1 U96 ( .IN1(n67), .IN2(n9), .IN3(n141), .IN4(n50), .Q(n51) );
  NOR2X0 U97 ( .IN1(in2[9]), .IN2(n53), .QN(n57) );
  AO21X1 U98 ( .IN1(in2[9]), .IN2(n53), .IN3(n57), .Q(n58) );
  OA22X1 U99 ( .IN1(n9), .IN2(n130), .IN3(n140), .IN4(n58), .Q(n56) );
  AOI22X1 U100 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n54), .QN(n55) );
  OA21X1 U101 ( .IN1(n57), .IN2(n10), .IN3(n61), .Q(n62) );
  AOI22X1 U102 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n62), .QN(n60) );
  OA22X1 U103 ( .IN1(n67), .IN2(n10), .IN3(n141), .IN4(n58), .Q(n59) );
  NOR2X0 U104 ( .IN1(in2[11]), .IN2(n61), .QN(n65) );
  AO21X1 U105 ( .IN1(in2[11]), .IN2(n61), .IN3(n65), .Q(n66) );
  OA22X1 U106 ( .IN1(n10), .IN2(n130), .IN3(n140), .IN4(n66), .Q(n64) );
  AOI22X1 U107 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n62), .QN(n63) );
  OA21X1 U108 ( .IN1(n65), .IN2(n11), .IN3(n77), .Q(n70) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n70), .QN(n69) );
  OA22X1 U110 ( .IN1(n67), .IN2(n11), .IN3(n141), .IN4(n66), .Q(n68) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n12), .S(n71), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n11), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n13), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n12), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n12), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n14), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n13), .IN4(n85), .IN5(n84), 
        .Q(out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n15), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n14), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n14), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n16), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n15), .IN4(n97), .IN5(n96), 
        .Q(out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n17), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n16), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n16), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n18), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n17), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n19), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n18), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n18), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n20), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n19), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n21), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n20), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n20), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n21), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_12 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n33), .IN2(n7), .QN(n37) );
  NAND2X0 U4 ( .IN1(n41), .IN2(n8), .QN(n45) );
  NAND2X0 U5 ( .IN1(n49), .IN2(n9), .QN(n53) );
  NAND2X0 U6 ( .IN1(n57), .IN2(n10), .QN(n61) );
  NAND2X0 U7 ( .IN1(n25), .IN2(n6), .QN(n30) );
  NAND2X0 U8 ( .IN1(n65), .IN2(n11), .QN(n77) );
  NAND2X0 U9 ( .IN1(n81), .IN2(n13), .QN(n89) );
  NAND2X0 U10 ( .IN1(n93), .IN2(n15), .QN(n101) );
  NAND2X0 U11 ( .IN1(n118), .IN2(n19), .QN(n125) );
  NAND2X0 U12 ( .IN1(n105), .IN2(n17), .QN(n114) );
  NAND2X0 U13 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U14 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U15 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U16 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U17 ( .IN1(n40), .IN2(n39), .QN(out1[5]) );
  NAND2X0 U18 ( .IN1(n44), .IN2(n43), .QN(out1[6]) );
  NAND2X0 U19 ( .IN1(in1[2]), .IN2(n77), .QN(n71) );
  NAND2X0 U20 ( .IN1(n70), .IN2(n132), .QN(n74) );
  NAND2X0 U21 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U22 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U23 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U24 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U25 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U26 ( .IN1(n23), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U27 ( .IN1(in1[2]), .IN2(n22), .QN(n23) );
  NAND2X0 U28 ( .IN1(n36), .IN2(n35), .QN(out1[4]) );
  NAND2X0 U29 ( .IN1(n32), .IN2(n31), .QN(out1[3]) );
  NAND2X0 U30 ( .IN1(n27), .IN2(n132), .QN(n4) );
  NAND2X0 U31 ( .IN1(n48), .IN2(n47), .QN(out1[7]) );
  NAND2X0 U32 ( .IN1(n52), .IN2(n51), .QN(out1[8]) );
  NAND2X0 U33 ( .IN1(n56), .IN2(n55), .QN(out1[9]) );
  NAND2X0 U34 ( .IN1(n60), .IN2(n59), .QN(out1[10]) );
  NAND2X0 U35 ( .IN1(n64), .IN2(n63), .QN(out1[11]) );
  NAND2X0 U36 ( .IN1(n69), .IN2(n68), .QN(out1[12]) );
  NAND2X0 U37 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U38 ( .IN1(n141), .IN2(n130), .QN(n24) );
  NAND2X0 U39 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NOR2X0 U40 ( .IN1(n28), .IN2(n26), .QN(n3) );
  NOR2X0 U41 ( .IN1(n142), .IN2(n21), .QN(n1) );
  INVX0 U42 ( .INP(n132), .ZN(n141) );
  INVX0 U43 ( .INP(n130), .ZN(n137) );
  NAND3X0 U44 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  NOR2X0 U45 ( .IN1(n142), .IN2(n111), .QN(n138) );
  MUX21X1 U46 ( .IN1(n22), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  NOR3X0 U47 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  INVX0 U48 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U49 ( .INP(in2[2]), .ZN(n6) );
  INVX0 U50 ( .INP(in2[4]), .ZN(n7) );
  INVX0 U51 ( .INP(in2[6]), .ZN(n8) );
  INVX0 U52 ( .INP(in2[8]), .ZN(n9) );
  INVX0 U53 ( .INP(in2[10]), .ZN(n10) );
  INVX0 U54 ( .INP(in2[12]), .ZN(n11) );
  INVX0 U55 ( .INP(in2[13]), .ZN(n12) );
  INVX0 U56 ( .INP(in2[14]), .ZN(n13) );
  INVX0 U57 ( .INP(in2[15]), .ZN(n14) );
  INVX0 U58 ( .INP(in2[16]), .ZN(n15) );
  INVX0 U59 ( .INP(in2[17]), .ZN(n16) );
  INVX0 U60 ( .INP(in2[18]), .ZN(n17) );
  INVX0 U61 ( .INP(in2[19]), .ZN(n18) );
  INVX0 U62 ( .INP(in2[20]), .ZN(n19) );
  INVX0 U63 ( .INP(in2[21]), .ZN(n20) );
  INVX0 U64 ( .INP(in2[22]), .ZN(n21) );
  INVX0 U65 ( .INP(in1[1]), .ZN(n22) );
  INVX0 U66 ( .INP(in1[2]), .ZN(n111) );
  INVX0 U67 ( .INP(n138), .ZN(n140) );
  NOR2X0 U68 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n25) );
  AOI21X1 U69 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n25), .QN(n27) );
  NOR2X0 U70 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U71 ( .IN1(n24), .IN2(in2[0]), .IN3(n138), .IN4(n27), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U72 ( .INP(n133), .ZN(n67) );
  NOR2X0 U73 ( .IN1(n67), .IN2(n6), .QN(n28) );
  OA21X1 U74 ( .IN1(n25), .IN2(n6), .IN3(n30), .Q(n29) );
  AO22X1 U75 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n29), .Q(n26) );
  AOI22X1 U76 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n29), .QN(n32) );
  NOR2X0 U77 ( .IN1(in2[3]), .IN2(n30), .QN(n33) );
  AO21X1 U78 ( .IN1(in2[3]), .IN2(n30), .IN3(n33), .Q(n34) );
  OA22X1 U79 ( .IN1(n6), .IN2(n130), .IN3(n140), .IN4(n34), .Q(n31) );
  OA21X1 U80 ( .IN1(n33), .IN2(n7), .IN3(n37), .Q(n38) );
  AOI22X1 U81 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n38), .QN(n36) );
  OA22X1 U82 ( .IN1(n67), .IN2(n7), .IN3(n141), .IN4(n34), .Q(n35) );
  NOR2X0 U83 ( .IN1(in2[5]), .IN2(n37), .QN(n41) );
  AO21X1 U84 ( .IN1(in2[5]), .IN2(n37), .IN3(n41), .Q(n42) );
  OA22X1 U85 ( .IN1(n7), .IN2(n130), .IN3(n140), .IN4(n42), .Q(n40) );
  AOI22X1 U86 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n38), .QN(n39) );
  OA21X1 U87 ( .IN1(n41), .IN2(n8), .IN3(n45), .Q(n46) );
  AOI22X1 U88 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n46), .QN(n44) );
  OA22X1 U89 ( .IN1(n67), .IN2(n8), .IN3(n141), .IN4(n42), .Q(n43) );
  NOR2X0 U90 ( .IN1(in2[7]), .IN2(n45), .QN(n49) );
  AO21X1 U91 ( .IN1(in2[7]), .IN2(n45), .IN3(n49), .Q(n50) );
  OA22X1 U92 ( .IN1(n8), .IN2(n130), .IN3(n140), .IN4(n50), .Q(n48) );
  AOI22X1 U93 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n46), .QN(n47) );
  OA21X1 U94 ( .IN1(n49), .IN2(n9), .IN3(n53), .Q(n54) );
  AOI22X1 U95 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n54), .QN(n52) );
  OA22X1 U96 ( .IN1(n67), .IN2(n9), .IN3(n141), .IN4(n50), .Q(n51) );
  NOR2X0 U97 ( .IN1(in2[9]), .IN2(n53), .QN(n57) );
  AO21X1 U98 ( .IN1(in2[9]), .IN2(n53), .IN3(n57), .Q(n58) );
  OA22X1 U99 ( .IN1(n9), .IN2(n130), .IN3(n140), .IN4(n58), .Q(n56) );
  AOI22X1 U100 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n54), .QN(n55) );
  OA21X1 U101 ( .IN1(n57), .IN2(n10), .IN3(n61), .Q(n62) );
  AOI22X1 U102 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n62), .QN(n60) );
  OA22X1 U103 ( .IN1(n67), .IN2(n10), .IN3(n141), .IN4(n58), .Q(n59) );
  NOR2X0 U104 ( .IN1(in2[11]), .IN2(n61), .QN(n65) );
  AO21X1 U105 ( .IN1(in2[11]), .IN2(n61), .IN3(n65), .Q(n66) );
  OA22X1 U106 ( .IN1(n10), .IN2(n130), .IN3(n140), .IN4(n66), .Q(n64) );
  AOI22X1 U107 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n62), .QN(n63) );
  OA21X1 U108 ( .IN1(n65), .IN2(n11), .IN3(n77), .Q(n70) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n70), .QN(n69) );
  OA22X1 U110 ( .IN1(n67), .IN2(n11), .IN3(n141), .IN4(n66), .Q(n68) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n12), .S(n71), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n11), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n13), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n12), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n12), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n14), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n13), .IN4(n85), .IN5(n84), 
        .Q(out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n15), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n14), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n14), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n16), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n15), .IN4(n97), .IN5(n96), 
        .Q(out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n17), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n16), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n16), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n18), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n17), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n19), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n18), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n18), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n20), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n19), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n21), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n20), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n20), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n21), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_13 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93;

  NAND2X0 U3 ( .IN1(n30), .IN2(n7), .QN(n32) );
  NAND2X0 U4 ( .IN1(n34), .IN2(n8), .QN(n36) );
  NAND2X0 U5 ( .IN1(n38), .IN2(n9), .QN(n40) );
  NAND2X0 U6 ( .IN1(n42), .IN2(n10), .QN(n47) );
  NAND2X0 U7 ( .IN1(n78), .IN2(n18), .QN(n82) );
  NAND2X0 U8 ( .IN1(n26), .IN2(n6), .QN(n28) );
  NAND2X0 U9 ( .IN1(in1[2]), .IN2(n47), .QN(n44) );
  NAND2X0 U10 ( .IN1(n52), .IN2(n12), .QN(n55) );
  NAND2X0 U11 ( .IN1(in1[2]), .IN2(n55), .QN(n51) );
  NAND2X0 U12 ( .IN1(n60), .IN2(n14), .QN(n63) );
  NAND2X0 U13 ( .IN1(in1[2]), .IN2(n63), .QN(n59) );
  NAND2X0 U14 ( .IN1(n68), .IN2(n16), .QN(n71) );
  NAND2X0 U15 ( .IN1(in1[2]), .IN2(n71), .QN(n67) );
  NAND2X0 U16 ( .IN1(in1[2]), .IN2(n82), .QN(n77) );
  NAND2X0 U17 ( .IN1(in2[21]), .IN2(n82), .QN(n83) );
  NAND2X0 U18 ( .IN1(n75), .IN2(in1[2]), .QN(n86) );
  NAND2X0 U19 ( .IN1(n3), .IN2(n4), .QN(n22) );
  NAND2X0 U20 ( .IN1(in2[1]), .IN2(in2[0]), .QN(n4) );
  NAND2X0 U21 ( .IN1(n23), .IN2(n22), .QN(out1[2]) );
  INVX0 U22 ( .INP(n86), .ZN(n89) );
  NOR2X0 U23 ( .IN1(n21), .IN2(n86), .QN(n3) );
  NOR2X0 U24 ( .IN1(in1[2]), .IN2(n75), .QN(n90) );
  NBUFFX2 U25 ( .INP(in1[2]), .Z(out1[25]) );
  NOR2X0 U26 ( .IN1(n75), .IN2(n72), .QN(n92) );
  NBUFFX2 U27 ( .INP(in1[2]), .Z(out1[26]) );
  INVX0 U28 ( .INP(in2[2]), .ZN(n5) );
  INVX0 U29 ( .INP(in2[4]), .ZN(n6) );
  INVX0 U30 ( .INP(in2[6]), .ZN(n7) );
  INVX0 U31 ( .INP(in2[8]), .ZN(n8) );
  INVX0 U32 ( .INP(in2[10]), .ZN(n9) );
  INVX0 U33 ( .INP(in2[12]), .ZN(n10) );
  INVX0 U34 ( .INP(in2[13]), .ZN(n11) );
  INVX0 U35 ( .INP(in2[14]), .ZN(n12) );
  INVX0 U36 ( .INP(in2[15]), .ZN(n13) );
  INVX0 U37 ( .INP(in2[16]), .ZN(n14) );
  INVX0 U38 ( .INP(in2[17]), .ZN(n15) );
  INVX0 U39 ( .INP(in2[18]), .ZN(n16) );
  INVX0 U40 ( .INP(in2[19]), .ZN(n17) );
  INVX0 U41 ( .INP(in2[20]), .ZN(n18) );
  INVX0 U42 ( .INP(in2[21]), .ZN(n19) );
  INVX0 U43 ( .INP(in2[22]), .ZN(n20) );
  INVX0 U44 ( .INP(in1[1]), .ZN(n75) );
  INVX0 U45 ( .INP(in1[2]), .ZN(n72) );
  NOR2X0 U46 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n21) );
  OR3X1 U47 ( .IN1(in2[2]), .IN2(in2[0]), .IN3(in2[1]), .Q(n24) );
  OA21X1 U48 ( .IN1(n21), .IN2(n5), .IN3(n24), .Q(n25) );
  AOI22X1 U49 ( .IN1(in2[2]), .IN2(n90), .IN3(n92), .IN4(n25), .QN(n23) );
  NOR2X0 U50 ( .IN1(in2[3]), .IN2(n24), .QN(n26) );
  AOI21X1 U51 ( .IN1(in2[3]), .IN2(n24), .IN3(n26), .QN(n27) );
  AO222X1 U52 ( .IN1(in2[3]), .IN2(n90), .IN3(n92), .IN4(n27), .IN5(n89), 
        .IN6(n25), .Q(out1[3]) );
  OA21X1 U53 ( .IN1(n26), .IN2(n6), .IN3(n28), .Q(n29) );
  AO222X1 U54 ( .IN1(in2[4]), .IN2(n90), .IN3(n92), .IN4(n29), .IN5(n89), 
        .IN6(n27), .Q(out1[4]) );
  NOR2X0 U55 ( .IN1(in2[5]), .IN2(n28), .QN(n30) );
  AOI21X1 U56 ( .IN1(in2[5]), .IN2(n28), .IN3(n30), .QN(n31) );
  AO222X1 U57 ( .IN1(in2[5]), .IN2(n90), .IN3(n92), .IN4(n31), .IN5(n89), 
        .IN6(n29), .Q(out1[5]) );
  OA21X1 U58 ( .IN1(n30), .IN2(n7), .IN3(n32), .Q(n33) );
  AO222X1 U59 ( .IN1(in2[6]), .IN2(n90), .IN3(n92), .IN4(n33), .IN5(n89), 
        .IN6(n31), .Q(out1[6]) );
  NOR2X0 U60 ( .IN1(in2[7]), .IN2(n32), .QN(n34) );
  AOI21X1 U61 ( .IN1(in2[7]), .IN2(n32), .IN3(n34), .QN(n35) );
  AO222X1 U62 ( .IN1(in2[7]), .IN2(n90), .IN3(n92), .IN4(n35), .IN5(n89), 
        .IN6(n33), .Q(out1[7]) );
  OA21X1 U63 ( .IN1(n34), .IN2(n8), .IN3(n36), .Q(n37) );
  AO222X1 U64 ( .IN1(in2[8]), .IN2(n90), .IN3(n92), .IN4(n37), .IN5(n89), 
        .IN6(n35), .Q(out1[8]) );
  NOR2X0 U65 ( .IN1(in2[9]), .IN2(n36), .QN(n38) );
  AOI21X1 U66 ( .IN1(in2[9]), .IN2(n36), .IN3(n38), .QN(n39) );
  AO222X1 U67 ( .IN1(in2[9]), .IN2(n90), .IN3(n92), .IN4(n39), .IN5(n89), 
        .IN6(n37), .Q(out1[9]) );
  OA21X1 U68 ( .IN1(n38), .IN2(n9), .IN3(n40), .Q(n41) );
  AO222X1 U69 ( .IN1(in2[10]), .IN2(n90), .IN3(n92), .IN4(n41), .IN5(n89), 
        .IN6(n39), .Q(out1[10]) );
  NOR2X0 U70 ( .IN1(in2[11]), .IN2(n40), .QN(n42) );
  AOI21X1 U71 ( .IN1(in2[11]), .IN2(n40), .IN3(n42), .QN(n43) );
  AO222X1 U72 ( .IN1(in2[11]), .IN2(n90), .IN3(n92), .IN4(n43), .IN5(n89), 
        .IN6(n41), .Q(out1[11]) );
  OA21X1 U73 ( .IN1(n42), .IN2(n10), .IN3(n47), .Q(n45) );
  AO222X1 U74 ( .IN1(in2[12]), .IN2(n90), .IN3(n92), .IN4(n45), .IN5(n89), 
        .IN6(n43), .Q(out1[12]) );
  MUX21X1 U75 ( .IN1(n11), .IN2(in2[13]), .S(n44), .Q(n46) );
  AO22X1 U76 ( .IN1(in1[1]), .IN2(n46), .IN3(n89), .IN4(n45), .Q(out1[13]) );
  NOR2X0 U77 ( .IN1(in2[13]), .IN2(n47), .QN(n52) );
  AO21X1 U78 ( .IN1(in2[13]), .IN2(n47), .IN3(n86), .Q(n50) );
  NOR2X0 U79 ( .IN1(n52), .IN2(n72), .QN(n48) );
  MUX21X1 U80 ( .IN1(n12), .IN2(in2[14]), .S(n48), .Q(n49) );
  OAI22X1 U81 ( .IN1(n52), .IN2(n50), .IN3(n75), .IN4(n49), .QN(out1[14]) );
  MUX21X1 U82 ( .IN1(n13), .IN2(in2[15]), .S(n51), .Q(n54) );
  OA21X1 U83 ( .IN1(n52), .IN2(n12), .IN3(n89), .Q(n53) );
  AO22X1 U84 ( .IN1(in1[1]), .IN2(n54), .IN3(n53), .IN4(n55), .Q(out1[15]) );
  NOR2X0 U85 ( .IN1(in2[15]), .IN2(n55), .QN(n60) );
  AO21X1 U86 ( .IN1(in2[15]), .IN2(n55), .IN3(n86), .Q(n58) );
  NOR2X0 U87 ( .IN1(n60), .IN2(n72), .QN(n56) );
  MUX21X1 U88 ( .IN1(n14), .IN2(in2[16]), .S(n56), .Q(n57) );
  OAI22X1 U89 ( .IN1(n60), .IN2(n58), .IN3(n75), .IN4(n57), .QN(out1[16]) );
  MUX21X1 U90 ( .IN1(n15), .IN2(in2[17]), .S(n59), .Q(n62) );
  OA21X1 U91 ( .IN1(n60), .IN2(n14), .IN3(n89), .Q(n61) );
  AO22X1 U92 ( .IN1(in1[1]), .IN2(n62), .IN3(n61), .IN4(n63), .Q(out1[17]) );
  NOR2X0 U93 ( .IN1(in2[17]), .IN2(n63), .QN(n68) );
  AO21X1 U94 ( .IN1(in2[17]), .IN2(n63), .IN3(n86), .Q(n66) );
  NOR2X0 U95 ( .IN1(n68), .IN2(n72), .QN(n64) );
  MUX21X1 U96 ( .IN1(n16), .IN2(in2[18]), .S(n64), .Q(n65) );
  OAI22X1 U97 ( .IN1(n68), .IN2(n66), .IN3(n75), .IN4(n65), .QN(out1[18]) );
  MUX21X1 U98 ( .IN1(n17), .IN2(in2[19]), .S(n67), .Q(n70) );
  OA21X1 U99 ( .IN1(n68), .IN2(n16), .IN3(n89), .Q(n69) );
  AO22X1 U100 ( .IN1(in1[1]), .IN2(n70), .IN3(n69), .IN4(n71), .Q(out1[19]) );
  NOR2X0 U101 ( .IN1(in2[19]), .IN2(n71), .QN(n78) );
  AO21X1 U102 ( .IN1(in2[19]), .IN2(n71), .IN3(n86), .Q(n76) );
  NOR2X0 U103 ( .IN1(n78), .IN2(n72), .QN(n73) );
  MUX21X1 U104 ( .IN1(n18), .IN2(in2[20]), .S(n73), .Q(n74) );
  OAI22X1 U105 ( .IN1(n78), .IN2(n76), .IN3(n75), .IN4(n74), .QN(out1[20]) );
  MUX21X1 U106 ( .IN1(n19), .IN2(in2[21]), .S(n77), .Q(n80) );
  MUX21X1 U107 ( .IN1(n18), .IN2(in2[20]), .S(n78), .Q(n79) );
  AO22X1 U108 ( .IN1(in1[1]), .IN2(n80), .IN3(n89), .IN4(n79), .Q(out1[21]) );
  INVX0 U109 ( .INP(n92), .ZN(n81) );
  OR2X1 U110 ( .IN1(n82), .IN2(in2[21]), .Q(n88) );
  NOR2X0 U111 ( .IN1(n81), .IN2(n88), .QN(n87) );
  NOR2X0 U112 ( .IN1(in2[22]), .IN2(n81), .QN(n84) );
  OA221X1 U113 ( .IN1(n84), .IN2(n89), .IN3(n84), .IN4(n83), .IN5(n88), .Q(n85) );
  AO221X1 U114 ( .IN1(in2[22]), .IN2(n87), .IN3(in2[22]), .IN4(n90), .IN5(n85), 
        .Q(out1[22]) );
  NOR2X0 U115 ( .IN1(n86), .IN2(n88), .QN(n93) );
  AO21X1 U116 ( .IN1(n89), .IN2(n88), .IN3(n87), .Q(n91) );
  AO221X1 U117 ( .IN1(in2[22]), .IN2(n93), .IN3(n20), .IN4(n91), .IN5(n90), 
        .Q(out1[23]) );
  AO21X1 U118 ( .IN1(n93), .IN2(n20), .IN3(n92), .Q(out1[24]) );
endmodule


module mul26_1 ( clk, rst_n, in1, in2, en, mulout );
  input [25:0] in1;
  input [25:0] in2;
  output [50:0] mulout;
  input clk, rst_n, en;
  wire   N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24,
         N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38,
         N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N62, N63,
         N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77,
         N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91,
         N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n128,
         n129, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22,
         SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24,
         SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26,
         SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28,
         SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30,
         SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32,
         SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34,
         SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36,
         SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38,
         SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40,
         SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42,
         SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44,
         SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46,
         SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48,
         SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50,
         SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52,
         SYNOPSYS_UNCONNECTED_53, SYNOPSYS_UNCONNECTED_54,
         SYNOPSYS_UNCONNECTED_55, SYNOPSYS_UNCONNECTED_56,
         SYNOPSYS_UNCONNECTED_57, SYNOPSYS_UNCONNECTED_58,
         SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_60,
         SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_62,
         SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_64,
         SYNOPSYS_UNCONNECTED_65, SYNOPSYS_UNCONNECTED_66,
         SYNOPSYS_UNCONNECTED_67, SYNOPSYS_UNCONNECTED_68,
         SYNOPSYS_UNCONNECTED_69, SYNOPSYS_UNCONNECTED_70,
         SYNOPSYS_UNCONNECTED_71, SYNOPSYS_UNCONNECTED_72,
         SYNOPSYS_UNCONNECTED_73, SYNOPSYS_UNCONNECTED_74,
         SYNOPSYS_UNCONNECTED_75, SYNOPSYS_UNCONNECTED_76,
         SYNOPSYS_UNCONNECTED_77, SYNOPSYS_UNCONNECTED_78,
         SYNOPSYS_UNCONNECTED_79, SYNOPSYS_UNCONNECTED_80,
         SYNOPSYS_UNCONNECTED_81, SYNOPSYS_UNCONNECTED_82,
         SYNOPSYS_UNCONNECTED_83, SYNOPSYS_UNCONNECTED_84,
         SYNOPSYS_UNCONNECTED_85, SYNOPSYS_UNCONNECTED_86,
         SYNOPSYS_UNCONNECTED_87, SYNOPSYS_UNCONNECTED_88,
         SYNOPSYS_UNCONNECTED_89, SYNOPSYS_UNCONNECTED_90,
         SYNOPSYS_UNCONNECTED_91, SYNOPSYS_UNCONNECTED_92,
         SYNOPSYS_UNCONNECTED_93, SYNOPSYS_UNCONNECTED_94,
         SYNOPSYS_UNCONNECTED_95, SYNOPSYS_UNCONNECTED_96,
         SYNOPSYS_UNCONNECTED_97, SYNOPSYS_UNCONNECTED_98,
         SYNOPSYS_UNCONNECTED_99, SYNOPSYS_UNCONNECTED_100,
         SYNOPSYS_UNCONNECTED_101, SYNOPSYS_UNCONNECTED_102,
         SYNOPSYS_UNCONNECTED_103, SYNOPSYS_UNCONNECTED_104,
         SYNOPSYS_UNCONNECTED_105, SYNOPSYS_UNCONNECTED_106,
         SYNOPSYS_UNCONNECTED_107, SYNOPSYS_UNCONNECTED_108,
         SYNOPSYS_UNCONNECTED_109, SYNOPSYS_UNCONNECTED_110,
         SYNOPSYS_UNCONNECTED_111, SYNOPSYS_UNCONNECTED_112,
         SYNOPSYS_UNCONNECTED_113, SYNOPSYS_UNCONNECTED_114,
         SYNOPSYS_UNCONNECTED_115, SYNOPSYS_UNCONNECTED_116,
         SYNOPSYS_UNCONNECTED_117, SYNOPSYS_UNCONNECTED_118,
         SYNOPSYS_UNCONNECTED_119, SYNOPSYS_UNCONNECTED_120,
         SYNOPSYS_UNCONNECTED_121, SYNOPSYS_UNCONNECTED_122,
         SYNOPSYS_UNCONNECTED_123, SYNOPSYS_UNCONNECTED_124,
         SYNOPSYS_UNCONNECTED_125, SYNOPSYS_UNCONNECTED_126,
         SYNOPSYS_UNCONNECTED_127, SYNOPSYS_UNCONNECTED_128,
         SYNOPSYS_UNCONNECTED_129, SYNOPSYS_UNCONNECTED_130,
         SYNOPSYS_UNCONNECTED_131, SYNOPSYS_UNCONNECTED_132,
         SYNOPSYS_UNCONNECTED_133, SYNOPSYS_UNCONNECTED_134,
         SYNOPSYS_UNCONNECTED_135, SYNOPSYS_UNCONNECTED_136,
         SYNOPSYS_UNCONNECTED_137, SYNOPSYS_UNCONNECTED_138,
         SYNOPSYS_UNCONNECTED_139, SYNOPSYS_UNCONNECTED_140,
         SYNOPSYS_UNCONNECTED_141, SYNOPSYS_UNCONNECTED_142,
         SYNOPSYS_UNCONNECTED_143, SYNOPSYS_UNCONNECTED_144,
         SYNOPSYS_UNCONNECTED_145, SYNOPSYS_UNCONNECTED_146,
         SYNOPSYS_UNCONNECTED_147, SYNOPSYS_UNCONNECTED_148,
         SYNOPSYS_UNCONNECTED_149, SYNOPSYS_UNCONNECTED_150,
         SYNOPSYS_UNCONNECTED_151, SYNOPSYS_UNCONNECTED_152,
         SYNOPSYS_UNCONNECTED_153, SYNOPSYS_UNCONNECTED_154,
         SYNOPSYS_UNCONNECTED_155, SYNOPSYS_UNCONNECTED_156,
         SYNOPSYS_UNCONNECTED_157, SYNOPSYS_UNCONNECTED_158,
         SYNOPSYS_UNCONNECTED_159, SYNOPSYS_UNCONNECTED_160,
         SYNOPSYS_UNCONNECTED_161, SYNOPSYS_UNCONNECTED_162,
         SYNOPSYS_UNCONNECTED_163, SYNOPSYS_UNCONNECTED_164,
         SYNOPSYS_UNCONNECTED_165, SYNOPSYS_UNCONNECTED_166,
         SYNOPSYS_UNCONNECTED_167, SYNOPSYS_UNCONNECTED_168,
         SYNOPSYS_UNCONNECTED_169, SYNOPSYS_UNCONNECTED_170,
         SYNOPSYS_UNCONNECTED_171, SYNOPSYS_UNCONNECTED_172,
         SYNOPSYS_UNCONNECTED_173, SYNOPSYS_UNCONNECTED_174,
         SYNOPSYS_UNCONNECTED_175, SYNOPSYS_UNCONNECTED_176,
         SYNOPSYS_UNCONNECTED_177, SYNOPSYS_UNCONNECTED_178,
         SYNOPSYS_UNCONNECTED_179, SYNOPSYS_UNCONNECTED_180,
         SYNOPSYS_UNCONNECTED_181, SYNOPSYS_UNCONNECTED_182,
         SYNOPSYS_UNCONNECTED_183, SYNOPSYS_UNCONNECTED_184,
         SYNOPSYS_UNCONNECTED_185, SYNOPSYS_UNCONNECTED_186,
         SYNOPSYS_UNCONNECTED_187, SYNOPSYS_UNCONNECTED_188,
         SYNOPSYS_UNCONNECTED_189, SYNOPSYS_UNCONNECTED_190,
         SYNOPSYS_UNCONNECTED_191, SYNOPSYS_UNCONNECTED_192,
         SYNOPSYS_UNCONNECTED_193, SYNOPSYS_UNCONNECTED_194,
         SYNOPSYS_UNCONNECTED_195, SYNOPSYS_UNCONNECTED_196,
         SYNOPSYS_UNCONNECTED_197, SYNOPSYS_UNCONNECTED_198,
         SYNOPSYS_UNCONNECTED_199, SYNOPSYS_UNCONNECTED_200,
         SYNOPSYS_UNCONNECTED_201, SYNOPSYS_UNCONNECTED_202,
         SYNOPSYS_UNCONNECTED_203, SYNOPSYS_UNCONNECTED_204,
         SYNOPSYS_UNCONNECTED_205, SYNOPSYS_UNCONNECTED_206,
         SYNOPSYS_UNCONNECTED_207, SYNOPSYS_UNCONNECTED_208,
         SYNOPSYS_UNCONNECTED_209, SYNOPSYS_UNCONNECTED_210,
         SYNOPSYS_UNCONNECTED_211, SYNOPSYS_UNCONNECTED_212,
         SYNOPSYS_UNCONNECTED_213, SYNOPSYS_UNCONNECTED_214,
         SYNOPSYS_UNCONNECTED_215, SYNOPSYS_UNCONNECTED_216,
         SYNOPSYS_UNCONNECTED_217, SYNOPSYS_UNCONNECTED_218,
         SYNOPSYS_UNCONNECTED_219, SYNOPSYS_UNCONNECTED_220,
         SYNOPSYS_UNCONNECTED_221, SYNOPSYS_UNCONNECTED_222,
         SYNOPSYS_UNCONNECTED_223, SYNOPSYS_UNCONNECTED_224,
         SYNOPSYS_UNCONNECTED_225, SYNOPSYS_UNCONNECTED_226,
         SYNOPSYS_UNCONNECTED_227, SYNOPSYS_UNCONNECTED_228,
         SYNOPSYS_UNCONNECTED_229, SYNOPSYS_UNCONNECTED_230,
         SYNOPSYS_UNCONNECTED_231, SYNOPSYS_UNCONNECTED_232,
         SYNOPSYS_UNCONNECTED_233, SYNOPSYS_UNCONNECTED_234,
         SYNOPSYS_UNCONNECTED_235, SYNOPSYS_UNCONNECTED_236,
         SYNOPSYS_UNCONNECTED_237, SYNOPSYS_UNCONNECTED_238,
         SYNOPSYS_UNCONNECTED_239, SYNOPSYS_UNCONNECTED_240,
         SYNOPSYS_UNCONNECTED_241, SYNOPSYS_UNCONNECTED_242,
         SYNOPSYS_UNCONNECTED_243, SYNOPSYS_UNCONNECTED_244,
         SYNOPSYS_UNCONNECTED_245, SYNOPSYS_UNCONNECTED_246,
         SYNOPSYS_UNCONNECTED_247, SYNOPSYS_UNCONNECTED_248,
         SYNOPSYS_UNCONNECTED_249, SYNOPSYS_UNCONNECTED_250,
         SYNOPSYS_UNCONNECTED_251, SYNOPSYS_UNCONNECTED_252,
         SYNOPSYS_UNCONNECTED_253, SYNOPSYS_UNCONNECTED_254,
         SYNOPSYS_UNCONNECTED_255, SYNOPSYS_UNCONNECTED_256,
         SYNOPSYS_UNCONNECTED_257, SYNOPSYS_UNCONNECTED_258,
         SYNOPSYS_UNCONNECTED_259, SYNOPSYS_UNCONNECTED_260,
         SYNOPSYS_UNCONNECTED_261, SYNOPSYS_UNCONNECTED_262,
         SYNOPSYS_UNCONNECTED_263, SYNOPSYS_UNCONNECTED_264,
         SYNOPSYS_UNCONNECTED_265, SYNOPSYS_UNCONNECTED_266,
         SYNOPSYS_UNCONNECTED_267, SYNOPSYS_UNCONNECTED_268,
         SYNOPSYS_UNCONNECTED_269, SYNOPSYS_UNCONNECTED_270,
         SYNOPSYS_UNCONNECTED_271, SYNOPSYS_UNCONNECTED_272,
         SYNOPSYS_UNCONNECTED_273, SYNOPSYS_UNCONNECTED_274,
         SYNOPSYS_UNCONNECTED_275, SYNOPSYS_UNCONNECTED_276,
         SYNOPSYS_UNCONNECTED_277, SYNOPSYS_UNCONNECTED_278,
         SYNOPSYS_UNCONNECTED_279, SYNOPSYS_UNCONNECTED_280,
         SYNOPSYS_UNCONNECTED_281, SYNOPSYS_UNCONNECTED_282,
         SYNOPSYS_UNCONNECTED_283, SYNOPSYS_UNCONNECTED_284,
         SYNOPSYS_UNCONNECTED_285, SYNOPSYS_UNCONNECTED_286,
         SYNOPSYS_UNCONNECTED_287, SYNOPSYS_UNCONNECTED_288,
         SYNOPSYS_UNCONNECTED_289, SYNOPSYS_UNCONNECTED_290,
         SYNOPSYS_UNCONNECTED_291, SYNOPSYS_UNCONNECTED_292,
         SYNOPSYS_UNCONNECTED_293, SYNOPSYS_UNCONNECTED_294,
         SYNOPSYS_UNCONNECTED_295, SYNOPSYS_UNCONNECTED_296,
         SYNOPSYS_UNCONNECTED_297, SYNOPSYS_UNCONNECTED_298,
         SYNOPSYS_UNCONNECTED_299, SYNOPSYS_UNCONNECTED_300,
         SYNOPSYS_UNCONNECTED_301, SYNOPSYS_UNCONNECTED_302,
         SYNOPSYS_UNCONNECTED_303, SYNOPSYS_UNCONNECTED_304,
         SYNOPSYS_UNCONNECTED_305, SYNOPSYS_UNCONNECTED_306,
         SYNOPSYS_UNCONNECTED_307, SYNOPSYS_UNCONNECTED_308,
         SYNOPSYS_UNCONNECTED_309, SYNOPSYS_UNCONNECTED_310,
         SYNOPSYS_UNCONNECTED_311, SYNOPSYS_UNCONNECTED_312,
         SYNOPSYS_UNCONNECTED_313, SYNOPSYS_UNCONNECTED_314,
         SYNOPSYS_UNCONNECTED_315, SYNOPSYS_UNCONNECTED_316,
         SYNOPSYS_UNCONNECTED_317, SYNOPSYS_UNCONNECTED_318,
         SYNOPSYS_UNCONNECTED_319, SYNOPSYS_UNCONNECTED_320,
         SYNOPSYS_UNCONNECTED_321, SYNOPSYS_UNCONNECTED_322,
         SYNOPSYS_UNCONNECTED_323, SYNOPSYS_UNCONNECTED_324,
         SYNOPSYS_UNCONNECTED_325, SYNOPSYS_UNCONNECTED_326,
         SYNOPSYS_UNCONNECTED_327, SYNOPSYS_UNCONNECTED_328,
         SYNOPSYS_UNCONNECTED_329, SYNOPSYS_UNCONNECTED_330,
         SYNOPSYS_UNCONNECTED_331, SYNOPSYS_UNCONNECTED_332,
         SYNOPSYS_UNCONNECTED_333, SYNOPSYS_UNCONNECTED_334,
         SYNOPSYS_UNCONNECTED_335, SYNOPSYS_UNCONNECTED_336,
         SYNOPSYS_UNCONNECTED_337, SYNOPSYS_UNCONNECTED_338,
         SYNOPSYS_UNCONNECTED_339, SYNOPSYS_UNCONNECTED_340,
         SYNOPSYS_UNCONNECTED_341, SYNOPSYS_UNCONNECTED_342,
         SYNOPSYS_UNCONNECTED_343, SYNOPSYS_UNCONNECTED_344,
         SYNOPSYS_UNCONNECTED_345, SYNOPSYS_UNCONNECTED_346,
         SYNOPSYS_UNCONNECTED_347, SYNOPSYS_UNCONNECTED_348,
         SYNOPSYS_UNCONNECTED_349, SYNOPSYS_UNCONNECTED_350,
         SYNOPSYS_UNCONNECTED_351, SYNOPSYS_UNCONNECTED_352,
         SYNOPSYS_UNCONNECTED_353, SYNOPSYS_UNCONNECTED_354,
         SYNOPSYS_UNCONNECTED_355, SYNOPSYS_UNCONNECTED_356,
         SYNOPSYS_UNCONNECTED_357, SYNOPSYS_UNCONNECTED_358,
         SYNOPSYS_UNCONNECTED_359, SYNOPSYS_UNCONNECTED_360,
         SYNOPSYS_UNCONNECTED_361, SYNOPSYS_UNCONNECTED_362,
         SYNOPSYS_UNCONNECTED_363, SYNOPSYS_UNCONNECTED_364,
         SYNOPSYS_UNCONNECTED_365, SYNOPSYS_UNCONNECTED_366,
         SYNOPSYS_UNCONNECTED_367, SYNOPSYS_UNCONNECTED_368,
         SYNOPSYS_UNCONNECTED_369, SYNOPSYS_UNCONNECTED_370,
         SYNOPSYS_UNCONNECTED_371, SYNOPSYS_UNCONNECTED_372,
         SYNOPSYS_UNCONNECTED_373, SYNOPSYS_UNCONNECTED_374,
         SYNOPSYS_UNCONNECTED_375, SYNOPSYS_UNCONNECTED_376,
         SYNOPSYS_UNCONNECTED_377, SYNOPSYS_UNCONNECTED_378,
         SYNOPSYS_UNCONNECTED_379, SYNOPSYS_UNCONNECTED_380,
         SYNOPSYS_UNCONNECTED_381, SYNOPSYS_UNCONNECTED_382,
         SYNOPSYS_UNCONNECTED_383, SYNOPSYS_UNCONNECTED_384,
         SYNOPSYS_UNCONNECTED_385, SYNOPSYS_UNCONNECTED_386,
         SYNOPSYS_UNCONNECTED_387, SYNOPSYS_UNCONNECTED_388,
         SYNOPSYS_UNCONNECTED_389, SYNOPSYS_UNCONNECTED_390,
         SYNOPSYS_UNCONNECTED_391, SYNOPSYS_UNCONNECTED_392,
         SYNOPSYS_UNCONNECTED_393, SYNOPSYS_UNCONNECTED_394,
         SYNOPSYS_UNCONNECTED_395, SYNOPSYS_UNCONNECTED_396,
         SYNOPSYS_UNCONNECTED_397, SYNOPSYS_UNCONNECTED_398,
         SYNOPSYS_UNCONNECTED_399, SYNOPSYS_UNCONNECTED_400,
         SYNOPSYS_UNCONNECTED_401, SYNOPSYS_UNCONNECTED_402,
         SYNOPSYS_UNCONNECTED_403, SYNOPSYS_UNCONNECTED_404,
         SYNOPSYS_UNCONNECTED_405, SYNOPSYS_UNCONNECTED_406,
         SYNOPSYS_UNCONNECTED_407, SYNOPSYS_UNCONNECTED_408,
         SYNOPSYS_UNCONNECTED_409, SYNOPSYS_UNCONNECTED_410,
         SYNOPSYS_UNCONNECTED_411, SYNOPSYS_UNCONNECTED_412;
  wire   [26:2] boothout1;
  wire   [26:0] boothout2;
  wire   [26:0] boothout3;
  wire   [26:0] boothout4;
  wire   [26:0] boothout5;
  wire   [26:0] boothout6;
  wire   [26:0] boothout7;
  wire   [26:0] boothout8;
  wire   [26:0] boothout9;
  wire   [26:0] boothout10;
  wire   [26:0] boothout11;
  wire   [25:0] boothout12;
  wire   [22:0] boothout13;
  wire   [29:2] cout1;
  wire   [31:3] mulout1;
  wire   [35:8] cout2;
  wire   [37:6] mulout2;
  wire   [41:14] cout3;
  wire   [42:12] mulout3;
  wire   [46:20] cout4;
  wire   [47:18] mulout4;
  wire   [31:3] cout5;
  wire   [46:4] mulout5;
  wire   [37:9] cout6;
  wire   [42:6] mulout6;
  wire   [46:18] cout7;
  wire   [47:12] mulout7;
  wire   [38:4] cout8;
  wire   [46:5] mulout8;
  wire   [46:12] cout9;
  wire   [47:6] mulout9;
  wire   [46:5] cout10;
  wire   [47:6] mulout10;
  wire   [46:6] cout11;
  wire   [47:7] mulout11;
  wire   [47:0] a;
  wire   [47:8] b;

  booth27_13 booth1 ( .out1({boothout1, SYNOPSYS_UNCONNECTED_1, 
        SYNOPSYS_UNCONNECTED_2}), .in1({in1[1:0], 1'b0}), .in2({1'b0, 1'b0, 
        1'b1, n31, n30, n29, n28, in2[18], n27, n26, in2[15], n25, n24, n23, 
        in2[11:8], n21, in2[6], n20, in2[4], n19, in2[2], n18, n17}) );
  booth27_12 booth2 ( .out1(boothout2), .in1(in1[3:1]), .in2({1'b0, 1'b0, 1'b1, 
        n31, n30, n29, n28, in2[18], n27, n26, in2[15], n25, n24, n23, 
        in2[11:8], n21, in2[6], n20, in2[4], n19, in2[2], n18, n17}) );
  booth27_11 booth3 ( .out1(boothout3), .in1(in1[5:3]), .in2({1'b0, 1'b0, 1'b1, 
        n31, n30, n29, n28, in2[18], n27, n26, in2[15], n25, n24, n23, 
        in2[11:6], n20, in2[4], n19, in2[2], n18, n17}) );
  booth27_10 booth4 ( .out1(boothout4), .in1(in1[7:5]), .in2({1'b0, 1'b0, 1'b1, 
        n31, n30, n29, n28, in2[18], n27, n26, in2[15], n25, n24, n23, 
        in2[11:8], n21, in2[6], n20, in2[4], n19, in2[2], n18, n17}) );
  booth27_9 booth5 ( .out1(boothout5), .in1(in1[9:7]), .in2({1'b0, 1'b0, 1'b1, 
        n31, n30, n29, n28, in2[18], n27, n26, in2[15], n25, n24, n23, 
        in2[11:6], n20, in2[4], n19, in2[2], n18, n17}) );
  booth27_8 booth6 ( .out1(boothout6), .in1(in1[11:9]), .in2({1'b0, 1'b0, 1'b1, 
        n31, n30, n29, n28, in2[18], n27, n26, in2[15], n25, n24, n23, 
        in2[11:6], n20, in2[4], n19, in2[2], n18, n17}) );
  booth27_7 booth7 ( .out1(boothout7), .in1(in1[13:11]), .in2({1'b0, 1'b0, 
        1'b1, n31, n30, n29, n28, in2[18], n27, n26, in2[15], n25, n24, n23, 
        in2[11:6], n20, in2[4], n19, in2[2], n18, n17}) );
  booth27_6 booth8 ( .out1(boothout8), .in1(in1[15:13]), .in2({1'b0, 1'b0, 
        1'b1, n31, n30, n29, n28, in2[18], n27, n26, in2[15], n25, n24, n23, 
        in2[11:6], n20, in2[4], n19, in2[2], n18, n17}) );
  booth27_5 booth9 ( .out1(boothout9), .in1(in1[17:15]), .in2({1'b0, 1'b0, 
        1'b1, n31, n30, n29, n28, in2[18], n27, n26, in2[15], n25, n24, n23, 
        in2[11:6], n20, in2[4], n19, in2[2], n18, n17}) );
  booth27_4 booth10 ( .out1(boothout10), .in1(in1[19:17]), .in2({1'b0, 1'b0, 
        1'b1, n31, n30, n29, n28, in2[18], n27, n26, in2[15], n25, n24, n23, 
        in2[11:6], n20, in2[4], n19, in2[2], n18, n17}) );
  booth27_3 booth11 ( .out1(boothout11), .in1(in1[21:19]), .in2({1'b0, 1'b0, 
        1'b1, n31, n30, n29, n28, in2[18], n27, n26, in2[15], n25, n24, n23, 
        in2[11:6], n20, in2[4], n19, in2[2], n18, n17}) );
  booth27_2 booth12 ( .out1({SYNOPSYS_UNCONNECTED_3, boothout12}), .in1({1'b1, 
        in1[22:21]}), .in2({1'b0, 1'b0, 1'b1, n31, n30, n29, n28, in2[18], n27, 
        n26, in2[15], n25, n24, n23, in2[11:8], n21, in2[6], n20, in2[4], n19, 
        in2[2], n18, n17}) );
  booth27_1 booth13 ( .out1({SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, 
        SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, boothout13}), .in1({
        1'b0, 1'b0, 1'b1}), .in2({1'b0, 1'b0, 1'b1, n31, n30, n29, n28, 
        in2[18], n27, n26, in2[15], n25, n24, n23, in2[11:8], n21, in2[6], n20, 
        in2[4], n19, in2[2], n18, n17}) );
  csa51squ_12 csa51squ1 ( .cout({SYNOPSYS_UNCONNECTED_8, 
        SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10, 
        SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12, 
        SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14, 
        SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16, 
        SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18, 
        SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20, 
        SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22, 
        SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24, 
        SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26, 
        SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28, cout1, 
        SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30}), .sumout({
        SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32, 
        SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34, 
        SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36, 
        SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38, 
        SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40, 
        SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42, 
        SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44, 
        SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46, 
        SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48, 
        SYNOPSYS_UNCONNECTED_49, mulout1[31], SYNOPSYS_UNCONNECTED_50, 
        mulout1[29:3], SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52, 
        SYNOPSYS_UNCONNECTED_53}), .in1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, boothout1, 1'b0, 1'b0}), .in2({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, boothout2, 
        1'b0, 1'b0}), .in3({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n129, 
        1'b0, boothout3[25:0], 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_11 csa51squ2 ( .cout({SYNOPSYS_UNCONNECTED_54, 
        SYNOPSYS_UNCONNECTED_55, SYNOPSYS_UNCONNECTED_56, 
        SYNOPSYS_UNCONNECTED_57, SYNOPSYS_UNCONNECTED_58, 
        SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_60, 
        SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_62, 
        SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_64, 
        SYNOPSYS_UNCONNECTED_65, SYNOPSYS_UNCONNECTED_66, 
        SYNOPSYS_UNCONNECTED_67, SYNOPSYS_UNCONNECTED_68, cout2, 
        SYNOPSYS_UNCONNECTED_69, SYNOPSYS_UNCONNECTED_70, 
        SYNOPSYS_UNCONNECTED_71, SYNOPSYS_UNCONNECTED_72, 
        SYNOPSYS_UNCONNECTED_73, SYNOPSYS_UNCONNECTED_74, 
        SYNOPSYS_UNCONNECTED_75, SYNOPSYS_UNCONNECTED_76}), .sumout({
        SYNOPSYS_UNCONNECTED_77, SYNOPSYS_UNCONNECTED_78, 
        SYNOPSYS_UNCONNECTED_79, SYNOPSYS_UNCONNECTED_80, 
        SYNOPSYS_UNCONNECTED_81, SYNOPSYS_UNCONNECTED_82, 
        SYNOPSYS_UNCONNECTED_83, SYNOPSYS_UNCONNECTED_84, 
        SYNOPSYS_UNCONNECTED_85, SYNOPSYS_UNCONNECTED_86, 
        SYNOPSYS_UNCONNECTED_87, SYNOPSYS_UNCONNECTED_88, 
        SYNOPSYS_UNCONNECTED_89, mulout2[37], SYNOPSYS_UNCONNECTED_90, 
        mulout2[35:6], SYNOPSYS_UNCONNECTED_91, SYNOPSYS_UNCONNECTED_92, 
        SYNOPSYS_UNCONNECTED_93, SYNOPSYS_UNCONNECTED_94, 
        SYNOPSYS_UNCONNECTED_95, SYNOPSYS_UNCONNECTED_96}), .in1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, boothout4, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, boothout5, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .in3({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n128, 1'b0, boothout6[25:0], 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_10 csa51squ3 ( .cout({SYNOPSYS_UNCONNECTED_97, 
        SYNOPSYS_UNCONNECTED_98, SYNOPSYS_UNCONNECTED_99, 
        SYNOPSYS_UNCONNECTED_100, SYNOPSYS_UNCONNECTED_101, 
        SYNOPSYS_UNCONNECTED_102, SYNOPSYS_UNCONNECTED_103, 
        SYNOPSYS_UNCONNECTED_104, SYNOPSYS_UNCONNECTED_105, cout3, 
        SYNOPSYS_UNCONNECTED_106, SYNOPSYS_UNCONNECTED_107, 
        SYNOPSYS_UNCONNECTED_108, SYNOPSYS_UNCONNECTED_109, 
        SYNOPSYS_UNCONNECTED_110, SYNOPSYS_UNCONNECTED_111, 
        SYNOPSYS_UNCONNECTED_112, SYNOPSYS_UNCONNECTED_113, 
        SYNOPSYS_UNCONNECTED_114, SYNOPSYS_UNCONNECTED_115, 
        SYNOPSYS_UNCONNECTED_116, SYNOPSYS_UNCONNECTED_117, 
        SYNOPSYS_UNCONNECTED_118, SYNOPSYS_UNCONNECTED_119}), .sumout({
        SYNOPSYS_UNCONNECTED_120, SYNOPSYS_UNCONNECTED_121, 
        SYNOPSYS_UNCONNECTED_122, SYNOPSYS_UNCONNECTED_123, 
        SYNOPSYS_UNCONNECTED_124, SYNOPSYS_UNCONNECTED_125, 
        SYNOPSYS_UNCONNECTED_126, SYNOPSYS_UNCONNECTED_127, mulout3, 
        SYNOPSYS_UNCONNECTED_128, SYNOPSYS_UNCONNECTED_129, 
        SYNOPSYS_UNCONNECTED_130, SYNOPSYS_UNCONNECTED_131, 
        SYNOPSYS_UNCONNECTED_132, SYNOPSYS_UNCONNECTED_133, 
        SYNOPSYS_UNCONNECTED_134, SYNOPSYS_UNCONNECTED_135, 
        SYNOPSYS_UNCONNECTED_136, SYNOPSYS_UNCONNECTED_137, 
        SYNOPSYS_UNCONNECTED_138, SYNOPSYS_UNCONNECTED_139}), .in1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, boothout7, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, boothout8, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .in3({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        boothout9, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_9 csa51squ4 ( .cout({SYNOPSYS_UNCONNECTED_140, 
        SYNOPSYS_UNCONNECTED_141, SYNOPSYS_UNCONNECTED_142, 
        SYNOPSYS_UNCONNECTED_143, cout4, SYNOPSYS_UNCONNECTED_144, 
        SYNOPSYS_UNCONNECTED_145, SYNOPSYS_UNCONNECTED_146, 
        SYNOPSYS_UNCONNECTED_147, SYNOPSYS_UNCONNECTED_148, 
        SYNOPSYS_UNCONNECTED_149, SYNOPSYS_UNCONNECTED_150, 
        SYNOPSYS_UNCONNECTED_151, SYNOPSYS_UNCONNECTED_152, 
        SYNOPSYS_UNCONNECTED_153, SYNOPSYS_UNCONNECTED_154, 
        SYNOPSYS_UNCONNECTED_155, SYNOPSYS_UNCONNECTED_156, 
        SYNOPSYS_UNCONNECTED_157, SYNOPSYS_UNCONNECTED_158, 
        SYNOPSYS_UNCONNECTED_159, SYNOPSYS_UNCONNECTED_160, 
        SYNOPSYS_UNCONNECTED_161, SYNOPSYS_UNCONNECTED_162, 
        SYNOPSYS_UNCONNECTED_163}), .sumout({SYNOPSYS_UNCONNECTED_164, 
        SYNOPSYS_UNCONNECTED_165, SYNOPSYS_UNCONNECTED_166, mulout4, 
        SYNOPSYS_UNCONNECTED_167, SYNOPSYS_UNCONNECTED_168, 
        SYNOPSYS_UNCONNECTED_169, SYNOPSYS_UNCONNECTED_170, 
        SYNOPSYS_UNCONNECTED_171, SYNOPSYS_UNCONNECTED_172, 
        SYNOPSYS_UNCONNECTED_173, SYNOPSYS_UNCONNECTED_174, 
        SYNOPSYS_UNCONNECTED_175, SYNOPSYS_UNCONNECTED_176, 
        SYNOPSYS_UNCONNECTED_177, SYNOPSYS_UNCONNECTED_178, 
        SYNOPSYS_UNCONNECTED_179, SYNOPSYS_UNCONNECTED_180, 
        SYNOPSYS_UNCONNECTED_181, SYNOPSYS_UNCONNECTED_182, 
        SYNOPSYS_UNCONNECTED_183, SYNOPSYS_UNCONNECTED_184}), .in1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, boothout10, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 1'b0, 1'b0, 1'b0, boothout11, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .in3({1'b0, 1'b0, 1'b0, boothout12, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_8 csa51squ5 ( .cout({SYNOPSYS_UNCONNECTED_185, 
        SYNOPSYS_UNCONNECTED_186, SYNOPSYS_UNCONNECTED_187, 
        SYNOPSYS_UNCONNECTED_188, SYNOPSYS_UNCONNECTED_189, 
        SYNOPSYS_UNCONNECTED_190, SYNOPSYS_UNCONNECTED_191, 
        SYNOPSYS_UNCONNECTED_192, SYNOPSYS_UNCONNECTED_193, 
        SYNOPSYS_UNCONNECTED_194, SYNOPSYS_UNCONNECTED_195, 
        SYNOPSYS_UNCONNECTED_196, SYNOPSYS_UNCONNECTED_197, 
        SYNOPSYS_UNCONNECTED_198, SYNOPSYS_UNCONNECTED_199, 
        SYNOPSYS_UNCONNECTED_200, SYNOPSYS_UNCONNECTED_201, 
        SYNOPSYS_UNCONNECTED_202, SYNOPSYS_UNCONNECTED_203, cout5, 
        SYNOPSYS_UNCONNECTED_204, SYNOPSYS_UNCONNECTED_205, 
        SYNOPSYS_UNCONNECTED_206}), .sumout({SYNOPSYS_UNCONNECTED_207, 
        SYNOPSYS_UNCONNECTED_208, SYNOPSYS_UNCONNECTED_209, 
        SYNOPSYS_UNCONNECTED_210, mulout5, SYNOPSYS_UNCONNECTED_211, 
        SYNOPSYS_UNCONNECTED_212, SYNOPSYS_UNCONNECTED_213, 
        SYNOPSYS_UNCONNECTED_214}), .in1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, cout1, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, mulout1[31], 1'b0, mulout1[29:3], 1'b0, 1'b0, 1'b0}), 
        .in3({1'b0, 1'b0, 1'b0, 1'b1, boothout13, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_7 csa51squ6 ( .cout({SYNOPSYS_UNCONNECTED_215, 
        SYNOPSYS_UNCONNECTED_216, SYNOPSYS_UNCONNECTED_217, 
        SYNOPSYS_UNCONNECTED_218, SYNOPSYS_UNCONNECTED_219, 
        SYNOPSYS_UNCONNECTED_220, SYNOPSYS_UNCONNECTED_221, 
        SYNOPSYS_UNCONNECTED_222, SYNOPSYS_UNCONNECTED_223, 
        SYNOPSYS_UNCONNECTED_224, SYNOPSYS_UNCONNECTED_225, 
        SYNOPSYS_UNCONNECTED_226, SYNOPSYS_UNCONNECTED_227, cout6, 
        SYNOPSYS_UNCONNECTED_228, SYNOPSYS_UNCONNECTED_229, 
        SYNOPSYS_UNCONNECTED_230, SYNOPSYS_UNCONNECTED_231, 
        SYNOPSYS_UNCONNECTED_232, SYNOPSYS_UNCONNECTED_233, 
        SYNOPSYS_UNCONNECTED_234, SYNOPSYS_UNCONNECTED_235, 
        SYNOPSYS_UNCONNECTED_236}), .sumout({SYNOPSYS_UNCONNECTED_237, 
        SYNOPSYS_UNCONNECTED_238, SYNOPSYS_UNCONNECTED_239, 
        SYNOPSYS_UNCONNECTED_240, SYNOPSYS_UNCONNECTED_241, 
        SYNOPSYS_UNCONNECTED_242, SYNOPSYS_UNCONNECTED_243, 
        SYNOPSYS_UNCONNECTED_244, mulout6, SYNOPSYS_UNCONNECTED_245, 
        SYNOPSYS_UNCONNECTED_246, SYNOPSYS_UNCONNECTED_247, 
        SYNOPSYS_UNCONNECTED_248, SYNOPSYS_UNCONNECTED_249, 
        SYNOPSYS_UNCONNECTED_250}), .in1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, cout2, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        mulout2[37], 1'b0, mulout2[35:6], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .in3({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, cout3, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  csa51squ_6 csa51squ7 ( .cout({SYNOPSYS_UNCONNECTED_251, 
        SYNOPSYS_UNCONNECTED_252, SYNOPSYS_UNCONNECTED_253, 
        SYNOPSYS_UNCONNECTED_254, cout7, SYNOPSYS_UNCONNECTED_255, 
        SYNOPSYS_UNCONNECTED_256, SYNOPSYS_UNCONNECTED_257, 
        SYNOPSYS_UNCONNECTED_258, SYNOPSYS_UNCONNECTED_259, 
        SYNOPSYS_UNCONNECTED_260, SYNOPSYS_UNCONNECTED_261, 
        SYNOPSYS_UNCONNECTED_262, SYNOPSYS_UNCONNECTED_263, 
        SYNOPSYS_UNCONNECTED_264, SYNOPSYS_UNCONNECTED_265, 
        SYNOPSYS_UNCONNECTED_266, SYNOPSYS_UNCONNECTED_267, 
        SYNOPSYS_UNCONNECTED_268, SYNOPSYS_UNCONNECTED_269, 
        SYNOPSYS_UNCONNECTED_270, SYNOPSYS_UNCONNECTED_271, 
        SYNOPSYS_UNCONNECTED_272}), .sumout({SYNOPSYS_UNCONNECTED_273, 
        SYNOPSYS_UNCONNECTED_274, SYNOPSYS_UNCONNECTED_275, mulout7, 
        SYNOPSYS_UNCONNECTED_276, SYNOPSYS_UNCONNECTED_277, 
        SYNOPSYS_UNCONNECTED_278, SYNOPSYS_UNCONNECTED_279, 
        SYNOPSYS_UNCONNECTED_280, SYNOPSYS_UNCONNECTED_281, 
        SYNOPSYS_UNCONNECTED_282, SYNOPSYS_UNCONNECTED_283, 
        SYNOPSYS_UNCONNECTED_284, SYNOPSYS_UNCONNECTED_285, 
        SYNOPSYS_UNCONNECTED_286, SYNOPSYS_UNCONNECTED_287}), .in1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mulout3, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 1'b0, 
        1'b0, cout4, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in3({1'b0, 1'b0, 1'b0, mulout4, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_5 csa51squ8 ( .cout({SYNOPSYS_UNCONNECTED_288, 
        SYNOPSYS_UNCONNECTED_289, SYNOPSYS_UNCONNECTED_290, 
        SYNOPSYS_UNCONNECTED_291, SYNOPSYS_UNCONNECTED_292, 
        SYNOPSYS_UNCONNECTED_293, SYNOPSYS_UNCONNECTED_294, 
        SYNOPSYS_UNCONNECTED_295, SYNOPSYS_UNCONNECTED_296, 
        SYNOPSYS_UNCONNECTED_297, SYNOPSYS_UNCONNECTED_298, 
        SYNOPSYS_UNCONNECTED_299, cout8, SYNOPSYS_UNCONNECTED_300, 
        SYNOPSYS_UNCONNECTED_301, SYNOPSYS_UNCONNECTED_302, 
        SYNOPSYS_UNCONNECTED_303}), .sumout({SYNOPSYS_UNCONNECTED_304, 
        SYNOPSYS_UNCONNECTED_305, SYNOPSYS_UNCONNECTED_306, 
        SYNOPSYS_UNCONNECTED_307, mulout8, SYNOPSYS_UNCONNECTED_308, 
        SYNOPSYS_UNCONNECTED_309, SYNOPSYS_UNCONNECTED_310, 
        SYNOPSYS_UNCONNECTED_311, SYNOPSYS_UNCONNECTED_312}), .in1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, cout5, 1'b0, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 
        1'b0, 1'b0, 1'b1, mulout5, 1'b0, 1'b0, 1'b0, 1'b0}), .in3({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, cout6, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_4 csa51squ9 ( .cout({SYNOPSYS_UNCONNECTED_313, 
        SYNOPSYS_UNCONNECTED_314, SYNOPSYS_UNCONNECTED_315, 
        SYNOPSYS_UNCONNECTED_316, cout9, SYNOPSYS_UNCONNECTED_317, 
        SYNOPSYS_UNCONNECTED_318, SYNOPSYS_UNCONNECTED_319, 
        SYNOPSYS_UNCONNECTED_320, SYNOPSYS_UNCONNECTED_321, 
        SYNOPSYS_UNCONNECTED_322, SYNOPSYS_UNCONNECTED_323, 
        SYNOPSYS_UNCONNECTED_324, SYNOPSYS_UNCONNECTED_325, 
        SYNOPSYS_UNCONNECTED_326, SYNOPSYS_UNCONNECTED_327, 
        SYNOPSYS_UNCONNECTED_328}), .sumout({SYNOPSYS_UNCONNECTED_329, 
        SYNOPSYS_UNCONNECTED_330, SYNOPSYS_UNCONNECTED_331, mulout9, 
        SYNOPSYS_UNCONNECTED_332, SYNOPSYS_UNCONNECTED_333, 
        SYNOPSYS_UNCONNECTED_334, SYNOPSYS_UNCONNECTED_335, 
        SYNOPSYS_UNCONNECTED_336, SYNOPSYS_UNCONNECTED_337}), .in1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mulout6, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .in2({1'b0, 1'b0, 1'b0, cout7, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .in3({1'b0, 1'b0, 1'b0, mulout7, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_3 csa51squ10 ( .cout({SYNOPSYS_UNCONNECTED_338, 
        SYNOPSYS_UNCONNECTED_339, SYNOPSYS_UNCONNECTED_340, 
        SYNOPSYS_UNCONNECTED_341, cout10, SYNOPSYS_UNCONNECTED_342, 
        SYNOPSYS_UNCONNECTED_343, SYNOPSYS_UNCONNECTED_344, 
        SYNOPSYS_UNCONNECTED_345, SYNOPSYS_UNCONNECTED_346}), .sumout({
        SYNOPSYS_UNCONNECTED_347, SYNOPSYS_UNCONNECTED_348, 
        SYNOPSYS_UNCONNECTED_349, mulout10, SYNOPSYS_UNCONNECTED_350, 
        SYNOPSYS_UNCONNECTED_351, SYNOPSYS_UNCONNECTED_352, 
        SYNOPSYS_UNCONNECTED_353, SYNOPSYS_UNCONNECTED_354, 
        SYNOPSYS_UNCONNECTED_355}), .in1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, cout8, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .in2({1'b0, 1'b0, 1'b0, 1'b1, mulout8, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .in3({1'b0, 1'b0, 1'b0, cout9, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_2 csa51squ11 ( .cout({SYNOPSYS_UNCONNECTED_356, 
        SYNOPSYS_UNCONNECTED_357, SYNOPSYS_UNCONNECTED_358, 
        SYNOPSYS_UNCONNECTED_359, cout11, SYNOPSYS_UNCONNECTED_360, 
        SYNOPSYS_UNCONNECTED_361, SYNOPSYS_UNCONNECTED_362, 
        SYNOPSYS_UNCONNECTED_363, SYNOPSYS_UNCONNECTED_364, 
        SYNOPSYS_UNCONNECTED_365}), .sumout({SYNOPSYS_UNCONNECTED_366, 
        SYNOPSYS_UNCONNECTED_367, SYNOPSYS_UNCONNECTED_368, mulout11, 
        SYNOPSYS_UNCONNECTED_369, SYNOPSYS_UNCONNECTED_370, 
        SYNOPSYS_UNCONNECTED_371, SYNOPSYS_UNCONNECTED_372, 
        SYNOPSYS_UNCONNECTED_373, SYNOPSYS_UNCONNECTED_374, 
        SYNOPSYS_UNCONNECTED_375}), .in1({1'b0, 1'b0, 1'b0, mulout9, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 1'b0, 1'b0, cout10, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in3({1'b0, 1'b0, 1'b0, mulout10, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_1 csa51squ12 ( .sumout({SYNOPSYS_UNCONNECTED_376, 
        SYNOPSYS_UNCONNECTED_377, SYNOPSYS_UNCONNECTED_378, N101, N100, N99, 
        N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, 
        N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, 
        N70, N69, N68, N67, N66, N65, N64, N63, N62, SYNOPSYS_UNCONNECTED_379, 
        SYNOPSYS_UNCONNECTED_380, SYNOPSYS_UNCONNECTED_381, 
        SYNOPSYS_UNCONNECTED_382, SYNOPSYS_UNCONNECTED_383, 
        SYNOPSYS_UNCONNECTED_384, SYNOPSYS_UNCONNECTED_385, 
        SYNOPSYS_UNCONNECTED_386}), .in1({1'b0, 1'b0, 1'b0, mulout11, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 1'b0, 1'b0, cout11, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in3({1'b1, 1'b0, 1'b1, 
        1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 
        1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .cout_46_(N50), .cout_44_(N48), .cout_42_(N46), .cout_40_(N44), .cout_38_(
        N42), .cout_36_(N40), .cout_34_(N38), .cout_32_(N36), .cout_30_(N34), 
        .cout_28_(N32), .cout_27_(N31), .cout_7__BAR(N11), .cout_8__BAR(N12), 
        .cout_9__BAR(N13), .cout_10__BAR(N14), .cout_11__BAR(N15), 
        .cout_12__BAR(N16), .cout_13__BAR(N17), .cout_14__BAR(N18), 
        .cout_15__BAR(N19), .cout_16__BAR(N20), .cout_17__BAR(N21), 
        .cout_18__BAR(N22), .cout_19__BAR(N23), .cout_20__BAR(N24), 
        .cout_21__BAR(N25), .cout_22__BAR(N26), .cout_23__BAR(N27), 
        .cout_24__BAR(N28), .cout_25__BAR(N29), .cout_26__BAR(N30), 
        .cout_29__BAR(N33), .cout_31__BAR(N35), .cout_33__BAR(N37), 
        .cout_35__BAR(N39), .cout_37__BAR(N41), .cout_39__BAR(N43), 
        .cout_41__BAR(N45), .cout_43__BAR(N47), .cout_45__BAR(N49) );
  cla51squ_1 cla51squ ( .out({SYNOPSYS_UNCONNECTED_387, 
        SYNOPSYS_UNCONNECTED_388, SYNOPSYS_UNCONNECTED_389, mulout[47:23], 
        SYNOPSYS_UNCONNECTED_390, SYNOPSYS_UNCONNECTED_391, 
        SYNOPSYS_UNCONNECTED_392, SYNOPSYS_UNCONNECTED_393, 
        SYNOPSYS_UNCONNECTED_394, SYNOPSYS_UNCONNECTED_395, 
        SYNOPSYS_UNCONNECTED_396, SYNOPSYS_UNCONNECTED_397, 
        SYNOPSYS_UNCONNECTED_398, SYNOPSYS_UNCONNECTED_399, 
        SYNOPSYS_UNCONNECTED_400, SYNOPSYS_UNCONNECTED_401, 
        SYNOPSYS_UNCONNECTED_402, SYNOPSYS_UNCONNECTED_403, 
        SYNOPSYS_UNCONNECTED_404, SYNOPSYS_UNCONNECTED_405, 
        SYNOPSYS_UNCONNECTED_406, SYNOPSYS_UNCONNECTED_407, 
        SYNOPSYS_UNCONNECTED_408, SYNOPSYS_UNCONNECTED_409, 
        SYNOPSYS_UNCONNECTED_410, SYNOPSYS_UNCONNECTED_411, 
        SYNOPSYS_UNCONNECTED_412}), .a({1'b0, 1'b0, 1'b0, a[47:8], 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({1'b0, 1'b0, 1'b0, b, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  DFFARX1 b_reg_47_ ( .D(N101), .CLK(clk), .RSTB(rst_n), .Q(b[47]) );
  DFFARX1 b_reg_46_ ( .D(N100), .CLK(clk), .RSTB(rst_n), .Q(b[46]) );
  DFFARX1 b_reg_45_ ( .D(N99), .CLK(clk), .RSTB(rst_n), .Q(b[45]) );
  DFFARX1 b_reg_44_ ( .D(N98), .CLK(clk), .RSTB(rst_n), .Q(b[44]) );
  DFFARX1 b_reg_43_ ( .D(N97), .CLK(clk), .RSTB(rst_n), .Q(b[43]) );
  DFFARX1 b_reg_42_ ( .D(N96), .CLK(clk), .RSTB(rst_n), .Q(b[42]) );
  DFFARX1 b_reg_41_ ( .D(N95), .CLK(clk), .RSTB(rst_n), .Q(b[41]) );
  DFFARX1 b_reg_40_ ( .D(N94), .CLK(clk), .RSTB(rst_n), .Q(b[40]) );
  DFFARX1 b_reg_39_ ( .D(N93), .CLK(clk), .RSTB(rst_n), .Q(b[39]) );
  DFFARX1 b_reg_38_ ( .D(N92), .CLK(clk), .RSTB(rst_n), .Q(b[38]) );
  DFFARX1 b_reg_37_ ( .D(N91), .CLK(clk), .RSTB(rst_n), .Q(b[37]) );
  DFFARX1 b_reg_36_ ( .D(N90), .CLK(clk), .RSTB(rst_n), .Q(b[36]) );
  DFFARX1 b_reg_35_ ( .D(N89), .CLK(clk), .RSTB(rst_n), .Q(b[35]) );
  DFFARX1 b_reg_34_ ( .D(N88), .CLK(clk), .RSTB(rst_n), .Q(b[34]) );
  DFFARX1 b_reg_33_ ( .D(N87), .CLK(clk), .RSTB(rst_n), .Q(b[33]) );
  DFFARX1 b_reg_32_ ( .D(N86), .CLK(clk), .RSTB(rst_n), .Q(b[32]) );
  DFFARX1 b_reg_31_ ( .D(N85), .CLK(clk), .RSTB(rst_n), .Q(b[31]) );
  DFFARX1 b_reg_30_ ( .D(N84), .CLK(clk), .RSTB(rst_n), .Q(b[30]) );
  DFFARX1 b_reg_29_ ( .D(N83), .CLK(clk), .RSTB(rst_n), .Q(b[29]) );
  DFFARX1 b_reg_28_ ( .D(N82), .CLK(clk), .RSTB(rst_n), .Q(b[28]) );
  DFFARX1 b_reg_27_ ( .D(N81), .CLK(clk), .RSTB(rst_n), .Q(b[27]) );
  DFFARX1 b_reg_26_ ( .D(N80), .CLK(clk), .RSTB(rst_n), .Q(b[26]) );
  DFFARX1 b_reg_25_ ( .D(N79), .CLK(clk), .RSTB(rst_n), .Q(b[25]) );
  DFFARX1 b_reg_24_ ( .D(N78), .CLK(clk), .RSTB(rst_n), .Q(b[24]) );
  DFFARX1 b_reg_23_ ( .D(N77), .CLK(clk), .RSTB(rst_n), .Q(b[23]) );
  DFFARX1 b_reg_22_ ( .D(N76), .CLK(clk), .RSTB(rst_n), .Q(b[22]) );
  DFFARX1 b_reg_21_ ( .D(N75), .CLK(clk), .RSTB(rst_n), .Q(b[21]) );
  DFFARX1 b_reg_20_ ( .D(N74), .CLK(clk), .RSTB(rst_n), .Q(b[20]) );
  DFFARX1 b_reg_19_ ( .D(N73), .CLK(clk), .RSTB(rst_n), .Q(b[19]) );
  DFFARX1 b_reg_18_ ( .D(N72), .CLK(clk), .RSTB(rst_n), .Q(b[18]) );
  DFFARX1 b_reg_17_ ( .D(N71), .CLK(clk), .RSTB(rst_n), .Q(b[17]) );
  DFFARX1 b_reg_16_ ( .D(N70), .CLK(clk), .RSTB(rst_n), .Q(b[16]) );
  DFFARX1 b_reg_15_ ( .D(N69), .CLK(clk), .RSTB(rst_n), .Q(b[15]) );
  DFFARX1 b_reg_14_ ( .D(N68), .CLK(clk), .RSTB(rst_n), .Q(b[14]) );
  DFFARX1 b_reg_13_ ( .D(N67), .CLK(clk), .RSTB(rst_n), .Q(b[13]) );
  DFFARX1 b_reg_12_ ( .D(N66), .CLK(clk), .RSTB(rst_n), .Q(b[12]) );
  DFFARX1 b_reg_11_ ( .D(N65), .CLK(clk), .RSTB(rst_n), .Q(b[11]) );
  DFFARX1 b_reg_10_ ( .D(N64), .CLK(clk), .RSTB(rst_n), .Q(b[10]) );
  DFFARX1 b_reg_9_ ( .D(N63), .CLK(clk), .RSTB(rst_n), .Q(b[9]) );
  DFFARX1 b_reg_8_ ( .D(N62), .CLK(clk), .RSTB(rst_n), .Q(b[8]) );
  DFFARX1 a_reg_47_ ( .D(N50), .CLK(clk), .RSTB(rst_n), .Q(a[47]) );
  DFFARX1 a_reg_46_ ( .D(n60), .CLK(clk), .RSTB(rst_n), .Q(a[46]) );
  DFFARX1 a_reg_45_ ( .D(N48), .CLK(clk), .RSTB(rst_n), .Q(a[45]) );
  DFFARX1 a_reg_44_ ( .D(n61), .CLK(clk), .RSTB(rst_n), .Q(a[44]) );
  DFFARX1 a_reg_43_ ( .D(N46), .CLK(clk), .RSTB(rst_n), .Q(a[43]) );
  DFFARX1 a_reg_42_ ( .D(n62), .CLK(clk), .RSTB(rst_n), .Q(a[42]) );
  DFFARX1 a_reg_41_ ( .D(N44), .CLK(clk), .RSTB(rst_n), .Q(a[41]) );
  DFFARX1 a_reg_40_ ( .D(n63), .CLK(clk), .RSTB(rst_n), .Q(a[40]) );
  DFFARX1 a_reg_39_ ( .D(N42), .CLK(clk), .RSTB(rst_n), .Q(a[39]) );
  DFFARX1 a_reg_38_ ( .D(n64), .CLK(clk), .RSTB(rst_n), .Q(a[38]) );
  DFFARX1 a_reg_37_ ( .D(N40), .CLK(clk), .RSTB(rst_n), .Q(a[37]) );
  DFFARX1 a_reg_36_ ( .D(n65), .CLK(clk), .RSTB(rst_n), .Q(a[36]) );
  DFFARX1 a_reg_35_ ( .D(N38), .CLK(clk), .RSTB(rst_n), .Q(a[35]) );
  DFFARX1 a_reg_34_ ( .D(n66), .CLK(clk), .RSTB(rst_n), .Q(a[34]) );
  DFFARX1 a_reg_33_ ( .D(N36), .CLK(clk), .RSTB(rst_n), .Q(a[33]) );
  DFFARX1 a_reg_32_ ( .D(n67), .CLK(clk), .RSTB(rst_n), .Q(a[32]) );
  DFFARX1 a_reg_31_ ( .D(N34), .CLK(clk), .RSTB(rst_n), .Q(a[31]) );
  DFFARX1 a_reg_30_ ( .D(n68), .CLK(clk), .RSTB(rst_n), .Q(a[30]) );
  DFFARX1 a_reg_29_ ( .D(N32), .CLK(clk), .RSTB(rst_n), .Q(a[29]) );
  DFFARX1 a_reg_28_ ( .D(N31), .CLK(clk), .RSTB(rst_n), .Q(a[28]) );
  DFFARX1 a_reg_27_ ( .D(n69), .CLK(clk), .RSTB(rst_n), .Q(a[27]) );
  DFFARX1 a_reg_26_ ( .D(n70), .CLK(clk), .RSTB(rst_n), .Q(a[26]) );
  DFFARX1 a_reg_25_ ( .D(n71), .CLK(clk), .RSTB(rst_n), .Q(a[25]) );
  DFFARX1 a_reg_24_ ( .D(n72), .CLK(clk), .RSTB(rst_n), .Q(a[24]) );
  DFFARX1 a_reg_23_ ( .D(n73), .CLK(clk), .RSTB(rst_n), .Q(a[23]) );
  DFFARX1 a_reg_22_ ( .D(n74), .CLK(clk), .RSTB(rst_n), .Q(a[22]) );
  DFFARX1 a_reg_21_ ( .D(n75), .CLK(clk), .RSTB(rst_n), .Q(a[21]) );
  DFFARX1 a_reg_20_ ( .D(n76), .CLK(clk), .RSTB(rst_n), .Q(a[20]) );
  DFFARX1 a_reg_19_ ( .D(n77), .CLK(clk), .RSTB(rst_n), .Q(a[19]) );
  DFFARX1 a_reg_18_ ( .D(n78), .CLK(clk), .RSTB(rst_n), .Q(a[18]) );
  DFFARX1 a_reg_17_ ( .D(n79), .CLK(clk), .RSTB(rst_n), .Q(a[17]) );
  DFFARX1 a_reg_16_ ( .D(n80), .CLK(clk), .RSTB(rst_n), .Q(a[16]) );
  DFFARX1 a_reg_15_ ( .D(n81), .CLK(clk), .RSTB(rst_n), .Q(a[15]) );
  DFFARX1 a_reg_14_ ( .D(n82), .CLK(clk), .RSTB(rst_n), .Q(a[14]) );
  DFFARX1 a_reg_13_ ( .D(n83), .CLK(clk), .RSTB(rst_n), .Q(a[13]) );
  DFFARX1 a_reg_12_ ( .D(n84), .CLK(clk), .RSTB(rst_n), .Q(a[12]) );
  DFFARX1 a_reg_11_ ( .D(n85), .CLK(clk), .RSTB(rst_n), .Q(a[11]) );
  DFFARX1 a_reg_10_ ( .D(n86), .CLK(clk), .RSTB(rst_n), .Q(a[10]) );
  DFFARX1 a_reg_9_ ( .D(n87), .CLK(clk), .RSTB(rst_n), .Q(a[9]) );
  DFFARX1 a_reg_8_ ( .D(n88), .CLK(clk), .RSTB(rst_n), .Q(a[8]) );
  INVX0 U5 ( .INP(boothout3[26]), .ZN(n129) );
  INVX0 U8 ( .INP(boothout6[26]), .ZN(n128) );
  NBUFFX8 U3 ( .INP(in2[16]), .Z(n26) );
  NBUFFX8 U4 ( .INP(in2[14]), .Z(n25) );
  NBUFFX8 U6 ( .INP(in2[20]), .Z(n29) );
  NBUFFX8 U7 ( .INP(in2[19]), .Z(n28) );
  NBUFFX8 U9 ( .INP(in2[13]), .Z(n24) );
  NBUFFX8 U10 ( .INP(in2[17]), .Z(n27) );
  NBUFFX8 U11 ( .INP(in2[21]), .Z(n30) );
  NBUFFX8 U12 ( .INP(in2[22]), .Z(n31) );
  NBUFFX8 U13 ( .INP(in2[3]), .Z(n19) );
  NBUFFX8 U14 ( .INP(in2[5]), .Z(n20) );
  INVX0 U15 ( .INP(n22), .ZN(n21) );
  NBUFFX2 U16 ( .INP(in2[12]), .Z(n23) );
  NBUFFX8 U17 ( .INP(in2[1]), .Z(n18) );
  NBUFFX8 U18 ( .INP(in2[0]), .Z(n17) );
  INVX0 U33 ( .INP(in2[7]), .ZN(n22) );
  INVX0 U69 ( .INP(N49), .ZN(n60) );
  INVX0 U70 ( .INP(N47), .ZN(n61) );
  INVX0 U71 ( .INP(N45), .ZN(n62) );
  INVX0 U72 ( .INP(N43), .ZN(n63) );
  INVX0 U73 ( .INP(N41), .ZN(n64) );
  INVX0 U74 ( .INP(N39), .ZN(n65) );
  INVX0 U75 ( .INP(N37), .ZN(n66) );
  INVX0 U76 ( .INP(N35), .ZN(n67) );
  INVX0 U77 ( .INP(N33), .ZN(n68) );
  INVX0 U78 ( .INP(N30), .ZN(n69) );
  INVX0 U79 ( .INP(N29), .ZN(n70) );
  INVX0 U80 ( .INP(N28), .ZN(n71) );
  INVX0 U81 ( .INP(N27), .ZN(n72) );
  INVX0 U82 ( .INP(N26), .ZN(n73) );
  INVX0 U83 ( .INP(N25), .ZN(n74) );
  INVX0 U84 ( .INP(N24), .ZN(n75) );
  INVX0 U85 ( .INP(N23), .ZN(n76) );
  INVX0 U86 ( .INP(N22), .ZN(n77) );
  INVX0 U87 ( .INP(N21), .ZN(n78) );
  INVX0 U88 ( .INP(N20), .ZN(n79) );
  INVX0 U89 ( .INP(N19), .ZN(n80) );
  INVX0 U90 ( .INP(N18), .ZN(n81) );
  INVX0 U91 ( .INP(N17), .ZN(n82) );
  INVX0 U92 ( .INP(N16), .ZN(n83) );
  INVX0 U93 ( .INP(N15), .ZN(n84) );
  INVX0 U94 ( .INP(N14), .ZN(n85) );
  INVX0 U95 ( .INP(N13), .ZN(n86) );
  INVX0 U96 ( .INP(N12), .ZN(n87) );
  INVX0 U97 ( .INP(N11), .ZN(n88) );
endmodule


module add_97 ( s, a, b, co, ci_BAR );
  input a, b, ci_BAR;
  output s, co;


  XOR2X1 U1 ( .IN1(a), .IN2(ci_BAR), .Q(s) );
endmodule


module add_98 ( s, a, b, ci, co_BAR );
  input a, b, ci;
  output s, co_BAR;


  NAND2X0 U1 ( .IN1(ci), .IN2(a), .QN(co_BAR) );
  OA21X1 U2 ( .IN1(ci), .IN2(a), .IN3(co_BAR), .Q(s) );
endmodule


module add_99 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_100 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_101 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_102 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_103 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  INVX0 U1 ( .INP(a), .ZN(s) );
  NBUFFX2 U2 ( .INP(a), .Z(co) );
endmodule


module add_104 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  NBUFFX2 U1 ( .INP(a), .Z(s) );
endmodule


module adder8_7 ( out, a, b, cin );
  output [7:0] out;
  input [7:0] a;
  input [7:0] b;
  input cin;

  wire   [6:1] c;

  add_104 add_01 ( .s(out[0]), .a(a[0]), .b(1'b1), .ci(1'b1) );
  add_103 add_02 ( .s(out[1]), .a(a[1]), .b(1'b0), .ci(1'b1), .co(c[1]) );
  add_102 add_03 ( .s(out[2]), .a(a[2]), .b(1'b0), .ci(c[1]), .co(c[2]) );
  add_101 add_04 ( .s(out[3]), .a(a[3]), .b(1'b0), .ci(c[2]), .co(c[3]) );
  add_100 add_05 ( .s(out[4]), .a(a[4]), .b(1'b0), .ci(c[3]), .co(c[4]) );
  add_99 add_06 ( .s(out[5]), .a(a[5]), .b(1'b0), .ci(c[4]), .co(c[5]) );
  add_98 add_07 ( .s(out[6]), .a(a[6]), .b(1'b0), .ci(c[5]), .co_BAR(c[6]) );
  add_97 add_08 ( .s(out[7]), .a(a[7]), .b(1'b1), .ci_BAR(c[6]) );
endmodule


module add_105 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  XOR3X1 U1 ( .IN1(b), .IN2(ci), .IN3(a), .Q(s) );
endmodule


module add_106 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_107 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_108 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_109 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_110 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_111 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_112 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(b), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(b), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module adder8_8 ( out, a, b, cin );
  output [7:0] out;
  input [7:0] a;
  input [7:0] b;
  input cin;

  wire   [6:0] c;

  add_112 add_01 ( .s(out[0]), .a(a[0]), .b(b[0]), .ci(1'b0), .co(c[0]) );
  add_111 add_02 ( .s(out[1]), .a(a[1]), .b(b[1]), .ci(c[0]), .co(c[1]) );
  add_110 add_03 ( .s(out[2]), .a(a[2]), .b(b[2]), .ci(c[1]), .co(c[2]) );
  add_109 add_04 ( .s(out[3]), .a(a[3]), .b(b[3]), .ci(c[2]), .co(c[3]) );
  add_108 add_05 ( .s(out[4]), .a(a[4]), .b(b[4]), .ci(c[3]), .co(c[4]) );
  add_107 add_06 ( .s(out[5]), .a(a[5]), .b(b[5]), .ci(c[4]), .co(c[5]) );
  add_106 add_07 ( .s(out[6]), .a(a[6]), .b(b[6]), .ci(c[5]), .co(c[6]) );
  add_105 add_08 ( .s(out[7]), .a(a[7]), .b(b[7]), .ci(c[6]) );
endmodule


module floating_point_multiple_1 ( clk, rst_n, input_factor_01, 
        input_factor_02, output_multiply );
  input [31:0] input_factor_01;
  input [31:0] input_factor_02;
  output [31:0] output_multiply;
  input clk, rst_n;
  wire   N5, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22,
         N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N48, N49, N50, N51,
         N52, N53, N54, N55, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22,
         SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24,
         SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26;
  wire   [47:23] base_multiply_result;
  wire   [47:23] mulout;
  wire   [7:0] exponent_factor_12;
  wire   [7:0] pre_mul_output_exponent;

  mul26_1 mul26_01 ( .clk(clk), .rst_n(rst_n), .in1({1'b0, 1'b0, 1'b1, 
        input_factor_01[22:0]}), .in2({1'b0, 1'b0, 1'b1, input_factor_02[22:0]}), .en(1'b1), .mulout({SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, 
        SYNOPSYS_UNCONNECTED_3, mulout, SYNOPSYS_UNCONNECTED_4, 
        SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, 
        SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, 
        SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11, 
        SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13, 
        SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, 
        SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17, 
        SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19, 
        SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21, 
        SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_23, 
        SYNOPSYS_UNCONNECTED_24, SYNOPSYS_UNCONNECTED_25, 
        SYNOPSYS_UNCONNECTED_26}) );
  adder8_8 adder8_01 ( .out(exponent_factor_12), .a(input_factor_01[30:23]), 
        .b(input_factor_02[30:23]), .cin(1'b0) );
  adder8_7 adder8_02 ( .out(pre_mul_output_exponent), .a(exponent_factor_12), 
        .b({1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0}), .cin(1'b1) );
  DFFARX1 mul_output_sign_reg ( .D(N5), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[31]) );
  DFFARX1 base_multiply_result_reg_47_ ( .D(mulout[47]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[47]) );
  DFFARX1 base_multiply_result_reg_46_ ( .D(mulout[46]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[46]) );
  DFFARX1 base_multiply_result_reg_45_ ( .D(mulout[45]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[45]) );
  DFFARX1 base_multiply_result_reg_44_ ( .D(mulout[44]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[44]) );
  DFFARX1 base_multiply_result_reg_43_ ( .D(mulout[43]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[43]) );
  DFFARX1 base_multiply_result_reg_42_ ( .D(mulout[42]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[42]) );
  DFFARX1 base_multiply_result_reg_41_ ( .D(mulout[41]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[41]) );
  DFFARX1 base_multiply_result_reg_40_ ( .D(mulout[40]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[40]) );
  DFFARX1 base_multiply_result_reg_39_ ( .D(mulout[39]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[39]) );
  DFFARX1 base_multiply_result_reg_38_ ( .D(mulout[38]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[38]) );
  DFFARX1 base_multiply_result_reg_37_ ( .D(mulout[37]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[37]) );
  DFFARX1 base_multiply_result_reg_36_ ( .D(mulout[36]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[36]) );
  DFFARX1 base_multiply_result_reg_35_ ( .D(mulout[35]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[35]) );
  DFFARX1 base_multiply_result_reg_34_ ( .D(mulout[34]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[34]) );
  DFFARX1 base_multiply_result_reg_33_ ( .D(mulout[33]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[33]) );
  DFFARX1 base_multiply_result_reg_32_ ( .D(mulout[32]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[32]) );
  DFFARX1 base_multiply_result_reg_31_ ( .D(mulout[31]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[31]) );
  DFFARX1 base_multiply_result_reg_30_ ( .D(mulout[30]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[30]) );
  DFFARX1 base_multiply_result_reg_29_ ( .D(mulout[29]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[29]) );
  DFFARX1 base_multiply_result_reg_28_ ( .D(mulout[28]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[28]) );
  DFFARX1 base_multiply_result_reg_27_ ( .D(mulout[27]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[27]) );
  DFFARX1 base_multiply_result_reg_26_ ( .D(mulout[26]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[26]) );
  DFFARX1 base_multiply_result_reg_25_ ( .D(mulout[25]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[25]) );
  DFFARX1 base_multiply_result_reg_24_ ( .D(mulout[24]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[24]) );
  DFFARX1 base_multiply_result_reg_23_ ( .D(mulout[23]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[23]) );
  DFFARX1 mul_output_significand_reg_22_ ( .D(N32), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[22]) );
  DFFARX1 mul_output_significand_reg_21_ ( .D(N31), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[21]) );
  DFFARX1 mul_output_significand_reg_20_ ( .D(N30), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[20]) );
  DFFARX1 mul_output_significand_reg_19_ ( .D(N29), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[19]) );
  DFFARX1 mul_output_significand_reg_18_ ( .D(N28), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[18]) );
  DFFARX1 mul_output_significand_reg_17_ ( .D(N27), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[17]) );
  DFFARX1 mul_output_significand_reg_16_ ( .D(N26), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[16]) );
  DFFARX1 mul_output_significand_reg_15_ ( .D(N25), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[15]) );
  DFFARX1 mul_output_significand_reg_14_ ( .D(N24), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[14]) );
  DFFARX1 mul_output_significand_reg_13_ ( .D(N23), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[13]) );
  DFFARX1 mul_output_significand_reg_12_ ( .D(N22), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[12]) );
  DFFARX1 mul_output_significand_reg_11_ ( .D(N21), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[11]) );
  DFFARX1 mul_output_significand_reg_10_ ( .D(N20), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[10]) );
  DFFARX1 mul_output_significand_reg_9_ ( .D(N19), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[9]) );
  DFFARX1 mul_output_significand_reg_8_ ( .D(N18), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[8]) );
  DFFARX1 mul_output_significand_reg_7_ ( .D(N17), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[7]) );
  DFFARX1 mul_output_significand_reg_6_ ( .D(N16), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[6]) );
  DFFARX1 mul_output_significand_reg_5_ ( .D(N15), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[5]) );
  DFFARX1 mul_output_significand_reg_4_ ( .D(N14), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[4]) );
  DFFARX1 mul_output_significand_reg_3_ ( .D(N13), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[3]) );
  DFFARX1 mul_output_significand_reg_2_ ( .D(N12), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[2]) );
  DFFARX1 mul_output_significand_reg_1_ ( .D(N11), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[1]) );
  DFFARX1 mul_output_significand_reg_0_ ( .D(N10), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[0]) );
  DFFARX1 mul_output_exponent_reg_7_ ( .D(N55), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[30]) );
  DFFARX1 mul_output_exponent_reg_6_ ( .D(N54), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[29]) );
  DFFARX1 mul_output_exponent_reg_5_ ( .D(N53), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[28]) );
  DFFARX1 mul_output_exponent_reg_4_ ( .D(N52), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[27]) );
  DFFARX1 mul_output_exponent_reg_3_ ( .D(N51), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[26]) );
  DFFARX1 mul_output_exponent_reg_2_ ( .D(N50), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[25]) );
  DFFARX1 mul_output_exponent_reg_1_ ( .D(N49), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[24]) );
  DFFARX1 mul_output_exponent_reg_0_ ( .D(N48), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[23]) );
  AND2X1 U3 ( .IN1(base_multiply_result[47]), .IN2(n35), .Q(n32) );
  INVX0 U4 ( .INP(n1), .ZN(n2) );
  OR2X1 U5 ( .IN1(base_multiply_result[47]), .IN2(n24), .Q(n1) );
  INVX0 U6 ( .INP(input_factor_02[31]), .ZN(n3) );
  NOR4X0 U7 ( .IN1(input_factor_01[0]), .IN2(input_factor_01[10]), .IN3(
        input_factor_01[11]), .IN4(input_factor_01[12]), .QN(n7) );
  NOR4X0 U8 ( .IN1(input_factor_01[13]), .IN2(input_factor_01[14]), .IN3(
        input_factor_01[15]), .IN4(input_factor_01[16]), .QN(n6) );
  NOR4X0 U9 ( .IN1(input_factor_01[17]), .IN2(input_factor_01[18]), .IN3(
        input_factor_01[19]), .IN4(input_factor_01[1]), .QN(n5) );
  NOR4X0 U10 ( .IN1(input_factor_01[20]), .IN2(input_factor_01[21]), .IN3(
        input_factor_01[22]), .IN4(input_factor_01[23]), .QN(n4) );
  NAND4X0 U11 ( .IN1(n7), .IN2(n6), .IN3(n5), .IN4(n4), .QN(n23) );
  NOR4X0 U12 ( .IN1(input_factor_01[24]), .IN2(input_factor_01[25]), .IN3(
        input_factor_01[26]), .IN4(input_factor_01[27]), .QN(n11) );
  NOR4X0 U13 ( .IN1(input_factor_01[28]), .IN2(input_factor_01[29]), .IN3(
        input_factor_01[2]), .IN4(input_factor_01[30]), .QN(n10) );
  NOR4X0 U14 ( .IN1(input_factor_01[31]), .IN2(input_factor_01[3]), .IN3(
        input_factor_01[4]), .IN4(input_factor_01[5]), .QN(n9) );
  NOR4X0 U15 ( .IN1(input_factor_01[6]), .IN2(input_factor_01[7]), .IN3(
        input_factor_01[8]), .IN4(input_factor_01[9]), .QN(n8) );
  NAND4X0 U16 ( .IN1(n11), .IN2(n10), .IN3(n9), .IN4(n8), .QN(n22) );
  NOR4X0 U17 ( .IN1(input_factor_02[0]), .IN2(input_factor_02[10]), .IN3(
        input_factor_02[11]), .IN4(input_factor_02[12]), .QN(n15) );
  NOR4X0 U18 ( .IN1(input_factor_02[13]), .IN2(input_factor_02[14]), .IN3(
        input_factor_02[15]), .IN4(input_factor_02[16]), .QN(n14) );
  NOR4X0 U19 ( .IN1(input_factor_02[17]), .IN2(input_factor_02[18]), .IN3(
        input_factor_02[19]), .IN4(input_factor_02[1]), .QN(n13) );
  NOR4X0 U20 ( .IN1(input_factor_02[20]), .IN2(input_factor_02[21]), .IN3(
        input_factor_02[22]), .IN4(input_factor_02[23]), .QN(n12) );
  NAND4X0 U21 ( .IN1(n15), .IN2(n14), .IN3(n13), .IN4(n12), .QN(n21) );
  NOR4X0 U22 ( .IN1(input_factor_02[24]), .IN2(input_factor_02[25]), .IN3(
        input_factor_02[26]), .IN4(input_factor_02[27]), .QN(n19) );
  NOR4X0 U23 ( .IN1(input_factor_02[28]), .IN2(input_factor_02[29]), .IN3(
        input_factor_02[2]), .IN4(input_factor_02[30]), .QN(n18) );
  NOR4X0 U24 ( .IN1(input_factor_02[31]), .IN2(input_factor_02[3]), .IN3(
        input_factor_02[4]), .IN4(input_factor_02[5]), .QN(n17) );
  NOR4X0 U25 ( .IN1(input_factor_02[6]), .IN2(input_factor_02[7]), .IN3(
        input_factor_02[8]), .IN4(input_factor_02[9]), .QN(n16) );
  NAND4X0 U26 ( .IN1(n19), .IN2(n18), .IN3(n17), .IN4(n16), .QN(n20) );
  OA22X1 U27 ( .IN1(n23), .IN2(n22), .IN3(n21), .IN4(n20), .Q(n35) );
  INVX0 U28 ( .INP(n35), .ZN(n24) );
  AO22X1 U29 ( .IN1(n2), .IN2(base_multiply_result[23]), .IN3(n32), .IN4(
        base_multiply_result[24]), .Q(N10) );
  AO22X1 U30 ( .IN1(n2), .IN2(base_multiply_result[24]), .IN3(n32), .IN4(
        base_multiply_result[25]), .Q(N11) );
  AO22X1 U31 ( .IN1(n2), .IN2(base_multiply_result[25]), .IN3(n32), .IN4(
        base_multiply_result[26]), .Q(N12) );
  AO22X1 U32 ( .IN1(n2), .IN2(base_multiply_result[26]), .IN3(n32), .IN4(
        base_multiply_result[27]), .Q(N13) );
  AO22X1 U33 ( .IN1(n2), .IN2(base_multiply_result[27]), .IN3(n32), .IN4(
        base_multiply_result[28]), .Q(N14) );
  AO22X1 U34 ( .IN1(n2), .IN2(base_multiply_result[28]), .IN3(n32), .IN4(
        base_multiply_result[29]), .Q(N15) );
  AO22X1 U35 ( .IN1(n2), .IN2(base_multiply_result[29]), .IN3(n32), .IN4(
        base_multiply_result[30]), .Q(N16) );
  AO22X1 U36 ( .IN1(n2), .IN2(base_multiply_result[30]), .IN3(n32), .IN4(
        base_multiply_result[31]), .Q(N17) );
  AO22X1 U37 ( .IN1(n2), .IN2(base_multiply_result[31]), .IN3(n32), .IN4(
        base_multiply_result[32]), .Q(N18) );
  AO22X1 U38 ( .IN1(n2), .IN2(base_multiply_result[32]), .IN3(n32), .IN4(
        base_multiply_result[33]), .Q(N19) );
  AO22X1 U39 ( .IN1(n2), .IN2(base_multiply_result[33]), .IN3(n32), .IN4(
        base_multiply_result[34]), .Q(N20) );
  AO22X1 U40 ( .IN1(n2), .IN2(base_multiply_result[34]), .IN3(n32), .IN4(
        base_multiply_result[35]), .Q(N21) );
  AO22X1 U41 ( .IN1(n2), .IN2(base_multiply_result[35]), .IN3(n32), .IN4(
        base_multiply_result[36]), .Q(N22) );
  AO22X1 U42 ( .IN1(n2), .IN2(base_multiply_result[36]), .IN3(n32), .IN4(
        base_multiply_result[37]), .Q(N23) );
  AO22X1 U43 ( .IN1(n2), .IN2(base_multiply_result[37]), .IN3(n32), .IN4(
        base_multiply_result[38]), .Q(N24) );
  AO22X1 U44 ( .IN1(n2), .IN2(base_multiply_result[38]), .IN3(n32), .IN4(
        base_multiply_result[39]), .Q(N25) );
  AO22X1 U45 ( .IN1(n2), .IN2(base_multiply_result[39]), .IN3(n32), .IN4(
        base_multiply_result[40]), .Q(N26) );
  AO22X1 U46 ( .IN1(n2), .IN2(base_multiply_result[40]), .IN3(n32), .IN4(
        base_multiply_result[41]), .Q(N27) );
  AO22X1 U47 ( .IN1(n2), .IN2(base_multiply_result[41]), .IN3(n32), .IN4(
        base_multiply_result[42]), .Q(N28) );
  AO22X1 U48 ( .IN1(n2), .IN2(base_multiply_result[42]), .IN3(n32), .IN4(
        base_multiply_result[43]), .Q(N29) );
  AO22X1 U49 ( .IN1(n2), .IN2(base_multiply_result[43]), .IN3(n32), .IN4(
        base_multiply_result[44]), .Q(N30) );
  AO22X1 U50 ( .IN1(n2), .IN2(base_multiply_result[44]), .IN3(n32), .IN4(
        base_multiply_result[45]), .Q(N31) );
  AO22X1 U51 ( .IN1(n2), .IN2(base_multiply_result[45]), .IN3(n32), .IN4(
        base_multiply_result[46]), .Q(N32) );
  MUX21X1 U52 ( .IN1(n2), .IN2(n32), .S(pre_mul_output_exponent[0]), .Q(N48)
         );
  AO21X1 U53 ( .IN1(pre_mul_output_exponent[0]), .IN2(n2), .IN3(n32), .Q(n25)
         );
  NOR3X0 U54 ( .IN1(pre_mul_output_exponent[1]), .IN2(
        pre_mul_output_exponent[0]), .IN3(n1), .QN(n27) );
  AO21X1 U55 ( .IN1(pre_mul_output_exponent[1]), .IN2(n25), .IN3(n27), .Q(N49)
         );
  INVX0 U56 ( .INP(input_factor_01[31]), .ZN(n26) );
  OA221X1 U57 ( .IN1(input_factor_01[31]), .IN2(input_factor_02[31]), .IN3(n26), .IN4(n3), .IN5(n35), .Q(N5) );
  AO221X1 U58 ( .IN1(n2), .IN2(pre_mul_output_exponent[1]), .IN3(n2), .IN4(
        pre_mul_output_exponent[0]), .IN5(n32), .Q(n28) );
  MUX21X1 U59 ( .IN1(n27), .IN2(n28), .S(pre_mul_output_exponent[2]), .Q(N50)
         );
  AND2X1 U60 ( .IN1(n2), .IN2(pre_mul_output_exponent[2]), .Q(n29) );
  OR4X1 U61 ( .IN1(pre_mul_output_exponent[1]), .IN2(
        pre_mul_output_exponent[0]), .IN3(pre_mul_output_exponent[3]), .IN4(
        pre_mul_output_exponent[2]), .Q(n34) );
  NOR2X0 U62 ( .IN1(n1), .IN2(n34), .QN(n31) );
  AO221X1 U63 ( .IN1(pre_mul_output_exponent[3]), .IN2(n29), .IN3(
        pre_mul_output_exponent[3]), .IN4(n28), .IN5(n31), .Q(N51) );
  OA21X1 U64 ( .IN1(base_multiply_result[47]), .IN2(n34), .IN3(n35), .Q(n30)
         );
  MUX21X1 U65 ( .IN1(n31), .IN2(n30), .S(pre_mul_output_exponent[4]), .Q(N52)
         );
  AO221X1 U66 ( .IN1(n2), .IN2(pre_mul_output_exponent[4]), .IN3(n2), .IN4(n34), .IN5(n32), .Q(n33) );
  NOR4X0 U67 ( .IN1(pre_mul_output_exponent[5]), .IN2(
        pre_mul_output_exponent[4]), .IN3(n34), .IN4(n1), .QN(n37) );
  AO21X1 U68 ( .IN1(pre_mul_output_exponent[5]), .IN2(n33), .IN3(n37), .Q(N53)
         );
  OR3X1 U69 ( .IN1(pre_mul_output_exponent[5]), .IN2(
        pre_mul_output_exponent[4]), .IN3(n34), .Q(n36) );
  OA21X1 U70 ( .IN1(base_multiply_result[47]), .IN2(n36), .IN3(n35), .Q(n39)
         );
  INVX0 U71 ( .INP(n37), .ZN(n38) );
  NOR2X0 U72 ( .IN1(pre_mul_output_exponent[6]), .IN2(n38), .QN(n41) );
  AO21X1 U73 ( .IN1(pre_mul_output_exponent[6]), .IN2(n39), .IN3(n41), .Q(N54)
         );
  AO21X1 U74 ( .IN1(n2), .IN2(pre_mul_output_exponent[6]), .IN3(n39), .Q(n40)
         );
  MUX21X1 U75 ( .IN1(n41), .IN2(n40), .S(pre_mul_output_exponent[7]), .Q(N55)
         );
endmodule


module cla51squ_2 ( out, a, b );
  output [50:0] out;
  input [50:0] a;
  input [50:0] b;
  wire   intadd_2_CI, intadd_2_n24, intadd_2_n23, intadd_2_n22, intadd_2_n21,
         intadd_2_n20, intadd_2_n19, intadd_2_n18, intadd_2_n17, intadd_2_n16,
         intadd_2_n15, intadd_2_n14, intadd_2_n13, intadd_2_n12, intadd_2_n11,
         intadd_2_n10, intadd_2_n9, intadd_2_n8, intadd_2_n7, intadd_2_n6,
         intadd_2_n5, intadd_2_n4, intadd_2_n3, intadd_2_n2, intadd_2_n1, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14;

  FADDX1 intadd_2_U25 ( .A(b[23]), .B(a[23]), .CI(intadd_2_CI), .CO(
        intadd_2_n24), .S(out[23]) );
  FADDX1 intadd_2_U24 ( .A(b[24]), .B(a[24]), .CI(intadd_2_n24), .CO(
        intadd_2_n23), .S(out[24]) );
  FADDX1 intadd_2_U23 ( .A(b[25]), .B(a[25]), .CI(intadd_2_n23), .CO(
        intadd_2_n22), .S(out[25]) );
  FADDX1 intadd_2_U22 ( .A(b[26]), .B(a[26]), .CI(intadd_2_n22), .CO(
        intadd_2_n21), .S(out[26]) );
  FADDX1 intadd_2_U21 ( .A(b[27]), .B(a[27]), .CI(intadd_2_n21), .CO(
        intadd_2_n20), .S(out[27]) );
  FADDX1 intadd_2_U20 ( .A(b[28]), .B(a[28]), .CI(intadd_2_n20), .CO(
        intadd_2_n19), .S(out[28]) );
  FADDX1 intadd_2_U19 ( .A(b[29]), .B(a[29]), .CI(intadd_2_n19), .CO(
        intadd_2_n18), .S(out[29]) );
  FADDX1 intadd_2_U18 ( .A(b[30]), .B(a[30]), .CI(intadd_2_n18), .CO(
        intadd_2_n17), .S(out[30]) );
  FADDX1 intadd_2_U17 ( .A(b[31]), .B(a[31]), .CI(intadd_2_n17), .CO(
        intadd_2_n16), .S(out[31]) );
  FADDX1 intadd_2_U16 ( .A(b[32]), .B(a[32]), .CI(intadd_2_n16), .CO(
        intadd_2_n15), .S(out[32]) );
  FADDX1 intadd_2_U15 ( .A(b[33]), .B(a[33]), .CI(intadd_2_n15), .CO(
        intadd_2_n14), .S(out[33]) );
  FADDX1 intadd_2_U14 ( .A(b[34]), .B(a[34]), .CI(intadd_2_n14), .CO(
        intadd_2_n13), .S(out[34]) );
  FADDX1 intadd_2_U13 ( .A(b[35]), .B(a[35]), .CI(intadd_2_n13), .CO(
        intadd_2_n12), .S(out[35]) );
  FADDX1 intadd_2_U12 ( .A(b[36]), .B(a[36]), .CI(intadd_2_n12), .CO(
        intadd_2_n11), .S(out[36]) );
  FADDX1 intadd_2_U11 ( .A(b[37]), .B(a[37]), .CI(intadd_2_n11), .CO(
        intadd_2_n10), .S(out[37]) );
  FADDX1 intadd_2_U10 ( .A(b[38]), .B(a[38]), .CI(intadd_2_n10), .CO(
        intadd_2_n9), .S(out[38]) );
  FADDX1 intadd_2_U9 ( .A(b[39]), .B(a[39]), .CI(intadd_2_n9), .CO(intadd_2_n8), .S(out[39]) );
  FADDX1 intadd_2_U8 ( .A(b[40]), .B(a[40]), .CI(intadd_2_n8), .CO(intadd_2_n7), .S(out[40]) );
  FADDX1 intadd_2_U7 ( .A(b[41]), .B(a[41]), .CI(intadd_2_n7), .CO(intadd_2_n6), .S(out[41]) );
  FADDX1 intadd_2_U6 ( .A(b[42]), .B(a[42]), .CI(intadd_2_n6), .CO(intadd_2_n5), .S(out[42]) );
  FADDX1 intadd_2_U5 ( .A(b[43]), .B(a[43]), .CI(intadd_2_n5), .CO(intadd_2_n4), .S(out[43]) );
  FADDX1 intadd_2_U4 ( .A(b[44]), .B(a[44]), .CI(intadd_2_n4), .CO(intadd_2_n3), .S(out[44]) );
  FADDX1 intadd_2_U3 ( .A(b[45]), .B(a[45]), .CI(intadd_2_n3), .CO(intadd_2_n2), .S(out[45]) );
  FADDX1 intadd_2_U2 ( .A(b[46]), .B(a[46]), .CI(intadd_2_n2), .CO(intadd_2_n1), .S(out[46]) );
  OA21X1 U2 ( .IN1(b[9]), .IN2(a[9]), .IN3(a[8]), .Q(n1) );
  AO22X1 U3 ( .IN1(b[9]), .IN2(a[9]), .IN3(b[8]), .IN4(n1), .Q(n2) );
  AO222X1 U4 ( .IN1(b[10]), .IN2(a[10]), .IN3(b[10]), .IN4(n2), .IN5(a[10]), 
        .IN6(n2), .Q(n3) );
  AO222X1 U5 ( .IN1(b[11]), .IN2(a[11]), .IN3(b[11]), .IN4(n3), .IN5(a[11]), 
        .IN6(n3), .Q(n4) );
  AO222X1 U6 ( .IN1(b[12]), .IN2(a[12]), .IN3(b[12]), .IN4(n4), .IN5(a[12]), 
        .IN6(n4), .Q(n5) );
  AO222X1 U7 ( .IN1(b[13]), .IN2(a[13]), .IN3(b[13]), .IN4(n5), .IN5(a[13]), 
        .IN6(n5), .Q(n6) );
  AO222X1 U8 ( .IN1(b[14]), .IN2(a[14]), .IN3(b[14]), .IN4(n6), .IN5(a[14]), 
        .IN6(n6), .Q(n7) );
  AO222X1 U9 ( .IN1(b[15]), .IN2(a[15]), .IN3(b[15]), .IN4(n7), .IN5(a[15]), 
        .IN6(n7), .Q(n8) );
  AO222X1 U10 ( .IN1(b[16]), .IN2(a[16]), .IN3(b[16]), .IN4(n8), .IN5(a[16]), 
        .IN6(n8), .Q(n9) );
  AO222X1 U11 ( .IN1(b[17]), .IN2(a[17]), .IN3(b[17]), .IN4(n9), .IN5(a[17]), 
        .IN6(n9), .Q(n10) );
  AO222X1 U12 ( .IN1(b[18]), .IN2(a[18]), .IN3(b[18]), .IN4(n10), .IN5(a[18]), 
        .IN6(n10), .Q(n11) );
  AO222X1 U13 ( .IN1(b[19]), .IN2(a[19]), .IN3(b[19]), .IN4(n11), .IN5(a[19]), 
        .IN6(n11), .Q(n12) );
  AO222X1 U14 ( .IN1(b[20]), .IN2(a[20]), .IN3(b[20]), .IN4(n12), .IN5(a[20]), 
        .IN6(n12), .Q(n13) );
  AO222X1 U15 ( .IN1(b[21]), .IN2(a[21]), .IN3(b[21]), .IN4(n13), .IN5(a[21]), 
        .IN6(n13), .Q(n14) );
  AO222X1 U16 ( .IN1(b[22]), .IN2(a[22]), .IN3(b[22]), .IN4(n14), .IN5(a[22]), 
        .IN6(n14), .Q(intadd_2_CI) );
  XOR3X1 U17 ( .IN1(intadd_2_n1), .IN2(a[47]), .IN3(b[47]), .Q(out[47]) );
endmodule


module csa51squ_13 ( sumout, in1, in2, in3, cout_50_, cout_49_, cout_48_, 
        cout_47_, cout_46_, cout_44_, cout_42_, cout_40_, cout_38_, cout_36_, 
        cout_34_, cout_32_, cout_30_, cout_28_, cout_27_, cout_7__BAR, cout_6_, 
        cout_5_, cout_4_, cout_3_, cout_2_, cout_1_, cout_0_, cout_8__BAR, 
        cout_9__BAR, cout_10__BAR, cout_11__BAR, cout_12__BAR, cout_13__BAR, 
        cout_14__BAR, cout_15__BAR, cout_16__BAR, cout_17__BAR, cout_18__BAR, 
        cout_19__BAR, cout_20__BAR, cout_21__BAR, cout_22__BAR, cout_23__BAR, 
        cout_24__BAR, cout_25__BAR, cout_26__BAR, cout_29__BAR, cout_31__BAR, 
        cout_33__BAR, cout_35__BAR, cout_37__BAR, cout_39__BAR, cout_41__BAR, 
        cout_43__BAR, cout_45__BAR );
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  output cout_50_, cout_49_, cout_48_, cout_47_, cout_46_, cout_44_, cout_42_,
         cout_40_, cout_38_, cout_36_, cout_34_, cout_32_, cout_30_, cout_28_,
         cout_27_, cout_7__BAR, cout_6_, cout_5_, cout_4_, cout_3_, cout_2_,
         cout_1_, cout_0_, cout_8__BAR, cout_9__BAR, cout_10__BAR,
         cout_11__BAR, cout_12__BAR, cout_13__BAR, cout_14__BAR, cout_15__BAR,
         cout_16__BAR, cout_17__BAR, cout_18__BAR, cout_19__BAR, cout_20__BAR,
         cout_21__BAR, cout_22__BAR, cout_23__BAR, cout_24__BAR, cout_25__BAR,
         cout_26__BAR, cout_29__BAR, cout_31__BAR, cout_33__BAR, cout_35__BAR,
         cout_37__BAR, cout_39__BAR, cout_41__BAR, cout_43__BAR, cout_45__BAR;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11;

  NAND2X0 U1 ( .IN1(in2[8]), .IN2(in1[8]), .QN(cout_8__BAR) );
  NAND2X0 U2 ( .IN1(in2[9]), .IN2(in1[9]), .QN(cout_9__BAR) );
  NAND2X0 U3 ( .IN1(in2[10]), .IN2(in1[10]), .QN(cout_10__BAR) );
  NAND2X0 U4 ( .IN1(in2[11]), .IN2(in1[11]), .QN(cout_11__BAR) );
  NAND2X0 U5 ( .IN1(in2[12]), .IN2(in1[12]), .QN(cout_12__BAR) );
  NAND2X0 U6 ( .IN1(in2[13]), .IN2(in1[13]), .QN(cout_13__BAR) );
  NAND2X0 U7 ( .IN1(in2[14]), .IN2(in1[14]), .QN(cout_14__BAR) );
  NAND2X0 U8 ( .IN1(in2[15]), .IN2(in1[15]), .QN(cout_15__BAR) );
  NAND2X0 U9 ( .IN1(in2[16]), .IN2(in1[16]), .QN(cout_16__BAR) );
  NAND2X0 U10 ( .IN1(in2[17]), .IN2(in1[17]), .QN(cout_17__BAR) );
  NAND2X0 U11 ( .IN1(in2[18]), .IN2(in1[18]), .QN(cout_18__BAR) );
  NAND2X0 U12 ( .IN1(in2[19]), .IN2(in1[19]), .QN(cout_19__BAR) );
  NAND2X0 U13 ( .IN1(in2[20]), .IN2(in1[20]), .QN(cout_20__BAR) );
  NAND2X0 U14 ( .IN1(in2[21]), .IN2(in1[21]), .QN(cout_21__BAR) );
  NAND2X0 U15 ( .IN1(in2[22]), .IN2(in1[22]), .QN(cout_22__BAR) );
  NAND2X0 U16 ( .IN1(in2[23]), .IN2(in1[23]), .QN(cout_23__BAR) );
  NAND2X0 U17 ( .IN1(in2[24]), .IN2(in1[24]), .QN(cout_24__BAR) );
  NAND2X0 U18 ( .IN1(in2[25]), .IN2(in1[25]), .QN(cout_25__BAR) );
  NAND2X0 U19 ( .IN1(in2[26]), .IN2(in1[26]), .QN(cout_26__BAR) );
  NAND2X0 U20 ( .IN1(in2[29]), .IN2(in1[29]), .QN(cout_29__BAR) );
  NAND2X0 U21 ( .IN1(in2[31]), .IN2(in1[31]), .QN(cout_31__BAR) );
  NAND2X0 U22 ( .IN1(in2[33]), .IN2(in1[33]), .QN(cout_33__BAR) );
  NAND2X0 U23 ( .IN1(in2[35]), .IN2(in1[35]), .QN(cout_35__BAR) );
  NAND2X0 U24 ( .IN1(in2[37]), .IN2(in1[37]), .QN(cout_37__BAR) );
  NAND2X0 U25 ( .IN1(in2[39]), .IN2(in1[39]), .QN(cout_39__BAR) );
  NAND2X0 U26 ( .IN1(in2[41]), .IN2(in1[41]), .QN(cout_41__BAR) );
  NAND2X0 U27 ( .IN1(in2[43]), .IN2(in1[43]), .QN(cout_43__BAR) );
  NAND2X0 U28 ( .IN1(in2[45]), .IN2(in1[45]), .QN(cout_45__BAR) );
  NAND2X0 U29 ( .IN1(in2[7]), .IN2(in1[7]), .QN(cout_7__BAR) );
  NAND2X0 U30 ( .IN1(n1), .IN2(cout_27_), .QN(sumout[27]) );
  NAND2X0 U31 ( .IN1(in1[27]), .IN2(in2[27]), .QN(n1) );
  NAND2X0 U32 ( .IN1(n2), .IN2(cout_28_), .QN(sumout[28]) );
  NAND2X0 U33 ( .IN1(in1[28]), .IN2(in2[28]), .QN(n2) );
  NAND2X0 U34 ( .IN1(n3), .IN2(cout_30_), .QN(sumout[30]) );
  NAND2X0 U35 ( .IN1(in1[30]), .IN2(in2[30]), .QN(n3) );
  NAND2X0 U36 ( .IN1(n4), .IN2(cout_32_), .QN(sumout[32]) );
  NAND2X0 U37 ( .IN1(in1[32]), .IN2(in2[32]), .QN(n4) );
  NAND2X0 U38 ( .IN1(n5), .IN2(cout_34_), .QN(sumout[34]) );
  NAND2X0 U39 ( .IN1(in1[34]), .IN2(in2[34]), .QN(n5) );
  NAND2X0 U40 ( .IN1(n6), .IN2(cout_36_), .QN(sumout[36]) );
  NAND2X0 U41 ( .IN1(in1[36]), .IN2(in2[36]), .QN(n6) );
  NAND2X0 U42 ( .IN1(n7), .IN2(cout_38_), .QN(sumout[38]) );
  NAND2X0 U43 ( .IN1(in1[38]), .IN2(in2[38]), .QN(n7) );
  NAND2X0 U44 ( .IN1(n8), .IN2(cout_40_), .QN(sumout[40]) );
  NAND2X0 U45 ( .IN1(in1[40]), .IN2(in2[40]), .QN(n8) );
  NAND2X0 U46 ( .IN1(n9), .IN2(cout_42_), .QN(sumout[42]) );
  NAND2X0 U47 ( .IN1(in1[42]), .IN2(in2[42]), .QN(n9) );
  NAND2X0 U48 ( .IN1(n10), .IN2(cout_44_), .QN(sumout[44]) );
  NAND2X0 U49 ( .IN1(in1[44]), .IN2(in2[44]), .QN(n10) );
  NAND2X0 U50 ( .IN1(n11), .IN2(cout_46_), .QN(sumout[46]) );
  NAND2X0 U51 ( .IN1(in1[46]), .IN2(in2[46]), .QN(n11) );
  OR2X1 U52 ( .IN1(in2[27]), .IN2(in1[27]), .Q(cout_27_) );
  OR2X1 U53 ( .IN1(in2[28]), .IN2(in1[28]), .Q(cout_28_) );
  OR2X1 U54 ( .IN1(in2[30]), .IN2(in1[30]), .Q(cout_30_) );
  OR2X1 U55 ( .IN1(in2[32]), .IN2(in1[32]), .Q(cout_32_) );
  OR2X1 U56 ( .IN1(in2[34]), .IN2(in1[34]), .Q(cout_34_) );
  OR2X1 U57 ( .IN1(in2[36]), .IN2(in1[36]), .Q(cout_36_) );
  OR2X1 U58 ( .IN1(in2[38]), .IN2(in1[38]), .Q(cout_38_) );
  OR2X1 U59 ( .IN1(in2[40]), .IN2(in1[40]), .Q(cout_40_) );
  OR2X1 U60 ( .IN1(in2[42]), .IN2(in1[42]), .Q(cout_42_) );
  OR2X1 U61 ( .IN1(in2[44]), .IN2(in1[44]), .Q(cout_44_) );
  OR2X1 U62 ( .IN1(in2[46]), .IN2(in1[46]), .Q(cout_46_) );
  OA21X1 U63 ( .IN1(in2[8]), .IN2(in1[8]), .IN3(cout_8__BAR), .Q(sumout[8]) );
  OA21X1 U64 ( .IN1(in2[9]), .IN2(in1[9]), .IN3(cout_9__BAR), .Q(sumout[9]) );
  OA21X1 U65 ( .IN1(in2[10]), .IN2(in1[10]), .IN3(cout_10__BAR), .Q(sumout[10]) );
  OA21X1 U66 ( .IN1(in2[11]), .IN2(in1[11]), .IN3(cout_11__BAR), .Q(sumout[11]) );
  OA21X1 U67 ( .IN1(in2[12]), .IN2(in1[12]), .IN3(cout_12__BAR), .Q(sumout[12]) );
  OA21X1 U68 ( .IN1(in2[13]), .IN2(in1[13]), .IN3(cout_13__BAR), .Q(sumout[13]) );
  OA21X1 U69 ( .IN1(in2[14]), .IN2(in1[14]), .IN3(cout_14__BAR), .Q(sumout[14]) );
  OA21X1 U70 ( .IN1(in2[15]), .IN2(in1[15]), .IN3(cout_15__BAR), .Q(sumout[15]) );
  OA21X1 U71 ( .IN1(in2[16]), .IN2(in1[16]), .IN3(cout_16__BAR), .Q(sumout[16]) );
  OA21X1 U72 ( .IN1(in2[17]), .IN2(in1[17]), .IN3(cout_17__BAR), .Q(sumout[17]) );
  OA21X1 U73 ( .IN1(in2[18]), .IN2(in1[18]), .IN3(cout_18__BAR), .Q(sumout[18]) );
  OA21X1 U74 ( .IN1(in2[19]), .IN2(in1[19]), .IN3(cout_19__BAR), .Q(sumout[19]) );
  OA21X1 U75 ( .IN1(in2[20]), .IN2(in1[20]), .IN3(cout_20__BAR), .Q(sumout[20]) );
  OA21X1 U76 ( .IN1(in2[21]), .IN2(in1[21]), .IN3(cout_21__BAR), .Q(sumout[21]) );
  OA21X1 U77 ( .IN1(in2[22]), .IN2(in1[22]), .IN3(cout_22__BAR), .Q(sumout[22]) );
  OA21X1 U78 ( .IN1(in2[23]), .IN2(in1[23]), .IN3(cout_23__BAR), .Q(sumout[23]) );
  OA21X1 U79 ( .IN1(in2[24]), .IN2(in1[24]), .IN3(cout_24__BAR), .Q(sumout[24]) );
  OA21X1 U80 ( .IN1(in2[25]), .IN2(in1[25]), .IN3(cout_25__BAR), .Q(sumout[25]) );
  OA21X1 U81 ( .IN1(in2[26]), .IN2(in1[26]), .IN3(cout_26__BAR), .Q(sumout[26]) );
  OA21X1 U82 ( .IN1(in2[29]), .IN2(in1[29]), .IN3(cout_29__BAR), .Q(sumout[29]) );
  OA21X1 U83 ( .IN1(in2[31]), .IN2(in1[31]), .IN3(cout_31__BAR), .Q(sumout[31]) );
  OA21X1 U84 ( .IN1(in2[33]), .IN2(in1[33]), .IN3(cout_33__BAR), .Q(sumout[33]) );
  OA21X1 U85 ( .IN1(in2[35]), .IN2(in1[35]), .IN3(cout_35__BAR), .Q(sumout[35]) );
  OA21X1 U86 ( .IN1(in2[37]), .IN2(in1[37]), .IN3(cout_37__BAR), .Q(sumout[37]) );
  OA21X1 U87 ( .IN1(in2[39]), .IN2(in1[39]), .IN3(cout_39__BAR), .Q(sumout[39]) );
  OA21X1 U88 ( .IN1(in2[41]), .IN2(in1[41]), .IN3(cout_41__BAR), .Q(sumout[41]) );
  OA21X1 U89 ( .IN1(in2[43]), .IN2(in1[43]), .IN3(cout_43__BAR), .Q(sumout[43]) );
  OA21X1 U90 ( .IN1(in2[45]), .IN2(in1[45]), .IN3(cout_45__BAR), .Q(sumout[45]) );
  XOR2X1 U91 ( .IN1(in1[47]), .IN2(in2[47]), .Q(sumout[47]) );
endmodule


module csa51squ_14 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;


  AO222X1 U1 ( .IN1(in2[6]), .IN2(in3[6]), .IN3(in2[6]), .IN4(in1[6]), .IN5(
        in3[6]), .IN6(in1[6]), .Q(cout[6]) );
  FADDX1 U2 ( .A(in1[10]), .B(in2[10]), .CI(in3[10]), .CO(cout[10]), .S(
        sumout[10]) );
  FADDX1 U3 ( .A(in1[11]), .B(in2[11]), .CI(in3[11]), .CO(cout[11]), .S(
        sumout[11]) );
  FADDX1 U4 ( .A(in1[12]), .B(in2[12]), .CI(in3[12]), .CO(cout[12]), .S(
        sumout[12]) );
  FADDX1 U5 ( .A(in1[13]), .B(in2[13]), .CI(in3[13]), .CO(cout[13]), .S(
        sumout[13]) );
  FADDX1 U6 ( .A(in1[14]), .B(in2[14]), .CI(in3[14]), .CO(cout[14]), .S(
        sumout[14]) );
  FADDX1 U7 ( .A(in1[15]), .B(in2[15]), .CI(in3[15]), .CO(cout[15]), .S(
        sumout[15]) );
  FADDX1 U8 ( .A(in1[16]), .B(in2[16]), .CI(in3[16]), .CO(cout[16]), .S(
        sumout[16]) );
  FADDX1 U9 ( .A(in1[17]), .B(in2[17]), .CI(in3[17]), .CO(cout[17]), .S(
        sumout[17]) );
  FADDX1 U10 ( .A(in1[18]), .B(in2[18]), .CI(in3[18]), .CO(cout[18]), .S(
        sumout[18]) );
  FADDX1 U11 ( .A(in1[19]), .B(in2[19]), .CI(in3[19]), .CO(cout[19]), .S(
        sumout[19]) );
  FADDX1 U12 ( .A(in1[20]), .B(in2[20]), .CI(in3[20]), .CO(cout[20]), .S(
        sumout[20]) );
  FADDX1 U13 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U14 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U15 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U16 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U17 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U18 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U19 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U20 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U21 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U22 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U23 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U24 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
  FADDX1 U25 ( .A(in1[33]), .B(in2[33]), .CI(in3[33]), .CO(cout[33]), .S(
        sumout[33]) );
  FADDX1 U26 ( .A(in1[34]), .B(in2[34]), .CI(in3[34]), .CO(cout[34]), .S(
        sumout[34]) );
  FADDX1 U27 ( .A(in1[35]), .B(in2[35]), .CI(in3[35]), .CO(cout[35]), .S(
        sumout[35]) );
  FADDX1 U28 ( .A(in1[36]), .B(in2[36]), .CI(in3[36]), .CO(cout[36]), .S(
        sumout[36]) );
  FADDX1 U29 ( .A(in1[37]), .B(in2[37]), .CI(in3[37]), .CO(cout[37]), .S(
        sumout[37]) );
  FADDX1 U30 ( .A(in1[38]), .B(in2[38]), .CI(in3[38]), .CO(cout[38]), .S(
        sumout[38]) );
  FADDX1 U31 ( .A(in1[39]), .B(in2[39]), .CI(in3[39]), .CO(cout[39]), .S(
        sumout[39]) );
  FADDX1 U32 ( .A(in1[40]), .B(in2[40]), .CI(in3[40]), .CO(cout[40]), .S(
        sumout[40]) );
  FADDX1 U33 ( .A(in1[41]), .B(in2[41]), .CI(in3[41]), .CO(cout[41]), .S(
        sumout[41]) );
  FADDX1 U34 ( .A(in1[42]), .B(in2[42]), .CI(in3[42]), .CO(cout[42]), .S(
        sumout[42]) );
  FADDX1 U35 ( .A(in1[43]), .B(in2[43]), .CI(in3[43]), .CO(cout[43]), .S(
        sumout[43]) );
  FADDX1 U36 ( .A(in1[44]), .B(in2[44]), .CI(in3[44]), .CO(cout[44]), .S(
        sumout[44]) );
  FADDX1 U37 ( .A(in1[45]), .B(in2[45]), .CI(in3[45]), .CO(cout[45]), .S(
        sumout[45]) );
  FADDX1 U38 ( .A(in1[46]), .B(in2[46]), .CI(in3[46]), .CO(cout[46]), .S(
        sumout[46]) );
  XOR3X1 U39 ( .IN1(in2[47]), .IN2(in3[47]), .IN3(in1[47]), .Q(sumout[47]) );
  FADDX1 U40 ( .A(in1[7]), .B(in2[7]), .CI(in3[7]), .CO(cout[7]), .S(sumout[7]) );
  FADDX1 U41 ( .A(in1[8]), .B(in2[8]), .CI(in3[8]), .CO(cout[8]), .S(sumout[8]) );
  FADDX1 U42 ( .A(in1[9]), .B(in2[9]), .CI(in3[9]), .CO(cout[9]), .S(sumout[9]) );
endmodule


module csa51squ_15 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14;

  AND2X1 U1 ( .IN1(in2[7]), .IN2(in1[7]), .Q(cout[7]) );
  NOR2X0 U2 ( .IN1(in2[7]), .IN2(in1[7]), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(cout[7]), .QN(sumout[7]) );
  AND2X1 U4 ( .IN1(in2[8]), .IN2(in1[8]), .Q(cout[8]) );
  NOR2X0 U5 ( .IN1(in2[8]), .IN2(in1[8]), .QN(n2) );
  NOR2X0 U6 ( .IN1(n2), .IN2(cout[8]), .QN(sumout[8]) );
  AND2X1 U7 ( .IN1(in2[9]), .IN2(in1[9]), .Q(cout[9]) );
  NOR2X0 U8 ( .IN1(in2[9]), .IN2(in1[9]), .QN(n3) );
  NOR2X0 U9 ( .IN1(n3), .IN2(cout[9]), .QN(sumout[9]) );
  AND2X1 U10 ( .IN1(in2[10]), .IN2(in1[10]), .Q(cout[10]) );
  NOR2X0 U11 ( .IN1(in2[10]), .IN2(in1[10]), .QN(n4) );
  NOR2X0 U12 ( .IN1(n4), .IN2(cout[10]), .QN(sumout[10]) );
  AND2X1 U13 ( .IN1(in2[11]), .IN2(in1[11]), .Q(cout[11]) );
  NOR2X0 U14 ( .IN1(in2[11]), .IN2(in1[11]), .QN(n5) );
  NOR2X0 U15 ( .IN1(n5), .IN2(cout[11]), .QN(sumout[11]) );
  AND2X1 U16 ( .IN1(in2[12]), .IN2(in1[12]), .Q(cout[12]) );
  NOR2X0 U17 ( .IN1(in2[12]), .IN2(in1[12]), .QN(n6) );
  NOR2X0 U18 ( .IN1(n6), .IN2(cout[12]), .QN(sumout[12]) );
  AND2X1 U19 ( .IN1(in3[40]), .IN2(in2[40]), .Q(cout[40]) );
  NOR2X0 U20 ( .IN1(in3[40]), .IN2(in2[40]), .QN(n7) );
  NOR2X0 U21 ( .IN1(n7), .IN2(cout[40]), .QN(sumout[40]) );
  AND2X1 U22 ( .IN1(in3[41]), .IN2(in2[41]), .Q(cout[41]) );
  NOR2X0 U23 ( .IN1(in3[41]), .IN2(in2[41]), .QN(n8) );
  NOR2X0 U24 ( .IN1(n8), .IN2(cout[41]), .QN(sumout[41]) );
  AND2X1 U25 ( .IN1(in3[42]), .IN2(in2[42]), .Q(cout[42]) );
  NOR2X0 U26 ( .IN1(in3[42]), .IN2(in2[42]), .QN(n9) );
  NOR2X0 U27 ( .IN1(n9), .IN2(cout[42]), .QN(sumout[42]) );
  AND2X1 U28 ( .IN1(in3[43]), .IN2(in2[43]), .Q(cout[43]) );
  NOR2X0 U29 ( .IN1(in3[43]), .IN2(in2[43]), .QN(n10) );
  NOR2X0 U30 ( .IN1(n10), .IN2(cout[43]), .QN(sumout[43]) );
  AND2X1 U31 ( .IN1(in3[44]), .IN2(in2[44]), .Q(cout[44]) );
  NOR2X0 U32 ( .IN1(in3[44]), .IN2(in2[44]), .QN(n11) );
  NOR2X0 U33 ( .IN1(n11), .IN2(cout[44]), .QN(sumout[44]) );
  AND2X1 U34 ( .IN1(in3[45]), .IN2(in2[45]), .Q(cout[45]) );
  NOR2X0 U35 ( .IN1(in3[45]), .IN2(in2[45]), .QN(n12) );
  NOR2X0 U36 ( .IN1(n12), .IN2(cout[45]), .QN(sumout[45]) );
  AND2X1 U37 ( .IN1(in3[46]), .IN2(in2[46]), .Q(cout[46]) );
  NOR2X0 U38 ( .IN1(in3[46]), .IN2(in2[46]), .QN(n13) );
  NOR2X0 U39 ( .IN1(n13), .IN2(cout[46]), .QN(sumout[46]) );
  INVX0 U40 ( .INP(in3[47]), .ZN(sumout[47]) );
  AND2X1 U41 ( .IN1(in2[5]), .IN2(in1[5]), .Q(cout[5]) );
  AND2X1 U42 ( .IN1(in2[6]), .IN2(in1[6]), .Q(cout[6]) );
  NOR2X0 U43 ( .IN1(in2[6]), .IN2(in1[6]), .QN(n14) );
  NOR2X0 U44 ( .IN1(n14), .IN2(cout[6]), .QN(sumout[6]) );
  FADDX1 U45 ( .A(in1[13]), .B(in2[13]), .CI(in3[13]), .CO(cout[13]), .S(
        sumout[13]) );
  FADDX1 U46 ( .A(in1[14]), .B(in2[14]), .CI(in3[14]), .CO(cout[14]), .S(
        sumout[14]) );
  FADDX1 U47 ( .A(in1[15]), .B(in2[15]), .CI(in3[15]), .CO(cout[15]), .S(
        sumout[15]) );
  FADDX1 U48 ( .A(in1[16]), .B(in2[16]), .CI(in3[16]), .CO(cout[16]), .S(
        sumout[16]) );
  FADDX1 U49 ( .A(in1[17]), .B(in2[17]), .CI(in3[17]), .CO(cout[17]), .S(
        sumout[17]) );
  FADDX1 U50 ( .A(in1[18]), .B(in2[18]), .CI(in3[18]), .CO(cout[18]), .S(
        sumout[18]) );
  FADDX1 U51 ( .A(in1[19]), .B(in2[19]), .CI(in3[19]), .CO(cout[19]), .S(
        sumout[19]) );
  FADDX1 U52 ( .A(in1[20]), .B(in2[20]), .CI(in3[20]), .CO(cout[20]), .S(
        sumout[20]) );
  FADDX1 U53 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U54 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U55 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U56 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U57 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U58 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U59 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U60 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U61 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U62 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U63 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U64 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
  FADDX1 U65 ( .A(in1[33]), .B(in2[33]), .CI(in3[33]), .CO(cout[33]), .S(
        sumout[33]) );
  FADDX1 U66 ( .A(in1[34]), .B(in2[34]), .CI(in3[34]), .CO(cout[34]), .S(
        sumout[34]) );
  FADDX1 U67 ( .A(in1[35]), .B(in2[35]), .CI(in3[35]), .CO(cout[35]), .S(
        sumout[35]) );
  FADDX1 U68 ( .A(in1[36]), .B(in2[36]), .CI(in3[36]), .CO(cout[36]), .S(
        sumout[36]) );
  FADDX1 U69 ( .A(in1[37]), .B(in2[37]), .CI(in3[37]), .CO(cout[37]), .S(
        sumout[37]) );
  FADDX1 U70 ( .A(in1[38]), .B(in2[38]), .CI(in3[38]), .CO(cout[38]), .S(
        sumout[38]) );
  FADDX1 U71 ( .A(in1[39]), .B(in2[39]), .CI(in3[39]), .CO(cout[39]), .S(
        sumout[39]) );
endmodule


module csa51squ_16 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17;

  NBUFFX2 U1 ( .INP(in1[6]), .Z(sumout[6]) );
  NBUFFX2 U2 ( .INP(in1[7]), .Z(sumout[7]) );
  NBUFFX2 U3 ( .INP(in1[8]), .Z(sumout[8]) );
  NBUFFX2 U4 ( .INP(in1[9]), .Z(sumout[9]) );
  NBUFFX2 U5 ( .INP(in1[10]), .Z(sumout[10]) );
  NBUFFX2 U6 ( .INP(in1[11]), .Z(sumout[11]) );
  AND2X1 U7 ( .IN1(in3[13]), .IN2(in1[13]), .Q(cout[13]) );
  NOR2X0 U8 ( .IN1(in3[13]), .IN2(in1[13]), .QN(n7) );
  NOR2X0 U9 ( .IN1(n7), .IN2(cout[13]), .QN(sumout[13]) );
  AND2X1 U10 ( .IN1(in3[15]), .IN2(in1[15]), .Q(cout[15]) );
  NOR2X0 U11 ( .IN1(in3[15]), .IN2(in1[15]), .QN(n8) );
  NOR2X0 U12 ( .IN1(n8), .IN2(cout[15]), .QN(sumout[15]) );
  AND2X1 U13 ( .IN1(in3[17]), .IN2(in1[17]), .Q(cout[17]) );
  NOR2X0 U14 ( .IN1(in3[17]), .IN2(in1[17]), .QN(n9) );
  NOR2X0 U15 ( .IN1(n9), .IN2(cout[17]), .QN(sumout[17]) );
  AND2X1 U16 ( .IN1(in3[43]), .IN2(in2[43]), .Q(cout[43]) );
  NOR2X0 U17 ( .IN1(in3[43]), .IN2(in2[43]), .QN(n10) );
  NOR2X0 U18 ( .IN1(n10), .IN2(cout[43]), .QN(sumout[43]) );
  AND2X1 U19 ( .IN1(in3[44]), .IN2(in2[44]), .Q(cout[44]) );
  NOR2X0 U20 ( .IN1(in3[44]), .IN2(in2[44]), .QN(n11) );
  NOR2X0 U21 ( .IN1(n11), .IN2(cout[44]), .QN(sumout[44]) );
  AND2X1 U22 ( .IN1(in3[45]), .IN2(in2[45]), .Q(cout[45]) );
  NOR2X0 U23 ( .IN1(in3[45]), .IN2(in2[45]), .QN(n12) );
  NOR2X0 U24 ( .IN1(n12), .IN2(cout[45]), .QN(sumout[45]) );
  AND2X1 U25 ( .IN1(in3[46]), .IN2(in2[46]), .Q(cout[46]) );
  NOR2X0 U26 ( .IN1(in3[46]), .IN2(in2[46]), .QN(n13) );
  NOR2X0 U27 ( .IN1(n13), .IN2(cout[46]), .QN(sumout[46]) );
  XOR2X1 U28 ( .IN1(in3[47]), .IN2(in2[47]), .Q(sumout[47]) );
  AND2X1 U29 ( .IN1(in3[12]), .IN2(in1[12]), .Q(cout[12]) );
  NOR2X0 U30 ( .IN1(in3[12]), .IN2(in1[12]), .QN(n14) );
  NOR2X0 U31 ( .IN1(n14), .IN2(cout[12]), .QN(sumout[12]) );
  AND2X1 U32 ( .IN1(in3[14]), .IN2(in1[14]), .Q(cout[14]) );
  NOR2X0 U33 ( .IN1(in3[14]), .IN2(in1[14]), .QN(n15) );
  NOR2X0 U34 ( .IN1(n15), .IN2(cout[14]), .QN(sumout[14]) );
  AND2X1 U35 ( .IN1(in3[16]), .IN2(in1[16]), .Q(cout[16]) );
  NOR2X0 U36 ( .IN1(in3[16]), .IN2(in1[16]), .QN(n16) );
  NOR2X0 U37 ( .IN1(n16), .IN2(cout[16]), .QN(sumout[16]) );
  AND2X1 U38 ( .IN1(in3[18]), .IN2(in1[18]), .Q(cout[18]) );
  NOR2X0 U39 ( .IN1(in3[18]), .IN2(in1[18]), .QN(n17) );
  NOR2X0 U40 ( .IN1(n17), .IN2(cout[18]), .QN(sumout[18]) );
  FADDX1 U41 ( .A(in1[19]), .B(in2[19]), .CI(in3[19]), .CO(cout[19]), .S(
        sumout[19]) );
  FADDX1 U42 ( .A(in1[20]), .B(in2[20]), .CI(in3[20]), .CO(cout[20]), .S(
        sumout[20]) );
  FADDX1 U43 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U44 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U45 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U46 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U47 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U48 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U49 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U50 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U51 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U52 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U53 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U54 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
  FADDX1 U55 ( .A(in1[33]), .B(in2[33]), .CI(in3[33]), .CO(cout[33]), .S(
        sumout[33]) );
  FADDX1 U56 ( .A(in1[34]), .B(in2[34]), .CI(in3[34]), .CO(cout[34]), .S(
        sumout[34]) );
  FADDX1 U57 ( .A(in1[35]), .B(in2[35]), .CI(in3[35]), .CO(cout[35]), .S(
        sumout[35]) );
  FADDX1 U58 ( .A(in1[36]), .B(in2[36]), .CI(in3[36]), .CO(cout[36]), .S(
        sumout[36]) );
  FADDX1 U59 ( .A(in1[37]), .B(in2[37]), .CI(in3[37]), .CO(cout[37]), .S(
        sumout[37]) );
  FADDX1 U60 ( .A(in1[38]), .B(in2[38]), .CI(in3[38]), .CO(cout[38]), .S(
        sumout[38]) );
  FADDX1 U61 ( .A(in1[39]), .B(in2[39]), .CI(in3[39]), .CO(cout[39]), .S(
        sumout[39]) );
  FADDX1 U62 ( .A(in1[40]), .B(in2[40]), .CI(in3[40]), .CO(cout[40]), .S(
        sumout[40]) );
  FADDX1 U63 ( .A(in1[41]), .B(in2[41]), .CI(in3[41]), .CO(cout[41]), .S(
        sumout[41]) );
  FADDX1 U64 ( .A(in1[42]), .B(in2[42]), .CI(in3[42]), .CO(cout[42]), .S(
        sumout[42]) );
endmodule


module csa51squ_17 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19;

  NBUFFX2 U1 ( .INP(in2[46]), .Z(sumout[46]) );
  NBUFFX2 U2 ( .INP(in2[45]), .Z(sumout[45]) );
  NBUFFX2 U3 ( .INP(in2[44]), .Z(sumout[44]) );
  NBUFFX2 U4 ( .INP(in2[43]), .Z(sumout[43]) );
  NBUFFX2 U5 ( .INP(in2[42]), .Z(sumout[42]) );
  NBUFFX2 U6 ( .INP(in2[41]), .Z(sumout[41]) );
  NBUFFX2 U7 ( .INP(in2[40]), .Z(sumout[40]) );
  NBUFFX2 U8 ( .INP(in2[39]), .Z(sumout[39]) );
  AND2X1 U9 ( .IN1(in2[7]), .IN2(in1[7]), .Q(cout[7]) );
  NOR2X0 U10 ( .IN1(in2[7]), .IN2(in1[7]), .QN(n9) );
  NOR2X0 U11 ( .IN1(n9), .IN2(cout[7]), .QN(sumout[7]) );
  AND2X1 U12 ( .IN1(in2[8]), .IN2(in1[8]), .Q(cout[8]) );
  NOR2X0 U13 ( .IN1(in2[8]), .IN2(in1[8]), .QN(n10) );
  NOR2X0 U14 ( .IN1(n10), .IN2(cout[8]), .QN(sumout[8]) );
  AND2X1 U15 ( .IN1(in2[9]), .IN2(in1[9]), .Q(cout[9]) );
  NOR2X0 U16 ( .IN1(in2[9]), .IN2(in1[9]), .QN(n11) );
  NOR2X0 U17 ( .IN1(n11), .IN2(cout[9]), .QN(sumout[9]) );
  AND2X1 U18 ( .IN1(in3[33]), .IN2(in2[33]), .Q(cout[33]) );
  NOR2X0 U19 ( .IN1(in3[33]), .IN2(in2[33]), .QN(n12) );
  NOR2X0 U20 ( .IN1(n12), .IN2(cout[33]), .QN(sumout[33]) );
  AND2X1 U21 ( .IN1(in3[34]), .IN2(in2[34]), .Q(cout[34]) );
  NOR2X0 U22 ( .IN1(in3[34]), .IN2(in2[34]), .QN(n13) );
  NOR2X0 U23 ( .IN1(n13), .IN2(cout[34]), .QN(sumout[34]) );
  AND2X1 U24 ( .IN1(in3[35]), .IN2(in2[35]), .Q(cout[35]) );
  NOR2X0 U25 ( .IN1(in3[35]), .IN2(in2[35]), .QN(n14) );
  NOR2X0 U26 ( .IN1(n14), .IN2(cout[35]), .QN(sumout[35]) );
  AND2X1 U27 ( .IN1(in3[36]), .IN2(in2[36]), .Q(cout[36]) );
  NOR2X0 U28 ( .IN1(in3[36]), .IN2(in2[36]), .QN(n15) );
  NOR2X0 U29 ( .IN1(n15), .IN2(cout[36]), .QN(sumout[36]) );
  AND2X1 U30 ( .IN1(in3[37]), .IN2(in2[37]), .Q(cout[37]) );
  NOR2X0 U31 ( .IN1(in3[37]), .IN2(in2[37]), .QN(n16) );
  NOR2X0 U32 ( .IN1(n16), .IN2(cout[37]), .QN(sumout[37]) );
  AND2X1 U33 ( .IN1(in3[38]), .IN2(in2[38]), .Q(cout[38]) );
  NOR2X0 U34 ( .IN1(in3[38]), .IN2(in2[38]), .QN(n17) );
  NOR2X0 U35 ( .IN1(n17), .IN2(cout[38]), .QN(sumout[38]) );
  AND2X1 U36 ( .IN1(in2[4]), .IN2(in1[4]), .Q(cout[4]) );
  AND2X1 U37 ( .IN1(in2[5]), .IN2(in1[5]), .Q(cout[5]) );
  NOR2X0 U38 ( .IN1(in2[5]), .IN2(in1[5]), .QN(n18) );
  NOR2X0 U39 ( .IN1(n18), .IN2(cout[5]), .QN(sumout[5]) );
  AND2X1 U40 ( .IN1(in2[6]), .IN2(in1[6]), .Q(cout[6]) );
  NOR2X0 U41 ( .IN1(in2[6]), .IN2(in1[6]), .QN(n19) );
  NOR2X0 U42 ( .IN1(n19), .IN2(cout[6]), .QN(sumout[6]) );
  FADDX1 U43 ( .A(in1[10]), .B(in2[10]), .CI(in3[10]), .CO(cout[10]), .S(
        sumout[10]) );
  FADDX1 U44 ( .A(in1[11]), .B(in2[11]), .CI(in3[11]), .CO(cout[11]), .S(
        sumout[11]) );
  FADDX1 U45 ( .A(in1[12]), .B(in2[12]), .CI(in3[12]), .CO(cout[12]), .S(
        sumout[12]) );
  FADDX1 U46 ( .A(in1[13]), .B(in2[13]), .CI(in3[13]), .CO(cout[13]), .S(
        sumout[13]) );
  FADDX1 U47 ( .A(in1[14]), .B(in2[14]), .CI(in3[14]), .CO(cout[14]), .S(
        sumout[14]) );
  FADDX1 U48 ( .A(in1[15]), .B(in2[15]), .CI(in3[15]), .CO(cout[15]), .S(
        sumout[15]) );
  FADDX1 U49 ( .A(in1[16]), .B(in2[16]), .CI(in3[16]), .CO(cout[16]), .S(
        sumout[16]) );
  FADDX1 U50 ( .A(in1[17]), .B(in2[17]), .CI(in3[17]), .CO(cout[17]), .S(
        sumout[17]) );
  FADDX1 U51 ( .A(in1[18]), .B(in2[18]), .CI(in3[18]), .CO(cout[18]), .S(
        sumout[18]) );
  FADDX1 U52 ( .A(in1[19]), .B(in2[19]), .CI(in3[19]), .CO(cout[19]), .S(
        sumout[19]) );
  FADDX1 U53 ( .A(in1[20]), .B(in2[20]), .CI(in3[20]), .CO(cout[20]), .S(
        sumout[20]) );
  FADDX1 U54 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U55 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U56 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U57 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U58 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U59 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U60 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U61 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U62 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U63 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U64 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U65 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
endmodule


module csa51squ_18 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n7, n8, n9, n10, n11, n12, n13;

  NBUFFX2 U1 ( .INP(in1[12]), .Z(sumout[12]) );
  NBUFFX2 U2 ( .INP(in1[13]), .Z(sumout[13]) );
  NBUFFX2 U3 ( .INP(in1[14]), .Z(sumout[14]) );
  NBUFFX2 U4 ( .INP(in1[15]), .Z(sumout[15]) );
  NBUFFX2 U5 ( .INP(in1[16]), .Z(sumout[16]) );
  NBUFFX2 U6 ( .INP(in1[17]), .Z(sumout[17]) );
  AND2X1 U7 ( .IN1(in3[19]), .IN2(in1[19]), .Q(cout[19]) );
  NOR2X0 U8 ( .IN1(in3[19]), .IN2(in1[19]), .QN(n7) );
  NOR2X0 U9 ( .IN1(n7), .IN2(cout[19]), .QN(sumout[19]) );
  AND2X1 U10 ( .IN1(in3[44]), .IN2(in2[44]), .Q(cout[44]) );
  NOR2X0 U11 ( .IN1(in3[44]), .IN2(in2[44]), .QN(n8) );
  NOR2X0 U12 ( .IN1(n8), .IN2(cout[44]), .QN(sumout[44]) );
  AND2X1 U13 ( .IN1(in3[45]), .IN2(in2[45]), .Q(cout[45]) );
  NOR2X0 U14 ( .IN1(in3[45]), .IN2(in2[45]), .QN(n9) );
  NOR2X0 U15 ( .IN1(n9), .IN2(cout[45]), .QN(sumout[45]) );
  AND2X1 U16 ( .IN1(in3[46]), .IN2(in2[46]), .Q(cout[46]) );
  NOR2X0 U17 ( .IN1(in3[46]), .IN2(in2[46]), .QN(n10) );
  NOR2X0 U18 ( .IN1(n10), .IN2(cout[46]), .QN(sumout[46]) );
  XOR2X1 U19 ( .IN1(in3[47]), .IN2(in2[47]), .Q(sumout[47]) );
  AND2X1 U20 ( .IN1(in3[18]), .IN2(in1[18]), .Q(cout[18]) );
  NOR2X0 U21 ( .IN1(in3[18]), .IN2(in1[18]), .QN(n11) );
  NOR2X0 U22 ( .IN1(n11), .IN2(cout[18]), .QN(sumout[18]) );
  AND2X1 U23 ( .IN1(in3[20]), .IN2(in1[20]), .Q(cout[20]) );
  NOR2X0 U24 ( .IN1(in3[20]), .IN2(in1[20]), .QN(n12) );
  NOR2X0 U25 ( .IN1(n12), .IN2(cout[20]), .QN(sumout[20]) );
  INVX0 U26 ( .INP(in1[42]), .ZN(n13) );
  FADDX1 U27 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U28 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U29 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U30 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U31 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U32 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U33 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U34 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U35 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U36 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U37 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U38 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
  FADDX1 U39 ( .A(in1[33]), .B(in2[33]), .CI(in3[33]), .CO(cout[33]), .S(
        sumout[33]) );
  FADDX1 U40 ( .A(in1[34]), .B(in2[34]), .CI(in3[34]), .CO(cout[34]), .S(
        sumout[34]) );
  FADDX1 U41 ( .A(in1[35]), .B(in2[35]), .CI(in3[35]), .CO(cout[35]), .S(
        sumout[35]) );
  FADDX1 U42 ( .A(in1[36]), .B(in2[36]), .CI(in3[36]), .CO(cout[36]), .S(
        sumout[36]) );
  FADDX1 U43 ( .A(in1[37]), .B(in2[37]), .CI(in3[37]), .CO(cout[37]), .S(
        sumout[37]) );
  FADDX1 U44 ( .A(in1[38]), .B(in2[38]), .CI(in3[38]), .CO(cout[38]), .S(
        sumout[38]) );
  FADDX1 U45 ( .A(in1[39]), .B(in2[39]), .CI(in3[39]), .CO(cout[39]), .S(
        sumout[39]) );
  FADDX1 U46 ( .A(in1[40]), .B(in2[40]), .CI(in3[40]), .CO(cout[40]), .S(
        sumout[40]) );
  FADDX1 U47 ( .A(in1[41]), .B(in2[41]), .CI(in3[41]), .CO(cout[41]), .S(
        sumout[41]) );
  FADDX1 U48 ( .A(in1[42]), .B(in2[42]), .CI(in3[42]), .CO(cout[42]), .S(
        sumout[42]) );
  FADDX1 U49 ( .A(in2[43]), .B(in3[43]), .CI(n13), .CO(cout[43]), .S(
        sumout[43]) );
endmodule


module csa51squ_19 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n9, n10, n11, n12, n13, n14, n15;

  NBUFFX2 U1 ( .INP(in2[6]), .Z(sumout[6]) );
  NBUFFX2 U2 ( .INP(in2[7]), .Z(sumout[7]) );
  NBUFFX2 U3 ( .INP(in2[8]), .Z(sumout[8]) );
  NBUFFX2 U4 ( .INP(in3[42]), .Z(sumout[42]) );
  NBUFFX2 U5 ( .INP(in3[41]), .Z(sumout[41]) );
  NBUFFX2 U6 ( .INP(in3[39]), .Z(sumout[39]) );
  NBUFFX2 U7 ( .INP(in3[38]), .Z(sumout[38]) );
  NBUFFX2 U8 ( .INP(in3[40]), .Z(sumout[40]) );
  AND2X1 U9 ( .IN1(in2[13]), .IN2(in1[13]), .Q(cout[13]) );
  NOR2X0 U10 ( .IN1(in2[13]), .IN2(in1[13]), .QN(n9) );
  NOR2X0 U11 ( .IN1(n9), .IN2(cout[13]), .QN(sumout[13]) );
  AND2X1 U12 ( .IN1(in2[37]), .IN2(in3[37]), .Q(cout[37]) );
  INVX0 U13 ( .INP(in2[37]), .ZN(n15) );
  MUX21X1 U14 ( .IN1(in2[37]), .IN2(n15), .S(in3[37]), .Q(sumout[37]) );
  AND2X1 U15 ( .IN1(in2[9]), .IN2(in1[9]), .Q(cout[9]) );
  NOR2X0 U16 ( .IN1(in2[9]), .IN2(in1[9]), .QN(n10) );
  NOR2X0 U17 ( .IN1(n10), .IN2(cout[9]), .QN(sumout[9]) );
  AND2X1 U18 ( .IN1(in2[10]), .IN2(in1[10]), .Q(cout[10]) );
  NOR2X0 U19 ( .IN1(in2[10]), .IN2(in1[10]), .QN(n11) );
  NOR2X0 U20 ( .IN1(n11), .IN2(cout[10]), .QN(sumout[10]) );
  AND2X1 U21 ( .IN1(in2[11]), .IN2(in1[11]), .Q(cout[11]) );
  NOR2X0 U22 ( .IN1(in2[11]), .IN2(in1[11]), .QN(n12) );
  NOR2X0 U23 ( .IN1(n12), .IN2(cout[11]), .QN(sumout[11]) );
  AND2X1 U24 ( .IN1(in2[12]), .IN2(in1[12]), .Q(cout[12]) );
  NOR2X0 U25 ( .IN1(in2[12]), .IN2(in1[12]), .QN(n13) );
  NOR2X0 U26 ( .IN1(n13), .IN2(cout[12]), .QN(sumout[12]) );
  AND2X1 U27 ( .IN1(in2[14]), .IN2(in1[14]), .Q(cout[14]) );
  NOR2X0 U28 ( .IN1(in2[14]), .IN2(in1[14]), .QN(n14) );
  NOR2X0 U29 ( .IN1(n14), .IN2(cout[14]), .QN(sumout[14]) );
  FADDX1 U30 ( .A(in1[15]), .B(in2[15]), .CI(in3[15]), .CO(cout[15]), .S(
        sumout[15]) );
  FADDX1 U31 ( .A(in1[16]), .B(in2[16]), .CI(in3[16]), .CO(cout[16]), .S(
        sumout[16]) );
  FADDX1 U32 ( .A(in1[17]), .B(in2[17]), .CI(in3[17]), .CO(cout[17]), .S(
        sumout[17]) );
  FADDX1 U33 ( .A(in1[18]), .B(in2[18]), .CI(in3[18]), .CO(cout[18]), .S(
        sumout[18]) );
  FADDX1 U34 ( .A(in1[19]), .B(in2[19]), .CI(in3[19]), .CO(cout[19]), .S(
        sumout[19]) );
  FADDX1 U35 ( .A(in1[20]), .B(in2[20]), .CI(in3[20]), .CO(cout[20]), .S(
        sumout[20]) );
  FADDX1 U36 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U37 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U38 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U39 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U40 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U41 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U42 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U43 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U44 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U45 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U46 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U47 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
  FADDX1 U48 ( .A(in1[33]), .B(in2[33]), .CI(in3[33]), .CO(cout[33]), .S(
        sumout[33]) );
  FADDX1 U49 ( .A(in1[34]), .B(in2[34]), .CI(in3[34]), .CO(cout[34]), .S(
        sumout[34]) );
  FADDX1 U50 ( .A(in1[35]), .B(in2[35]), .CI(in3[35]), .CO(cout[35]), .S(
        sumout[35]) );
  FADDX1 U51 ( .A(in1[36]), .B(in3[36]), .CI(n15), .CO(cout[36]), .S(
        sumout[36]) );
endmodule


module csa51squ_20 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36;

  NBUFFX2 U1 ( .INP(in3[46]), .Z(sumout[46]) );
  NBUFFX2 U2 ( .INP(in3[45]), .Z(sumout[45]) );
  NBUFFX2 U3 ( .INP(in3[44]), .Z(sumout[44]) );
  NBUFFX2 U4 ( .INP(in3[43]), .Z(sumout[43]) );
  NBUFFX2 U5 ( .INP(in3[42]), .Z(sumout[42]) );
  NBUFFX2 U6 ( .INP(in3[33]), .Z(sumout[33]) );
  NBUFFX2 U7 ( .INP(in3[32]), .Z(sumout[32]) );
  NBUFFX2 U8 ( .INP(in3[35]), .Z(sumout[35]) );
  NBUFFX2 U9 ( .INP(in3[34]), .Z(sumout[34]) );
  NBUFFX2 U10 ( .INP(in3[37]), .Z(sumout[37]) );
  NBUFFX2 U11 ( .INP(in3[36]), .Z(sumout[36]) );
  NBUFFX2 U12 ( .INP(in3[41]), .Z(sumout[41]) );
  NBUFFX2 U13 ( .INP(in3[40]), .Z(sumout[40]) );
  NBUFFX2 U14 ( .INP(in3[39]), .Z(sumout[39]) );
  NBUFFX2 U15 ( .INP(in3[38]), .Z(sumout[38]) );
  AND2X1 U16 ( .IN1(in2[31]), .IN2(in3[31]), .Q(cout[31]) );
  INVX0 U17 ( .INP(in2[31]), .ZN(n36) );
  MUX21X1 U18 ( .IN1(in2[31]), .IN2(n36), .S(in3[31]), .Q(sumout[31]) );
  AND2X1 U19 ( .IN1(in2[3]), .IN2(in1[3]), .Q(cout[3]) );
  AND2X1 U20 ( .IN1(in2[4]), .IN2(in1[4]), .Q(cout[4]) );
  NOR2X0 U21 ( .IN1(in2[4]), .IN2(in1[4]), .QN(n16) );
  NOR2X0 U22 ( .IN1(n16), .IN2(cout[4]), .QN(sumout[4]) );
  AND2X1 U23 ( .IN1(in2[5]), .IN2(in1[5]), .Q(cout[5]) );
  NOR2X0 U24 ( .IN1(in2[5]), .IN2(in1[5]), .QN(n17) );
  NOR2X0 U25 ( .IN1(n17), .IN2(cout[5]), .QN(sumout[5]) );
  AND2X1 U26 ( .IN1(in2[6]), .IN2(in1[6]), .Q(cout[6]) );
  NOR2X0 U27 ( .IN1(in2[6]), .IN2(in1[6]), .QN(n18) );
  NOR2X0 U28 ( .IN1(n18), .IN2(cout[6]), .QN(sumout[6]) );
  AND2X1 U29 ( .IN1(in2[7]), .IN2(in1[7]), .Q(cout[7]) );
  NOR2X0 U30 ( .IN1(in2[7]), .IN2(in1[7]), .QN(n19) );
  NOR2X0 U31 ( .IN1(n19), .IN2(cout[7]), .QN(sumout[7]) );
  AND2X1 U32 ( .IN1(in2[8]), .IN2(in1[8]), .Q(cout[8]) );
  NOR2X0 U33 ( .IN1(in2[8]), .IN2(in1[8]), .QN(n20) );
  NOR2X0 U34 ( .IN1(n20), .IN2(cout[8]), .QN(sumout[8]) );
  AND2X1 U35 ( .IN1(in2[9]), .IN2(in1[9]), .Q(cout[9]) );
  NOR2X0 U36 ( .IN1(in2[9]), .IN2(in1[9]), .QN(n21) );
  NOR2X0 U37 ( .IN1(n21), .IN2(cout[9]), .QN(sumout[9]) );
  AND2X1 U38 ( .IN1(in2[10]), .IN2(in1[10]), .Q(cout[10]) );
  NOR2X0 U39 ( .IN1(in2[10]), .IN2(in1[10]), .QN(n22) );
  NOR2X0 U40 ( .IN1(n22), .IN2(cout[10]), .QN(sumout[10]) );
  AND2X1 U41 ( .IN1(in2[11]), .IN2(in1[11]), .Q(cout[11]) );
  NOR2X0 U42 ( .IN1(in2[11]), .IN2(in1[11]), .QN(n23) );
  NOR2X0 U43 ( .IN1(n23), .IN2(cout[11]), .QN(sumout[11]) );
  AND2X1 U44 ( .IN1(in2[12]), .IN2(in1[12]), .Q(cout[12]) );
  NOR2X0 U45 ( .IN1(in2[12]), .IN2(in1[12]), .QN(n24) );
  NOR2X0 U46 ( .IN1(n24), .IN2(cout[12]), .QN(sumout[12]) );
  AND2X1 U47 ( .IN1(in2[13]), .IN2(in1[13]), .Q(cout[13]) );
  NOR2X0 U48 ( .IN1(in2[13]), .IN2(in1[13]), .QN(n25) );
  NOR2X0 U49 ( .IN1(n25), .IN2(cout[13]), .QN(sumout[13]) );
  AND2X1 U50 ( .IN1(in2[14]), .IN2(in1[14]), .Q(cout[14]) );
  NOR2X0 U51 ( .IN1(in2[14]), .IN2(in1[14]), .QN(n26) );
  NOR2X0 U52 ( .IN1(n26), .IN2(cout[14]), .QN(sumout[14]) );
  AND2X1 U53 ( .IN1(in2[15]), .IN2(in1[15]), .Q(cout[15]) );
  NOR2X0 U54 ( .IN1(in2[15]), .IN2(in1[15]), .QN(n27) );
  NOR2X0 U55 ( .IN1(n27), .IN2(cout[15]), .QN(sumout[15]) );
  AND2X1 U56 ( .IN1(in2[16]), .IN2(in1[16]), .Q(cout[16]) );
  NOR2X0 U57 ( .IN1(in2[16]), .IN2(in1[16]), .QN(n28) );
  NOR2X0 U58 ( .IN1(n28), .IN2(cout[16]), .QN(sumout[16]) );
  AND2X1 U59 ( .IN1(in2[17]), .IN2(in1[17]), .Q(cout[17]) );
  NOR2X0 U60 ( .IN1(in2[17]), .IN2(in1[17]), .QN(n29) );
  NOR2X0 U61 ( .IN1(n29), .IN2(cout[17]), .QN(sumout[17]) );
  AND2X1 U62 ( .IN1(in2[18]), .IN2(in1[18]), .Q(cout[18]) );
  NOR2X0 U63 ( .IN1(in2[18]), .IN2(in1[18]), .QN(n30) );
  NOR2X0 U64 ( .IN1(n30), .IN2(cout[18]), .QN(sumout[18]) );
  AND2X1 U65 ( .IN1(in2[19]), .IN2(in1[19]), .Q(cout[19]) );
  NOR2X0 U66 ( .IN1(in2[19]), .IN2(in1[19]), .QN(n31) );
  NOR2X0 U67 ( .IN1(n31), .IN2(cout[19]), .QN(sumout[19]) );
  AND2X1 U68 ( .IN1(in2[20]), .IN2(in1[20]), .Q(cout[20]) );
  NOR2X0 U69 ( .IN1(in2[20]), .IN2(in1[20]), .QN(n32) );
  NOR2X0 U70 ( .IN1(n32), .IN2(cout[20]), .QN(sumout[20]) );
  AND2X1 U71 ( .IN1(in2[21]), .IN2(in1[21]), .Q(cout[21]) );
  NOR2X0 U72 ( .IN1(in2[21]), .IN2(in1[21]), .QN(n33) );
  NOR2X0 U73 ( .IN1(n33), .IN2(cout[21]), .QN(sumout[21]) );
  AND2X1 U74 ( .IN1(in2[22]), .IN2(in1[22]), .Q(cout[22]) );
  NOR2X0 U75 ( .IN1(in2[22]), .IN2(in1[22]), .QN(n34) );
  NOR2X0 U76 ( .IN1(n34), .IN2(cout[22]), .QN(sumout[22]) );
  AND2X1 U77 ( .IN1(in2[23]), .IN2(in1[23]), .Q(cout[23]) );
  NOR2X0 U78 ( .IN1(in2[23]), .IN2(in1[23]), .QN(n35) );
  NOR2X0 U79 ( .IN1(n35), .IN2(cout[23]), .QN(sumout[23]) );
  FADDX1 U80 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U81 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U82 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U83 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U84 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U85 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U86 ( .A(in1[30]), .B(in3[30]), .CI(n36), .CO(cout[30]), .S(
        sumout[30]) );
endmodule


module csa51squ_21 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n3, n4, n5, n6, n7;

  NBUFFX2 U1 ( .INP(in1[18]), .Z(sumout[18]) );
  NBUFFX2 U2 ( .INP(in1[19]), .Z(sumout[19]) );
  AND2X1 U3 ( .IN1(in2[20]), .IN2(in1[20]), .Q(cout[20]) );
  NOR2X0 U4 ( .IN1(in2[20]), .IN2(in1[20]), .QN(n3) );
  NOR2X0 U5 ( .IN1(n3), .IN2(cout[20]), .QN(sumout[20]) );
  AND2X1 U6 ( .IN1(in2[21]), .IN2(in1[21]), .Q(cout[21]) );
  NOR2X0 U7 ( .IN1(in2[21]), .IN2(in1[21]), .QN(n4) );
  NOR2X0 U8 ( .IN1(n4), .IN2(cout[21]), .QN(sumout[21]) );
  AND2X1 U9 ( .IN1(in2[46]), .IN2(in3[46]), .Q(cout[46]) );
  NOR2X0 U10 ( .IN1(in2[46]), .IN2(in3[46]), .QN(n5) );
  NOR2X0 U11 ( .IN1(n5), .IN2(cout[46]), .QN(sumout[46]) );
  INVX0 U12 ( .INP(in2[46]), .ZN(n6) );
  MUX21X1 U13 ( .IN1(n6), .IN2(in2[46]), .S(in3[47]), .Q(sumout[47]) );
  INVX0 U14 ( .INP(in1[44]), .ZN(n7) );
  FADDX1 U15 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U16 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U17 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U18 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U19 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U20 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U21 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U22 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U23 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U24 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U25 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
  FADDX1 U26 ( .A(in1[33]), .B(in2[33]), .CI(in3[33]), .CO(cout[33]), .S(
        sumout[33]) );
  FADDX1 U27 ( .A(in1[34]), .B(in2[34]), .CI(in3[34]), .CO(cout[34]), .S(
        sumout[34]) );
  FADDX1 U28 ( .A(in1[35]), .B(in2[35]), .CI(in3[35]), .CO(cout[35]), .S(
        sumout[35]) );
  FADDX1 U29 ( .A(in1[36]), .B(in2[36]), .CI(in3[36]), .CO(cout[36]), .S(
        sumout[36]) );
  FADDX1 U30 ( .A(in1[37]), .B(in2[37]), .CI(in3[37]), .CO(cout[37]), .S(
        sumout[37]) );
  FADDX1 U31 ( .A(in1[38]), .B(in2[38]), .CI(in3[38]), .CO(cout[38]), .S(
        sumout[38]) );
  FADDX1 U32 ( .A(in1[39]), .B(in2[39]), .CI(in3[39]), .CO(cout[39]), .S(
        sumout[39]) );
  FADDX1 U33 ( .A(in1[40]), .B(in2[40]), .CI(in3[40]), .CO(cout[40]), .S(
        sumout[40]) );
  FADDX1 U34 ( .A(in1[41]), .B(in2[41]), .CI(in3[41]), .CO(cout[41]), .S(
        sumout[41]) );
  FADDX1 U35 ( .A(in1[42]), .B(in2[42]), .CI(in3[42]), .CO(cout[42]), .S(
        sumout[42]) );
  FADDX1 U36 ( .A(in1[43]), .B(in2[43]), .CI(in3[43]), .CO(cout[43]), .S(
        sumout[43]) );
  FADDX1 U37 ( .A(in1[44]), .B(in2[44]), .CI(in3[44]), .CO(cout[44]), .S(
        sumout[44]) );
  FADDX1 U38 ( .A(in2[45]), .B(in3[45]), .CI(n7), .CO(cout[45]), .S(sumout[45]) );
endmodule


module csa51squ_22 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n4, n5, n6, n7, n8;

  NBUFFX2 U1 ( .INP(in1[12]), .Z(sumout[12]) );
  NBUFFX2 U2 ( .INP(in1[13]), .Z(sumout[13]) );
  NBUFFX2 U3 ( .INP(in3[42]), .Z(sumout[42]) );
  AND2X1 U4 ( .IN1(in2[14]), .IN2(in1[14]), .Q(cout[14]) );
  NOR2X0 U5 ( .IN1(in2[14]), .IN2(in1[14]), .QN(n4) );
  NOR2X0 U6 ( .IN1(n4), .IN2(cout[14]), .QN(sumout[14]) );
  AND2X1 U7 ( .IN1(in2[15]), .IN2(in1[15]), .Q(cout[15]) );
  NOR2X0 U8 ( .IN1(in2[15]), .IN2(in1[15]), .QN(n5) );
  NOR2X0 U9 ( .IN1(n5), .IN2(cout[15]), .QN(sumout[15]) );
  AND2X1 U10 ( .IN1(in2[40]), .IN2(in3[40]), .Q(cout[40]) );
  NOR2X0 U11 ( .IN1(in2[40]), .IN2(in3[40]), .QN(n6) );
  NOR2X0 U12 ( .IN1(n6), .IN2(cout[40]), .QN(sumout[40]) );
  INVX0 U13 ( .INP(in3[41]), .ZN(n7) );
  NOR2X0 U14 ( .IN1(in2[40]), .IN2(n7), .QN(cout[41]) );
  MUX21X1 U15 ( .IN1(n7), .IN2(in3[41]), .S(in2[40]), .Q(sumout[41]) );
  INVX0 U16 ( .INP(in1[38]), .ZN(n8) );
  FADDX1 U17 ( .A(in1[16]), .B(in2[16]), .CI(in3[16]), .CO(cout[16]), .S(
        sumout[16]) );
  FADDX1 U18 ( .A(in1[17]), .B(in2[17]), .CI(in3[17]), .CO(cout[17]), .S(
        sumout[17]) );
  FADDX1 U19 ( .A(in1[18]), .B(in2[18]), .CI(in3[18]), .CO(cout[18]), .S(
        sumout[18]) );
  FADDX1 U20 ( .A(in1[19]), .B(in2[19]), .CI(in3[19]), .CO(cout[19]), .S(
        sumout[19]) );
  FADDX1 U21 ( .A(in1[20]), .B(in2[20]), .CI(in3[20]), .CO(cout[20]), .S(
        sumout[20]) );
  FADDX1 U22 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U23 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U24 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U25 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U26 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U27 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U28 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U29 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U30 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U31 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U32 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U33 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
  FADDX1 U34 ( .A(in1[33]), .B(in2[33]), .CI(in3[33]), .CO(cout[33]), .S(
        sumout[33]) );
  FADDX1 U35 ( .A(in1[34]), .B(in2[34]), .CI(in3[34]), .CO(cout[34]), .S(
        sumout[34]) );
  FADDX1 U36 ( .A(in1[35]), .B(in2[35]), .CI(in3[35]), .CO(cout[35]), .S(
        sumout[35]) );
  FADDX1 U37 ( .A(in1[36]), .B(in2[36]), .CI(in3[36]), .CO(cout[36]), .S(
        sumout[36]) );
  FADDX1 U38 ( .A(in1[37]), .B(in2[37]), .CI(in3[37]), .CO(cout[37]), .S(
        sumout[37]) );
  FADDX1 U39 ( .A(in1[38]), .B(in2[38]), .CI(in3[38]), .CO(cout[38]), .S(
        sumout[38]) );
  FADDX1 U40 ( .A(in2[39]), .B(in3[39]), .CI(n8), .CO(cout[39]), .S(sumout[39]) );
endmodule


module csa51squ_23 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n4, n5, n6, n7, n8;

  NBUFFX2 U1 ( .INP(in1[6]), .Z(sumout[6]) );
  NBUFFX2 U2 ( .INP(in1[7]), .Z(sumout[7]) );
  NBUFFX2 U3 ( .INP(in3[37]), .Z(sumout[37]) );
  AND2X1 U4 ( .IN1(in2[8]), .IN2(in1[8]), .Q(cout[8]) );
  NOR2X0 U5 ( .IN1(in2[8]), .IN2(in1[8]), .QN(n4) );
  NOR2X0 U6 ( .IN1(n4), .IN2(cout[8]), .QN(sumout[8]) );
  AND2X1 U7 ( .IN1(in2[9]), .IN2(in1[9]), .Q(cout[9]) );
  NOR2X0 U8 ( .IN1(in2[9]), .IN2(in1[9]), .QN(n5) );
  NOR2X0 U9 ( .IN1(n5), .IN2(cout[9]), .QN(sumout[9]) );
  AND2X1 U10 ( .IN1(in2[34]), .IN2(in3[34]), .Q(cout[34]) );
  NOR2X0 U11 ( .IN1(in2[34]), .IN2(in3[34]), .QN(n6) );
  NOR2X0 U12 ( .IN1(n6), .IN2(cout[34]), .QN(sumout[34]) );
  INVX0 U13 ( .INP(in3[35]), .ZN(n7) );
  NOR2X0 U14 ( .IN1(in2[34]), .IN2(n7), .QN(cout[35]) );
  MUX21X1 U15 ( .IN1(n7), .IN2(in3[35]), .S(in2[34]), .Q(sumout[35]) );
  INVX0 U16 ( .INP(in1[32]), .ZN(n8) );
  FADDX1 U17 ( .A(in1[10]), .B(in2[10]), .CI(in3[10]), .CO(cout[10]), .S(
        sumout[10]) );
  FADDX1 U18 ( .A(in1[11]), .B(in2[11]), .CI(in3[11]), .CO(cout[11]), .S(
        sumout[11]) );
  FADDX1 U19 ( .A(in1[12]), .B(in2[12]), .CI(in3[12]), .CO(cout[12]), .S(
        sumout[12]) );
  FADDX1 U20 ( .A(in1[13]), .B(in2[13]), .CI(in3[13]), .CO(cout[13]), .S(
        sumout[13]) );
  FADDX1 U21 ( .A(in1[14]), .B(in2[14]), .CI(in3[14]), .CO(cout[14]), .S(
        sumout[14]) );
  FADDX1 U22 ( .A(in1[15]), .B(in2[15]), .CI(in3[15]), .CO(cout[15]), .S(
        sumout[15]) );
  FADDX1 U23 ( .A(in1[16]), .B(in2[16]), .CI(in3[16]), .CO(cout[16]), .S(
        sumout[16]) );
  FADDX1 U24 ( .A(in1[17]), .B(in2[17]), .CI(in3[17]), .CO(cout[17]), .S(
        sumout[17]) );
  FADDX1 U25 ( .A(in1[18]), .B(in2[18]), .CI(in3[18]), .CO(cout[18]), .S(
        sumout[18]) );
  FADDX1 U26 ( .A(in1[19]), .B(in2[19]), .CI(in3[19]), .CO(cout[19]), .S(
        sumout[19]) );
  FADDX1 U27 ( .A(in1[20]), .B(in2[20]), .CI(in3[20]), .CO(cout[20]), .S(
        sumout[20]) );
  FADDX1 U28 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U29 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U30 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U31 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U32 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U33 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U34 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U35 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U36 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U37 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U38 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U39 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
  FADDX1 U40 ( .A(in2[33]), .B(in3[33]), .CI(n8), .CO(cout[33]), .S(sumout[33]) );
endmodule


module csa51squ_24 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n2, n3, n4, n5;

  NBUFFX2 U1 ( .INP(in3[31]), .Z(sumout[31]) );
  AND2X1 U2 ( .IN1(in2[2]), .IN2(in1[2]), .Q(cout[2]) );
  AND2X1 U3 ( .IN1(in2[3]), .IN2(in1[3]), .Q(cout[3]) );
  NOR2X0 U4 ( .IN1(in2[3]), .IN2(in1[3]), .QN(n2) );
  NOR2X0 U5 ( .IN1(n2), .IN2(cout[3]), .QN(sumout[3]) );
  AND2X1 U6 ( .IN1(in2[28]), .IN2(in3[28]), .Q(cout[28]) );
  NOR2X0 U7 ( .IN1(in2[28]), .IN2(in3[28]), .QN(n3) );
  NOR2X0 U8 ( .IN1(n3), .IN2(cout[28]), .QN(sumout[28]) );
  INVX0 U9 ( .INP(in3[29]), .ZN(n4) );
  NOR2X0 U10 ( .IN1(in2[28]), .IN2(n4), .QN(cout[29]) );
  MUX21X1 U11 ( .IN1(n4), .IN2(in3[29]), .S(in2[28]), .Q(sumout[29]) );
  INVX0 U12 ( .INP(in1[26]), .ZN(n5) );
  FADDX1 U13 ( .A(in1[10]), .B(in2[10]), .CI(in3[10]), .CO(cout[10]), .S(
        sumout[10]) );
  FADDX1 U14 ( .A(in1[11]), .B(in2[11]), .CI(in3[11]), .CO(cout[11]), .S(
        sumout[11]) );
  FADDX1 U15 ( .A(in1[12]), .B(in2[12]), .CI(in3[12]), .CO(cout[12]), .S(
        sumout[12]) );
  FADDX1 U16 ( .A(in1[13]), .B(in2[13]), .CI(in3[13]), .CO(cout[13]), .S(
        sumout[13]) );
  FADDX1 U17 ( .A(in1[14]), .B(in2[14]), .CI(in3[14]), .CO(cout[14]), .S(
        sumout[14]) );
  FADDX1 U18 ( .A(in1[15]), .B(in2[15]), .CI(in3[15]), .CO(cout[15]), .S(
        sumout[15]) );
  FADDX1 U19 ( .A(in1[16]), .B(in2[16]), .CI(in3[16]), .CO(cout[16]), .S(
        sumout[16]) );
  FADDX1 U20 ( .A(in1[17]), .B(in2[17]), .CI(in3[17]), .CO(cout[17]), .S(
        sumout[17]) );
  FADDX1 U21 ( .A(in1[18]), .B(in2[18]), .CI(in3[18]), .CO(cout[18]), .S(
        sumout[18]) );
  FADDX1 U22 ( .A(in1[19]), .B(in2[19]), .CI(in3[19]), .CO(cout[19]), .S(
        sumout[19]) );
  FADDX1 U23 ( .A(in1[20]), .B(in2[20]), .CI(in3[20]), .CO(cout[20]), .S(
        sumout[20]) );
  FADDX1 U24 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U25 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U26 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U27 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U28 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U29 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U30 ( .A(in2[27]), .B(in3[27]), .CI(n5), .CO(cout[27]), .S(sumout[27]) );
  FADDX1 U31 ( .A(in1[4]), .B(in2[4]), .CI(in3[4]), .CO(cout[4]), .S(sumout[4]) );
  FADDX1 U32 ( .A(in1[5]), .B(in2[5]), .CI(in3[5]), .CO(cout[5]), .S(sumout[5]) );
  FADDX1 U33 ( .A(in1[6]), .B(in2[6]), .CI(in3[6]), .CO(cout[6]), .S(sumout[6]) );
  FADDX1 U34 ( .A(in1[7]), .B(in2[7]), .CI(in3[7]), .CO(cout[7]), .S(sumout[7]) );
  FADDX1 U35 ( .A(in1[8]), .B(in2[8]), .CI(in3[8]), .CO(cout[8]), .S(sumout[8]) );
  FADDX1 U36 ( .A(in1[9]), .B(in2[9]), .CI(in3[9]), .CO(cout[9]), .S(sumout[9]) );
endmodule


module booth27_14 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;


  NBUFFX2 U3 ( .INP(in2[22]), .Z(out1[22]) );
  NBUFFX2 U4 ( .INP(in2[21]), .Z(out1[21]) );
  NBUFFX2 U5 ( .INP(in2[20]), .Z(out1[20]) );
  NBUFFX2 U6 ( .INP(in2[0]), .Z(out1[0]) );
  NBUFFX2 U7 ( .INP(in2[19]), .Z(out1[19]) );
  NBUFFX2 U8 ( .INP(in2[18]), .Z(out1[18]) );
  NBUFFX2 U9 ( .INP(in2[2]), .Z(out1[2]) );
  NBUFFX2 U10 ( .INP(in2[1]), .Z(out1[1]) );
  NBUFFX2 U11 ( .INP(in2[6]), .Z(out1[6]) );
  NBUFFX2 U12 ( .INP(in2[5]), .Z(out1[5]) );
  NBUFFX2 U13 ( .INP(in2[4]), .Z(out1[4]) );
  NBUFFX2 U14 ( .INP(in2[3]), .Z(out1[3]) );
  NBUFFX2 U15 ( .INP(in2[9]), .Z(out1[9]) );
  NBUFFX2 U16 ( .INP(in2[8]), .Z(out1[8]) );
  NBUFFX2 U17 ( .INP(in2[7]), .Z(out1[7]) );
  NBUFFX2 U18 ( .INP(in2[11]), .Z(out1[11]) );
  NBUFFX2 U19 ( .INP(in2[10]), .Z(out1[10]) );
  NBUFFX2 U20 ( .INP(in2[13]), .Z(out1[13]) );
  NBUFFX2 U21 ( .INP(in2[12]), .Z(out1[12]) );
  NBUFFX2 U22 ( .INP(in2[17]), .Z(out1[17]) );
  NBUFFX2 U23 ( .INP(in2[16]), .Z(out1[16]) );
  NBUFFX2 U24 ( .INP(in2[15]), .Z(out1[15]) );
  NBUFFX2 U25 ( .INP(in2[14]), .Z(out1[14]) );
endmodule


module booth27_15 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76;

  NAND2X0 U3 ( .IN1(n1), .IN2(n2), .QN(n8) );
  NAND2X0 U4 ( .IN1(n16), .IN2(in2[4]), .QN(n17) );
  NAND2X0 U5 ( .IN1(n19), .IN2(in2[5]), .QN(n20) );
  NAND2X0 U6 ( .IN1(n22), .IN2(in2[6]), .QN(n23) );
  NAND2X0 U7 ( .IN1(n25), .IN2(in2[7]), .QN(n26) );
  NAND2X0 U8 ( .IN1(n28), .IN2(in2[8]), .QN(n29) );
  NAND2X0 U9 ( .IN1(n31), .IN2(in2[9]), .QN(n32) );
  NAND2X0 U10 ( .IN1(n34), .IN2(in2[10]), .QN(n35) );
  NAND2X0 U11 ( .IN1(n37), .IN2(in2[11]), .QN(n38) );
  NAND2X0 U12 ( .IN1(n43), .IN2(in2[13]), .QN(n44) );
  NAND2X0 U13 ( .IN1(n46), .IN2(in2[14]), .QN(n47) );
  NAND2X0 U14 ( .IN1(n49), .IN2(in2[15]), .QN(n50) );
  NAND2X0 U15 ( .IN1(n52), .IN2(in2[16]), .QN(n53) );
  NAND2X0 U16 ( .IN1(n55), .IN2(in2[17]), .QN(n56) );
  NAND2X0 U17 ( .IN1(n7), .IN2(n15), .QN(out1[1]) );
  NAND2X0 U18 ( .IN1(n10), .IN2(n9), .QN(out1[2]) );
  NAND2X0 U19 ( .IN1(n58), .IN2(in2[18]), .QN(n59) );
  NAND2X0 U20 ( .IN1(n61), .IN2(in2[19]), .QN(n62) );
  NAND2X0 U21 ( .IN1(in1[1]), .IN2(in1[0]), .QN(out1[25]) );
  NOR2X0 U22 ( .IN1(in1[1]), .IN2(in1[0]), .QN(n71) );
  INVX0 U23 ( .INP(in2[0]), .ZN(n1) );
  INVX0 U24 ( .INP(in2[1]), .ZN(n2) );
  INVX0 U25 ( .INP(in2[3]), .ZN(n3) );
  INVX0 U26 ( .INP(in2[21]), .ZN(n4) );
  INVX0 U27 ( .INP(in2[22]), .ZN(n5) );
  INVX0 U28 ( .INP(in1[1]), .ZN(n6) );
  MUX21X1 U29 ( .IN1(in1[1]), .IN2(n6), .S(in1[0]), .Q(n74) );
  INVX0 U30 ( .INP(n74), .ZN(n76) );
  AO221X1 U31 ( .IN1(in2[0]), .IN2(in2[1]), .IN3(n1), .IN4(n2), .IN5(n76), .Q(
        n7) );
  NAND2X0 U32 ( .IN1(n71), .IN2(in2[0]), .QN(n15) );
  MUX21X1 U33 ( .IN1(n2), .IN2(n8), .S(in2[2]), .Q(n12) );
  AO221X1 U34 ( .IN1(n12), .IN2(in2[2]), .IN3(n12), .IN4(n1), .IN5(n76), .Q(
        n10) );
  INVX0 U35 ( .INP(n71), .ZN(n13) );
  AO221X1 U36 ( .IN1(in2[0]), .IN2(in2[1]), .IN3(n1), .IN4(n2), .IN5(n13), .Q(
        n9) );
  NOR3X0 U37 ( .IN1(in2[0]), .IN2(in2[2]), .IN3(in2[1]), .QN(n11) );
  OR4X1 U38 ( .IN1(in2[3]), .IN2(in2[0]), .IN3(in2[2]), .IN4(in2[1]), .Q(n16)
         );
  OA21X1 U39 ( .IN1(n11), .IN2(n3), .IN3(n16), .Q(n18) );
  INVX0 U40 ( .INP(n18), .ZN(n14) );
  OAI222X1 U41 ( .IN1(n15), .IN2(in2[2]), .IN3(n14), .IN4(n76), .IN5(n13), 
        .IN6(n12), .QN(out1[3]) );
  OR2X1 U42 ( .IN1(in2[4]), .IN2(n16), .Q(n19) );
  AND2X1 U43 ( .IN1(n19), .IN2(n17), .Q(n21) );
  AO22X1 U44 ( .IN1(n71), .IN2(n18), .IN3(n21), .IN4(n74), .Q(out1[4]) );
  OR2X1 U45 ( .IN1(in2[5]), .IN2(n19), .Q(n22) );
  AND2X1 U46 ( .IN1(n22), .IN2(n20), .Q(n24) );
  AO22X1 U47 ( .IN1(n71), .IN2(n21), .IN3(n24), .IN4(n74), .Q(out1[5]) );
  OR2X1 U48 ( .IN1(in2[6]), .IN2(n22), .Q(n25) );
  AND2X1 U49 ( .IN1(n25), .IN2(n23), .Q(n27) );
  AO22X1 U50 ( .IN1(n71), .IN2(n24), .IN3(n27), .IN4(n74), .Q(out1[6]) );
  OR2X1 U51 ( .IN1(in2[7]), .IN2(n25), .Q(n28) );
  AND2X1 U52 ( .IN1(n28), .IN2(n26), .Q(n30) );
  AO22X1 U53 ( .IN1(n71), .IN2(n27), .IN3(n30), .IN4(n74), .Q(out1[7]) );
  OR2X1 U54 ( .IN1(in2[8]), .IN2(n28), .Q(n31) );
  AND2X1 U55 ( .IN1(n31), .IN2(n29), .Q(n33) );
  AO22X1 U56 ( .IN1(n71), .IN2(n30), .IN3(n33), .IN4(n74), .Q(out1[8]) );
  OR2X1 U57 ( .IN1(in2[9]), .IN2(n31), .Q(n34) );
  AND2X1 U58 ( .IN1(n34), .IN2(n32), .Q(n36) );
  AO22X1 U59 ( .IN1(n71), .IN2(n33), .IN3(n36), .IN4(n74), .Q(out1[9]) );
  OR2X1 U60 ( .IN1(in2[10]), .IN2(n34), .Q(n37) );
  AND2X1 U61 ( .IN1(n37), .IN2(n35), .Q(n39) );
  AO22X1 U62 ( .IN1(n71), .IN2(n36), .IN3(n39), .IN4(n74), .Q(out1[10]) );
  OR2X1 U63 ( .IN1(in2[11]), .IN2(n37), .Q(n40) );
  AND2X1 U64 ( .IN1(n40), .IN2(n38), .Q(n42) );
  AO22X1 U65 ( .IN1(n71), .IN2(n39), .IN3(n42), .IN4(n74), .Q(out1[11]) );
  OR2X1 U66 ( .IN1(in2[12]), .IN2(n40), .Q(n43) );
  NAND2X0 U67 ( .IN1(n40), .IN2(in2[12]), .QN(n41) );
  AND2X1 U68 ( .IN1(n43), .IN2(n41), .Q(n45) );
  AO22X1 U69 ( .IN1(n71), .IN2(n42), .IN3(n45), .IN4(n74), .Q(out1[12]) );
  OR2X1 U70 ( .IN1(in2[13]), .IN2(n43), .Q(n46) );
  AND2X1 U71 ( .IN1(n46), .IN2(n44), .Q(n48) );
  AO22X1 U72 ( .IN1(n71), .IN2(n45), .IN3(n48), .IN4(n74), .Q(out1[13]) );
  OR2X1 U73 ( .IN1(in2[14]), .IN2(n46), .Q(n49) );
  AND2X1 U74 ( .IN1(n49), .IN2(n47), .Q(n51) );
  AO22X1 U75 ( .IN1(n71), .IN2(n48), .IN3(n51), .IN4(n74), .Q(out1[14]) );
  OR2X1 U76 ( .IN1(in2[15]), .IN2(n49), .Q(n52) );
  AND2X1 U77 ( .IN1(n52), .IN2(n50), .Q(n54) );
  AO22X1 U78 ( .IN1(n71), .IN2(n51), .IN3(n54), .IN4(n74), .Q(out1[15]) );
  OR2X1 U79 ( .IN1(in2[16]), .IN2(n52), .Q(n55) );
  AND2X1 U80 ( .IN1(n55), .IN2(n53), .Q(n57) );
  AO22X1 U81 ( .IN1(n71), .IN2(n54), .IN3(n57), .IN4(n74), .Q(out1[16]) );
  OR2X1 U82 ( .IN1(in2[17]), .IN2(n55), .Q(n58) );
  AND2X1 U83 ( .IN1(n58), .IN2(n56), .Q(n60) );
  AO22X1 U84 ( .IN1(n71), .IN2(n57), .IN3(n60), .IN4(n74), .Q(out1[17]) );
  OR2X1 U85 ( .IN1(in2[18]), .IN2(n58), .Q(n61) );
  AND2X1 U86 ( .IN1(n61), .IN2(n59), .Q(n63) );
  AO22X1 U87 ( .IN1(n71), .IN2(n60), .IN3(n63), .IN4(n74), .Q(out1[18]) );
  OR2X1 U88 ( .IN1(in2[19]), .IN2(n61), .Q(n64) );
  AND2X1 U89 ( .IN1(n64), .IN2(n62), .Q(n65) );
  AO22X1 U90 ( .IN1(n71), .IN2(n63), .IN3(n65), .IN4(n74), .Q(out1[19]) );
  NOR2X0 U91 ( .IN1(in2[20]), .IN2(n64), .QN(n72) );
  AOI21X1 U92 ( .IN1(in2[20]), .IN2(n64), .IN3(n72), .QN(n66) );
  AO22X1 U93 ( .IN1(n71), .IN2(n65), .IN3(n66), .IN4(n74), .Q(out1[20]) );
  MUX21X1 U94 ( .IN1(n4), .IN2(in2[21]), .S(n72), .Q(n69) );
  AO22X1 U95 ( .IN1(n71), .IN2(n66), .IN3(n69), .IN4(n74), .Q(out1[21]) );
  INVX0 U96 ( .INP(n72), .ZN(n67) );
  NOR2X0 U97 ( .IN1(in2[21]), .IN2(n67), .QN(n70) );
  MUX21X1 U98 ( .IN1(n5), .IN2(in2[22]), .S(n70), .Q(n68) );
  AO22X1 U99 ( .IN1(n71), .IN2(n69), .IN3(n68), .IN4(n74), .Q(out1[22]) );
  MUX21X1 U100 ( .IN1(n71), .IN2(n74), .S(n70), .Q(n73) );
  AND3X1 U101 ( .IN1(n72), .IN2(n71), .IN3(n4), .Q(n75) );
  MUX21X1 U102 ( .IN1(n73), .IN2(n75), .S(in2[22]), .Q(out1[23]) );
  AO21X1 U103 ( .IN1(n75), .IN2(n5), .IN3(n74), .Q(out1[24]) );
  NOR2X0 U104 ( .IN1(n76), .IN2(n1), .QN(out1[0]) );
endmodule


module booth27_16 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n25), .IN2(n6), .QN(n30) );
  NAND2X0 U4 ( .IN1(n33), .IN2(n7), .QN(n37) );
  NAND2X0 U5 ( .IN1(n41), .IN2(n8), .QN(n45) );
  NAND2X0 U6 ( .IN1(n49), .IN2(n9), .QN(n53) );
  NAND2X0 U7 ( .IN1(n57), .IN2(n10), .QN(n61) );
  NAND2X0 U8 ( .IN1(n65), .IN2(n11), .QN(n77) );
  NAND2X0 U9 ( .IN1(n81), .IN2(n13), .QN(n89) );
  NAND2X0 U10 ( .IN1(n93), .IN2(n15), .QN(n101) );
  NAND2X0 U11 ( .IN1(n105), .IN2(n17), .QN(n114) );
  NAND2X0 U12 ( .IN1(n27), .IN2(n132), .QN(n4) );
  NAND2X0 U13 ( .IN1(in1[2]), .IN2(n77), .QN(n71) );
  NAND2X0 U14 ( .IN1(n70), .IN2(n132), .QN(n74) );
  NAND2X0 U15 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U16 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U17 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U18 ( .IN1(n118), .IN2(n19), .QN(n125) );
  NAND2X0 U19 ( .IN1(n141), .IN2(n130), .QN(n24) );
  NAND2X0 U20 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NAND2X0 U21 ( .IN1(n32), .IN2(n31), .QN(out1[3]) );
  NAND2X0 U22 ( .IN1(n36), .IN2(n35), .QN(out1[4]) );
  NAND2X0 U23 ( .IN1(n40), .IN2(n39), .QN(out1[5]) );
  NAND2X0 U24 ( .IN1(n44), .IN2(n43), .QN(out1[6]) );
  NAND2X0 U25 ( .IN1(n48), .IN2(n47), .QN(out1[7]) );
  NAND2X0 U26 ( .IN1(n52), .IN2(n51), .QN(out1[8]) );
  NAND2X0 U27 ( .IN1(n56), .IN2(n55), .QN(out1[9]) );
  NAND2X0 U28 ( .IN1(n60), .IN2(n59), .QN(out1[10]) );
  NAND2X0 U29 ( .IN1(n64), .IN2(n63), .QN(out1[11]) );
  NAND2X0 U30 ( .IN1(n69), .IN2(n68), .QN(out1[12]) );
  NAND2X0 U31 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U32 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U33 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U34 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U35 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U36 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U37 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U38 ( .IN1(n23), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U39 ( .IN1(in1[2]), .IN2(n22), .QN(n23) );
  NOR2X0 U40 ( .IN1(n28), .IN2(n26), .QN(n3) );
  NOR2X0 U41 ( .IN1(n142), .IN2(n21), .QN(n1) );
  NOR2X0 U42 ( .IN1(n142), .IN2(n111), .QN(n138) );
  INVX0 U43 ( .INP(n130), .ZN(n137) );
  INVX0 U44 ( .INP(n132), .ZN(n141) );
  NOR3X0 U45 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  NAND3X0 U46 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  MUX21X1 U47 ( .IN1(n22), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  INVX0 U48 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U49 ( .INP(in2[2]), .ZN(n6) );
  INVX0 U50 ( .INP(in2[4]), .ZN(n7) );
  INVX0 U51 ( .INP(in2[6]), .ZN(n8) );
  INVX0 U52 ( .INP(in2[8]), .ZN(n9) );
  INVX0 U53 ( .INP(in2[10]), .ZN(n10) );
  INVX0 U54 ( .INP(in2[12]), .ZN(n11) );
  INVX0 U55 ( .INP(in2[13]), .ZN(n12) );
  INVX0 U56 ( .INP(in2[14]), .ZN(n13) );
  INVX0 U57 ( .INP(in2[15]), .ZN(n14) );
  INVX0 U58 ( .INP(in2[16]), .ZN(n15) );
  INVX0 U59 ( .INP(in2[17]), .ZN(n16) );
  INVX0 U60 ( .INP(in2[18]), .ZN(n17) );
  INVX0 U61 ( .INP(in2[19]), .ZN(n18) );
  INVX0 U62 ( .INP(in2[20]), .ZN(n19) );
  INVX0 U63 ( .INP(in2[21]), .ZN(n20) );
  INVX0 U64 ( .INP(in2[22]), .ZN(n21) );
  INVX0 U65 ( .INP(in1[1]), .ZN(n22) );
  INVX0 U66 ( .INP(in1[2]), .ZN(n111) );
  INVX0 U67 ( .INP(n138), .ZN(n140) );
  NOR2X0 U68 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n25) );
  AOI21X1 U69 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n25), .QN(n27) );
  NOR2X0 U70 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U71 ( .IN1(n24), .IN2(in2[0]), .IN3(n138), .IN4(n27), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U72 ( .INP(n133), .ZN(n67) );
  NOR2X0 U73 ( .IN1(n67), .IN2(n6), .QN(n28) );
  OA21X1 U74 ( .IN1(n25), .IN2(n6), .IN3(n30), .Q(n29) );
  AO22X1 U75 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n29), .Q(n26) );
  AOI22X1 U76 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n29), .QN(n32) );
  NOR2X0 U77 ( .IN1(in2[3]), .IN2(n30), .QN(n33) );
  AO21X1 U78 ( .IN1(in2[3]), .IN2(n30), .IN3(n33), .Q(n34) );
  OA22X1 U79 ( .IN1(n6), .IN2(n130), .IN3(n140), .IN4(n34), .Q(n31) );
  OA21X1 U80 ( .IN1(n33), .IN2(n7), .IN3(n37), .Q(n38) );
  AOI22X1 U81 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n38), .QN(n36) );
  OA22X1 U82 ( .IN1(n67), .IN2(n7), .IN3(n141), .IN4(n34), .Q(n35) );
  NOR2X0 U83 ( .IN1(in2[5]), .IN2(n37), .QN(n41) );
  AO21X1 U84 ( .IN1(in2[5]), .IN2(n37), .IN3(n41), .Q(n42) );
  OA22X1 U85 ( .IN1(n7), .IN2(n130), .IN3(n140), .IN4(n42), .Q(n40) );
  AOI22X1 U86 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n38), .QN(n39) );
  OA21X1 U87 ( .IN1(n41), .IN2(n8), .IN3(n45), .Q(n46) );
  AOI22X1 U88 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n46), .QN(n44) );
  OA22X1 U89 ( .IN1(n67), .IN2(n8), .IN3(n141), .IN4(n42), .Q(n43) );
  NOR2X0 U90 ( .IN1(in2[7]), .IN2(n45), .QN(n49) );
  AO21X1 U91 ( .IN1(in2[7]), .IN2(n45), .IN3(n49), .Q(n50) );
  OA22X1 U92 ( .IN1(n8), .IN2(n130), .IN3(n140), .IN4(n50), .Q(n48) );
  AOI22X1 U93 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n46), .QN(n47) );
  OA21X1 U94 ( .IN1(n49), .IN2(n9), .IN3(n53), .Q(n54) );
  AOI22X1 U95 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n54), .QN(n52) );
  OA22X1 U96 ( .IN1(n67), .IN2(n9), .IN3(n141), .IN4(n50), .Q(n51) );
  NOR2X0 U97 ( .IN1(in2[9]), .IN2(n53), .QN(n57) );
  AO21X1 U98 ( .IN1(in2[9]), .IN2(n53), .IN3(n57), .Q(n58) );
  OA22X1 U99 ( .IN1(n9), .IN2(n130), .IN3(n140), .IN4(n58), .Q(n56) );
  AOI22X1 U100 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n54), .QN(n55) );
  OA21X1 U101 ( .IN1(n57), .IN2(n10), .IN3(n61), .Q(n62) );
  AOI22X1 U102 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n62), .QN(n60) );
  OA22X1 U103 ( .IN1(n67), .IN2(n10), .IN3(n141), .IN4(n58), .Q(n59) );
  NOR2X0 U104 ( .IN1(in2[11]), .IN2(n61), .QN(n65) );
  AO21X1 U105 ( .IN1(in2[11]), .IN2(n61), .IN3(n65), .Q(n66) );
  OA22X1 U106 ( .IN1(n10), .IN2(n130), .IN3(n140), .IN4(n66), .Q(n64) );
  AOI22X1 U107 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n62), .QN(n63) );
  OA21X1 U108 ( .IN1(n65), .IN2(n11), .IN3(n77), .Q(n70) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n70), .QN(n69) );
  OA22X1 U110 ( .IN1(n67), .IN2(n11), .IN3(n141), .IN4(n66), .Q(n68) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n12), .S(n71), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n11), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n13), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n12), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n12), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n14), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n13), .IN4(n85), .IN5(n84), 
        .Q(out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n15), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n14), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n14), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n16), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n15), .IN4(n97), .IN5(n96), 
        .Q(out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n17), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n16), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n16), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n18), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n17), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n19), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n18), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n18), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n20), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n19), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n21), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n20), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n20), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n21), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_17 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n33), .IN2(n7), .QN(n37) );
  NAND2X0 U4 ( .IN1(n41), .IN2(n8), .QN(n45) );
  NAND2X0 U5 ( .IN1(n49), .IN2(n9), .QN(n53) );
  NAND2X0 U6 ( .IN1(n57), .IN2(n10), .QN(n61) );
  NAND2X0 U7 ( .IN1(n25), .IN2(n6), .QN(n30) );
  NAND2X0 U8 ( .IN1(n65), .IN2(n11), .QN(n77) );
  NAND2X0 U9 ( .IN1(n81), .IN2(n13), .QN(n89) );
  NAND2X0 U10 ( .IN1(n93), .IN2(n15), .QN(n101) );
  NAND2X0 U11 ( .IN1(n105), .IN2(n17), .QN(n114) );
  NAND2X0 U12 ( .IN1(n118), .IN2(n19), .QN(n125) );
  NAND2X0 U13 ( .IN1(in1[2]), .IN2(n77), .QN(n71) );
  NAND2X0 U14 ( .IN1(n70), .IN2(n132), .QN(n74) );
  NAND2X0 U15 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U16 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U17 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U18 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U19 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U20 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U21 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U22 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NAND2X0 U23 ( .IN1(n27), .IN2(n132), .QN(n4) );
  NAND2X0 U24 ( .IN1(n32), .IN2(n31), .QN(out1[3]) );
  NAND2X0 U25 ( .IN1(n36), .IN2(n35), .QN(out1[4]) );
  NAND2X0 U26 ( .IN1(n40), .IN2(n39), .QN(out1[5]) );
  NAND2X0 U27 ( .IN1(n44), .IN2(n43), .QN(out1[6]) );
  NAND2X0 U28 ( .IN1(n48), .IN2(n47), .QN(out1[7]) );
  NAND2X0 U29 ( .IN1(n52), .IN2(n51), .QN(out1[8]) );
  NAND2X0 U30 ( .IN1(n56), .IN2(n55), .QN(out1[9]) );
  NAND2X0 U31 ( .IN1(n60), .IN2(n59), .QN(out1[10]) );
  NAND2X0 U32 ( .IN1(n64), .IN2(n63), .QN(out1[11]) );
  NAND2X0 U33 ( .IN1(n69), .IN2(n68), .QN(out1[12]) );
  NAND2X0 U34 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U35 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U36 ( .IN1(n141), .IN2(n130), .QN(n24) );
  NAND2X0 U37 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U38 ( .IN1(n23), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U39 ( .IN1(in1[2]), .IN2(n22), .QN(n23) );
  NOR2X0 U40 ( .IN1(n28), .IN2(n26), .QN(n3) );
  NOR2X0 U41 ( .IN1(n142), .IN2(n111), .QN(n138) );
  NOR2X0 U42 ( .IN1(n142), .IN2(n21), .QN(n1) );
  INVX0 U43 ( .INP(n130), .ZN(n137) );
  INVX0 U44 ( .INP(n132), .ZN(n141) );
  NOR3X0 U45 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  NAND3X0 U46 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  MUX21X1 U47 ( .IN1(n22), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  INVX0 U48 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U49 ( .INP(in2[2]), .ZN(n6) );
  INVX0 U50 ( .INP(in2[4]), .ZN(n7) );
  INVX0 U51 ( .INP(in2[6]), .ZN(n8) );
  INVX0 U52 ( .INP(in2[8]), .ZN(n9) );
  INVX0 U53 ( .INP(in2[10]), .ZN(n10) );
  INVX0 U54 ( .INP(in2[12]), .ZN(n11) );
  INVX0 U55 ( .INP(in2[13]), .ZN(n12) );
  INVX0 U56 ( .INP(in2[14]), .ZN(n13) );
  INVX0 U57 ( .INP(in2[15]), .ZN(n14) );
  INVX0 U58 ( .INP(in2[16]), .ZN(n15) );
  INVX0 U59 ( .INP(in2[17]), .ZN(n16) );
  INVX0 U60 ( .INP(in2[18]), .ZN(n17) );
  INVX0 U61 ( .INP(in2[19]), .ZN(n18) );
  INVX0 U62 ( .INP(in2[20]), .ZN(n19) );
  INVX0 U63 ( .INP(in2[21]), .ZN(n20) );
  INVX0 U64 ( .INP(in2[22]), .ZN(n21) );
  INVX0 U65 ( .INP(in1[1]), .ZN(n22) );
  INVX0 U66 ( .INP(in1[2]), .ZN(n111) );
  INVX0 U67 ( .INP(n138), .ZN(n140) );
  NOR2X0 U68 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n25) );
  AOI21X1 U69 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n25), .QN(n27) );
  NOR2X0 U70 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U71 ( .IN1(n24), .IN2(in2[0]), .IN3(n138), .IN4(n27), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U72 ( .INP(n133), .ZN(n67) );
  NOR2X0 U73 ( .IN1(n67), .IN2(n6), .QN(n28) );
  OA21X1 U74 ( .IN1(n25), .IN2(n6), .IN3(n30), .Q(n29) );
  AO22X1 U75 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n29), .Q(n26) );
  AOI22X1 U76 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n29), .QN(n32) );
  NOR2X0 U77 ( .IN1(in2[3]), .IN2(n30), .QN(n33) );
  AO21X1 U78 ( .IN1(in2[3]), .IN2(n30), .IN3(n33), .Q(n34) );
  OA22X1 U79 ( .IN1(n6), .IN2(n130), .IN3(n140), .IN4(n34), .Q(n31) );
  OA21X1 U80 ( .IN1(n33), .IN2(n7), .IN3(n37), .Q(n38) );
  AOI22X1 U81 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n38), .QN(n36) );
  OA22X1 U82 ( .IN1(n67), .IN2(n7), .IN3(n141), .IN4(n34), .Q(n35) );
  NOR2X0 U83 ( .IN1(in2[5]), .IN2(n37), .QN(n41) );
  AO21X1 U84 ( .IN1(in2[5]), .IN2(n37), .IN3(n41), .Q(n42) );
  OA22X1 U85 ( .IN1(n7), .IN2(n130), .IN3(n140), .IN4(n42), .Q(n40) );
  AOI22X1 U86 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n38), .QN(n39) );
  OA21X1 U87 ( .IN1(n41), .IN2(n8), .IN3(n45), .Q(n46) );
  AOI22X1 U88 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n46), .QN(n44) );
  OA22X1 U89 ( .IN1(n67), .IN2(n8), .IN3(n141), .IN4(n42), .Q(n43) );
  NOR2X0 U90 ( .IN1(in2[7]), .IN2(n45), .QN(n49) );
  AO21X1 U91 ( .IN1(in2[7]), .IN2(n45), .IN3(n49), .Q(n50) );
  OA22X1 U92 ( .IN1(n8), .IN2(n130), .IN3(n140), .IN4(n50), .Q(n48) );
  AOI22X1 U93 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n46), .QN(n47) );
  OA21X1 U94 ( .IN1(n49), .IN2(n9), .IN3(n53), .Q(n54) );
  AOI22X1 U95 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n54), .QN(n52) );
  OA22X1 U96 ( .IN1(n67), .IN2(n9), .IN3(n141), .IN4(n50), .Q(n51) );
  NOR2X0 U97 ( .IN1(in2[9]), .IN2(n53), .QN(n57) );
  AO21X1 U98 ( .IN1(in2[9]), .IN2(n53), .IN3(n57), .Q(n58) );
  OA22X1 U99 ( .IN1(n9), .IN2(n130), .IN3(n140), .IN4(n58), .Q(n56) );
  AOI22X1 U100 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n54), .QN(n55) );
  OA21X1 U101 ( .IN1(n57), .IN2(n10), .IN3(n61), .Q(n62) );
  AOI22X1 U102 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n62), .QN(n60) );
  OA22X1 U103 ( .IN1(n67), .IN2(n10), .IN3(n141), .IN4(n58), .Q(n59) );
  NOR2X0 U104 ( .IN1(in2[11]), .IN2(n61), .QN(n65) );
  AO21X1 U105 ( .IN1(in2[11]), .IN2(n61), .IN3(n65), .Q(n66) );
  OA22X1 U106 ( .IN1(n10), .IN2(n130), .IN3(n140), .IN4(n66), .Q(n64) );
  AOI22X1 U107 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n62), .QN(n63) );
  OA21X1 U108 ( .IN1(n65), .IN2(n11), .IN3(n77), .Q(n70) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n70), .QN(n69) );
  OA22X1 U110 ( .IN1(n67), .IN2(n11), .IN3(n141), .IN4(n66), .Q(n68) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n12), .S(n71), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n11), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n13), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n12), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n12), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n14), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n13), .IN4(n85), .IN5(n84), 
        .Q(out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n15), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n14), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n14), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n16), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n15), .IN4(n97), .IN5(n96), 
        .Q(out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n17), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n16), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n16), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n18), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n17), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n19), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n18), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n18), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n20), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n19), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n21), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n20), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n20), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n21), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_18 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n41), .IN2(n8), .QN(n45) );
  NAND2X0 U4 ( .IN1(n49), .IN2(n9), .QN(n53) );
  NAND2X0 U5 ( .IN1(n57), .IN2(n10), .QN(n61) );
  NAND2X0 U6 ( .IN1(n33), .IN2(n7), .QN(n37) );
  NAND2X0 U7 ( .IN1(n25), .IN2(n6), .QN(n30) );
  NAND2X0 U8 ( .IN1(n65), .IN2(n11), .QN(n77) );
  NAND2X0 U9 ( .IN1(n81), .IN2(n13), .QN(n89) );
  NAND2X0 U10 ( .IN1(n93), .IN2(n15), .QN(n101) );
  NAND2X0 U11 ( .IN1(in1[2]), .IN2(n77), .QN(n71) );
  NAND2X0 U12 ( .IN1(n70), .IN2(n132), .QN(n74) );
  NAND2X0 U13 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U14 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U15 ( .IN1(n105), .IN2(n17), .QN(n114) );
  NAND2X0 U16 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U17 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U18 ( .IN1(n27), .IN2(n132), .QN(n4) );
  NAND2X0 U19 ( .IN1(n141), .IN2(n130), .QN(n24) );
  NAND2X0 U20 ( .IN1(n40), .IN2(n39), .QN(out1[5]) );
  NAND2X0 U21 ( .IN1(n44), .IN2(n43), .QN(out1[6]) );
  NAND2X0 U22 ( .IN1(n48), .IN2(n47), .QN(out1[7]) );
  NAND2X0 U23 ( .IN1(n52), .IN2(n51), .QN(out1[8]) );
  NAND2X0 U24 ( .IN1(n56), .IN2(n55), .QN(out1[9]) );
  NAND2X0 U25 ( .IN1(n60), .IN2(n59), .QN(out1[10]) );
  NAND2X0 U26 ( .IN1(n64), .IN2(n63), .QN(out1[11]) );
  NAND2X0 U27 ( .IN1(n69), .IN2(n68), .QN(out1[12]) );
  NAND2X0 U28 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U29 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U30 ( .IN1(n118), .IN2(n19), .QN(n125) );
  NAND2X0 U31 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U32 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U33 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U34 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U35 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NAND2X0 U36 ( .IN1(n32), .IN2(n31), .QN(out1[3]) );
  NAND2X0 U37 ( .IN1(n36), .IN2(n35), .QN(out1[4]) );
  NAND2X0 U38 ( .IN1(n23), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U39 ( .IN1(in1[2]), .IN2(n22), .QN(n23) );
  INVX0 U40 ( .INP(in1[2]), .ZN(n111) );
  NOR2X0 U41 ( .IN1(n28), .IN2(n26), .QN(n3) );
  NOR2X0 U42 ( .IN1(n142), .IN2(n21), .QN(n1) );
  INVX0 U43 ( .INP(n132), .ZN(n141) );
  INVX0 U44 ( .INP(n130), .ZN(n137) );
  NOR2X0 U45 ( .IN1(n142), .IN2(n111), .QN(n138) );
  MUX21X1 U46 ( .IN1(n22), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  NAND3X0 U47 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  NOR3X0 U48 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  INVX0 U49 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U50 ( .INP(in2[2]), .ZN(n6) );
  INVX0 U51 ( .INP(in2[4]), .ZN(n7) );
  INVX0 U52 ( .INP(in2[6]), .ZN(n8) );
  INVX0 U53 ( .INP(in2[8]), .ZN(n9) );
  INVX0 U54 ( .INP(in2[10]), .ZN(n10) );
  INVX0 U55 ( .INP(in2[12]), .ZN(n11) );
  INVX0 U56 ( .INP(in2[13]), .ZN(n12) );
  INVX0 U57 ( .INP(in2[14]), .ZN(n13) );
  INVX0 U58 ( .INP(in2[15]), .ZN(n14) );
  INVX0 U59 ( .INP(in2[16]), .ZN(n15) );
  INVX0 U60 ( .INP(in2[17]), .ZN(n16) );
  INVX0 U61 ( .INP(in2[18]), .ZN(n17) );
  INVX0 U62 ( .INP(in2[19]), .ZN(n18) );
  INVX0 U63 ( .INP(in2[20]), .ZN(n19) );
  INVX0 U64 ( .INP(in2[21]), .ZN(n20) );
  INVX0 U65 ( .INP(in2[22]), .ZN(n21) );
  INVX0 U66 ( .INP(in1[1]), .ZN(n22) );
  INVX0 U67 ( .INP(n138), .ZN(n140) );
  NOR2X0 U68 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n25) );
  AOI21X1 U69 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n25), .QN(n27) );
  NOR2X0 U70 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U71 ( .IN1(n24), .IN2(in2[0]), .IN3(n138), .IN4(n27), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U72 ( .INP(n133), .ZN(n67) );
  NOR2X0 U73 ( .IN1(n67), .IN2(n6), .QN(n28) );
  OA21X1 U74 ( .IN1(n25), .IN2(n6), .IN3(n30), .Q(n29) );
  AO22X1 U75 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n29), .Q(n26) );
  AOI22X1 U76 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n29), .QN(n32) );
  NOR2X0 U77 ( .IN1(in2[3]), .IN2(n30), .QN(n33) );
  AO21X1 U78 ( .IN1(in2[3]), .IN2(n30), .IN3(n33), .Q(n34) );
  OA22X1 U79 ( .IN1(n6), .IN2(n130), .IN3(n140), .IN4(n34), .Q(n31) );
  OA21X1 U80 ( .IN1(n33), .IN2(n7), .IN3(n37), .Q(n38) );
  AOI22X1 U81 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n38), .QN(n36) );
  OA22X1 U82 ( .IN1(n67), .IN2(n7), .IN3(n141), .IN4(n34), .Q(n35) );
  NOR2X0 U83 ( .IN1(in2[5]), .IN2(n37), .QN(n41) );
  AO21X1 U84 ( .IN1(in2[5]), .IN2(n37), .IN3(n41), .Q(n42) );
  OA22X1 U85 ( .IN1(n7), .IN2(n130), .IN3(n140), .IN4(n42), .Q(n40) );
  AOI22X1 U86 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n38), .QN(n39) );
  OA21X1 U87 ( .IN1(n41), .IN2(n8), .IN3(n45), .Q(n46) );
  AOI22X1 U88 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n46), .QN(n44) );
  OA22X1 U89 ( .IN1(n67), .IN2(n8), .IN3(n141), .IN4(n42), .Q(n43) );
  NOR2X0 U90 ( .IN1(in2[7]), .IN2(n45), .QN(n49) );
  AO21X1 U91 ( .IN1(in2[7]), .IN2(n45), .IN3(n49), .Q(n50) );
  OA22X1 U92 ( .IN1(n8), .IN2(n130), .IN3(n140), .IN4(n50), .Q(n48) );
  AOI22X1 U93 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n46), .QN(n47) );
  OA21X1 U94 ( .IN1(n49), .IN2(n9), .IN3(n53), .Q(n54) );
  AOI22X1 U95 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n54), .QN(n52) );
  OA22X1 U96 ( .IN1(n67), .IN2(n9), .IN3(n141), .IN4(n50), .Q(n51) );
  NOR2X0 U97 ( .IN1(in2[9]), .IN2(n53), .QN(n57) );
  AO21X1 U98 ( .IN1(in2[9]), .IN2(n53), .IN3(n57), .Q(n58) );
  OA22X1 U99 ( .IN1(n9), .IN2(n130), .IN3(n140), .IN4(n58), .Q(n56) );
  AOI22X1 U100 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n54), .QN(n55) );
  OA21X1 U101 ( .IN1(n57), .IN2(n10), .IN3(n61), .Q(n62) );
  AOI22X1 U102 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n62), .QN(n60) );
  OA22X1 U103 ( .IN1(n67), .IN2(n10), .IN3(n141), .IN4(n58), .Q(n59) );
  NOR2X0 U104 ( .IN1(in2[11]), .IN2(n61), .QN(n65) );
  AO21X1 U105 ( .IN1(in2[11]), .IN2(n61), .IN3(n65), .Q(n66) );
  OA22X1 U106 ( .IN1(n10), .IN2(n130), .IN3(n140), .IN4(n66), .Q(n64) );
  AOI22X1 U107 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n62), .QN(n63) );
  OA21X1 U108 ( .IN1(n65), .IN2(n11), .IN3(n77), .Q(n70) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n70), .QN(n69) );
  OA22X1 U110 ( .IN1(n67), .IN2(n11), .IN3(n141), .IN4(n66), .Q(n68) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n12), .S(n71), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n11), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n13), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n12), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n12), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n14), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n13), .IN4(n85), .IN5(n84), 
        .Q(out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n15), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n14), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n14), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n16), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n15), .IN4(n97), .IN5(n96), 
        .Q(out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n17), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n16), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n16), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n18), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n17), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n19), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n18), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n18), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n20), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n19), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n21), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n20), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n20), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n21), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_19 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n49), .IN2(n9), .QN(n53) );
  NAND2X0 U4 ( .IN1(n57), .IN2(n10), .QN(n61) );
  NAND2X0 U5 ( .IN1(n25), .IN2(n6), .QN(n30) );
  NAND2X0 U6 ( .IN1(n41), .IN2(n8), .QN(n45) );
  NAND2X0 U7 ( .IN1(n33), .IN2(n7), .QN(n37) );
  NAND2X0 U8 ( .IN1(n65), .IN2(n11), .QN(n77) );
  NAND2X0 U9 ( .IN1(n81), .IN2(n13), .QN(n89) );
  NAND2X0 U10 ( .IN1(n93), .IN2(n15), .QN(n101) );
  NAND2X0 U11 ( .IN1(n105), .IN2(n17), .QN(n114) );
  NAND2X0 U12 ( .IN1(in1[2]), .IN2(n77), .QN(n71) );
  NAND2X0 U13 ( .IN1(n70), .IN2(n132), .QN(n74) );
  NAND2X0 U14 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U15 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U16 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U17 ( .IN1(n118), .IN2(n19), .QN(n125) );
  NAND2X0 U18 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U19 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U20 ( .IN1(n27), .IN2(n132), .QN(n4) );
  NAND2X0 U21 ( .IN1(n48), .IN2(n47), .QN(out1[7]) );
  NAND2X0 U22 ( .IN1(n52), .IN2(n51), .QN(out1[8]) );
  NAND2X0 U23 ( .IN1(n56), .IN2(n55), .QN(out1[9]) );
  NAND2X0 U24 ( .IN1(n60), .IN2(n59), .QN(out1[10]) );
  NAND2X0 U25 ( .IN1(n64), .IN2(n63), .QN(out1[11]) );
  NAND2X0 U26 ( .IN1(n69), .IN2(n68), .QN(out1[12]) );
  NAND2X0 U27 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U28 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U29 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U30 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U31 ( .IN1(n141), .IN2(n130), .QN(n24) );
  NAND2X0 U32 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NAND2X0 U33 ( .IN1(n36), .IN2(n35), .QN(out1[4]) );
  NAND2X0 U34 ( .IN1(n32), .IN2(n31), .QN(out1[3]) );
  NAND2X0 U35 ( .IN1(n40), .IN2(n39), .QN(out1[5]) );
  NAND2X0 U36 ( .IN1(n44), .IN2(n43), .QN(out1[6]) );
  NAND2X0 U37 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U38 ( .IN1(n23), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U39 ( .IN1(in1[2]), .IN2(n22), .QN(n23) );
  NOR2X0 U40 ( .IN1(n28), .IN2(n26), .QN(n3) );
  INVX0 U41 ( .INP(n130), .ZN(n137) );
  NAND3X0 U42 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  NOR2X0 U43 ( .IN1(n142), .IN2(n21), .QN(n1) );
  NOR2X0 U44 ( .IN1(n142), .IN2(n111), .QN(n138) );
  MUX21X1 U45 ( .IN1(n22), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  INVX0 U46 ( .INP(n132), .ZN(n141) );
  NOR3X0 U47 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  INVX0 U48 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U49 ( .INP(in2[2]), .ZN(n6) );
  INVX0 U50 ( .INP(in2[4]), .ZN(n7) );
  INVX0 U51 ( .INP(in2[6]), .ZN(n8) );
  INVX0 U52 ( .INP(in2[8]), .ZN(n9) );
  INVX0 U53 ( .INP(in2[10]), .ZN(n10) );
  INVX0 U54 ( .INP(in2[12]), .ZN(n11) );
  INVX0 U55 ( .INP(in2[13]), .ZN(n12) );
  INVX0 U56 ( .INP(in2[14]), .ZN(n13) );
  INVX0 U57 ( .INP(in2[15]), .ZN(n14) );
  INVX0 U58 ( .INP(in2[16]), .ZN(n15) );
  INVX0 U59 ( .INP(in2[17]), .ZN(n16) );
  INVX0 U60 ( .INP(in2[18]), .ZN(n17) );
  INVX0 U61 ( .INP(in2[19]), .ZN(n18) );
  INVX0 U62 ( .INP(in2[20]), .ZN(n19) );
  INVX0 U63 ( .INP(in2[21]), .ZN(n20) );
  INVX0 U64 ( .INP(in2[22]), .ZN(n21) );
  INVX0 U65 ( .INP(in1[1]), .ZN(n22) );
  INVX0 U66 ( .INP(in1[2]), .ZN(n111) );
  INVX0 U67 ( .INP(n138), .ZN(n140) );
  NOR2X0 U68 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n25) );
  AOI21X1 U69 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n25), .QN(n27) );
  NOR2X0 U70 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U71 ( .IN1(n24), .IN2(in2[0]), .IN3(n138), .IN4(n27), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U72 ( .INP(n133), .ZN(n67) );
  NOR2X0 U73 ( .IN1(n67), .IN2(n6), .QN(n28) );
  OA21X1 U74 ( .IN1(n25), .IN2(n6), .IN3(n30), .Q(n29) );
  AO22X1 U75 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n29), .Q(n26) );
  AOI22X1 U76 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n29), .QN(n32) );
  NOR2X0 U77 ( .IN1(in2[3]), .IN2(n30), .QN(n33) );
  AO21X1 U78 ( .IN1(in2[3]), .IN2(n30), .IN3(n33), .Q(n34) );
  OA22X1 U79 ( .IN1(n6), .IN2(n130), .IN3(n140), .IN4(n34), .Q(n31) );
  OA21X1 U80 ( .IN1(n33), .IN2(n7), .IN3(n37), .Q(n38) );
  AOI22X1 U81 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n38), .QN(n36) );
  OA22X1 U82 ( .IN1(n67), .IN2(n7), .IN3(n141), .IN4(n34), .Q(n35) );
  NOR2X0 U83 ( .IN1(in2[5]), .IN2(n37), .QN(n41) );
  AO21X1 U84 ( .IN1(in2[5]), .IN2(n37), .IN3(n41), .Q(n42) );
  OA22X1 U85 ( .IN1(n7), .IN2(n130), .IN3(n140), .IN4(n42), .Q(n40) );
  AOI22X1 U86 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n38), .QN(n39) );
  OA21X1 U87 ( .IN1(n41), .IN2(n8), .IN3(n45), .Q(n46) );
  AOI22X1 U88 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n46), .QN(n44) );
  OA22X1 U89 ( .IN1(n67), .IN2(n8), .IN3(n141), .IN4(n42), .Q(n43) );
  NOR2X0 U90 ( .IN1(in2[7]), .IN2(n45), .QN(n49) );
  AO21X1 U91 ( .IN1(in2[7]), .IN2(n45), .IN3(n49), .Q(n50) );
  OA22X1 U92 ( .IN1(n8), .IN2(n130), .IN3(n140), .IN4(n50), .Q(n48) );
  AOI22X1 U93 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n46), .QN(n47) );
  OA21X1 U94 ( .IN1(n49), .IN2(n9), .IN3(n53), .Q(n54) );
  AOI22X1 U95 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n54), .QN(n52) );
  OA22X1 U96 ( .IN1(n67), .IN2(n9), .IN3(n141), .IN4(n50), .Q(n51) );
  NOR2X0 U97 ( .IN1(in2[9]), .IN2(n53), .QN(n57) );
  AO21X1 U98 ( .IN1(in2[9]), .IN2(n53), .IN3(n57), .Q(n58) );
  OA22X1 U99 ( .IN1(n9), .IN2(n130), .IN3(n140), .IN4(n58), .Q(n56) );
  AOI22X1 U100 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n54), .QN(n55) );
  OA21X1 U101 ( .IN1(n57), .IN2(n10), .IN3(n61), .Q(n62) );
  AOI22X1 U102 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n62), .QN(n60) );
  OA22X1 U103 ( .IN1(n67), .IN2(n10), .IN3(n141), .IN4(n58), .Q(n59) );
  NOR2X0 U104 ( .IN1(in2[11]), .IN2(n61), .QN(n65) );
  AO21X1 U105 ( .IN1(in2[11]), .IN2(n61), .IN3(n65), .Q(n66) );
  OA22X1 U106 ( .IN1(n10), .IN2(n130), .IN3(n140), .IN4(n66), .Q(n64) );
  AOI22X1 U107 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n62), .QN(n63) );
  OA21X1 U108 ( .IN1(n65), .IN2(n11), .IN3(n77), .Q(n70) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n70), .QN(n69) );
  OA22X1 U110 ( .IN1(n67), .IN2(n11), .IN3(n141), .IN4(n66), .Q(n68) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n12), .S(n71), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n11), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n13), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n12), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n12), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n14), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n13), .IN4(n85), .IN5(n84), 
        .Q(out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n15), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n14), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n14), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n16), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n15), .IN4(n97), .IN5(n96), 
        .Q(out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n17), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n16), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n16), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n18), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n17), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n19), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n18), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n18), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n20), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n19), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n21), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n20), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n20), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n21), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_20 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n57), .IN2(n10), .QN(n61) );
  NAND2X0 U4 ( .IN1(n33), .IN2(n7), .QN(n37) );
  NAND2X0 U5 ( .IN1(n49), .IN2(n9), .QN(n53) );
  NAND2X0 U6 ( .IN1(n41), .IN2(n8), .QN(n45) );
  NAND2X0 U7 ( .IN1(n65), .IN2(n11), .QN(n77) );
  NAND2X0 U8 ( .IN1(n81), .IN2(n13), .QN(n89) );
  NAND2X0 U9 ( .IN1(n93), .IN2(n15), .QN(n101) );
  NAND2X0 U10 ( .IN1(n105), .IN2(n17), .QN(n114) );
  NAND2X0 U11 ( .IN1(n118), .IN2(n19), .QN(n125) );
  NAND2X0 U12 ( .IN1(n25), .IN2(n6), .QN(n30) );
  NAND2X0 U13 ( .IN1(in1[2]), .IN2(n77), .QN(n71) );
  NAND2X0 U14 ( .IN1(n70), .IN2(n132), .QN(n74) );
  NAND2X0 U15 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U16 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U17 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U18 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U19 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U20 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U21 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U22 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U23 ( .IN1(n56), .IN2(n55), .QN(out1[9]) );
  NAND2X0 U24 ( .IN1(n60), .IN2(n59), .QN(out1[10]) );
  NAND2X0 U25 ( .IN1(n64), .IN2(n63), .QN(out1[11]) );
  NAND2X0 U26 ( .IN1(n69), .IN2(n68), .QN(out1[12]) );
  NAND2X0 U27 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U28 ( .IN1(n23), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U29 ( .IN1(in1[2]), .IN2(n22), .QN(n23) );
  NAND2X0 U30 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NAND2X0 U31 ( .IN1(n27), .IN2(n132), .QN(n4) );
  NAND2X0 U32 ( .IN1(n32), .IN2(n31), .QN(out1[3]) );
  NAND2X0 U33 ( .IN1(n36), .IN2(n35), .QN(out1[4]) );
  NAND2X0 U34 ( .IN1(n44), .IN2(n43), .QN(out1[6]) );
  NAND2X0 U35 ( .IN1(n40), .IN2(n39), .QN(out1[5]) );
  NAND2X0 U36 ( .IN1(n48), .IN2(n47), .QN(out1[7]) );
  NAND2X0 U37 ( .IN1(n52), .IN2(n51), .QN(out1[8]) );
  NAND2X0 U38 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U39 ( .IN1(n141), .IN2(n130), .QN(n24) );
  NOR2X0 U40 ( .IN1(n28), .IN2(n26), .QN(n3) );
  NOR2X0 U41 ( .IN1(n142), .IN2(n21), .QN(n1) );
  INVX0 U42 ( .INP(n132), .ZN(n141) );
  INVX0 U43 ( .INP(n130), .ZN(n137) );
  NAND3X0 U44 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  NOR3X0 U45 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  NOR2X0 U46 ( .IN1(n142), .IN2(n111), .QN(n138) );
  MUX21X1 U47 ( .IN1(n22), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  INVX0 U48 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U49 ( .INP(in2[2]), .ZN(n6) );
  INVX0 U50 ( .INP(in2[4]), .ZN(n7) );
  INVX0 U51 ( .INP(in2[6]), .ZN(n8) );
  INVX0 U52 ( .INP(in2[8]), .ZN(n9) );
  INVX0 U53 ( .INP(in2[10]), .ZN(n10) );
  INVX0 U54 ( .INP(in2[12]), .ZN(n11) );
  INVX0 U55 ( .INP(in2[13]), .ZN(n12) );
  INVX0 U56 ( .INP(in2[14]), .ZN(n13) );
  INVX0 U57 ( .INP(in2[15]), .ZN(n14) );
  INVX0 U58 ( .INP(in2[16]), .ZN(n15) );
  INVX0 U59 ( .INP(in2[17]), .ZN(n16) );
  INVX0 U60 ( .INP(in2[18]), .ZN(n17) );
  INVX0 U61 ( .INP(in2[19]), .ZN(n18) );
  INVX0 U62 ( .INP(in2[20]), .ZN(n19) );
  INVX0 U63 ( .INP(in2[21]), .ZN(n20) );
  INVX0 U64 ( .INP(in2[22]), .ZN(n21) );
  INVX0 U65 ( .INP(in1[1]), .ZN(n22) );
  INVX0 U66 ( .INP(in1[2]), .ZN(n111) );
  INVX0 U67 ( .INP(n138), .ZN(n140) );
  NOR2X0 U68 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n25) );
  AOI21X1 U69 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n25), .QN(n27) );
  NOR2X0 U70 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U71 ( .IN1(n24), .IN2(in2[0]), .IN3(n138), .IN4(n27), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U72 ( .INP(n133), .ZN(n67) );
  NOR2X0 U73 ( .IN1(n67), .IN2(n6), .QN(n28) );
  OA21X1 U74 ( .IN1(n25), .IN2(n6), .IN3(n30), .Q(n29) );
  AO22X1 U75 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n29), .Q(n26) );
  AOI22X1 U76 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n29), .QN(n32) );
  NOR2X0 U77 ( .IN1(in2[3]), .IN2(n30), .QN(n33) );
  AO21X1 U78 ( .IN1(in2[3]), .IN2(n30), .IN3(n33), .Q(n34) );
  OA22X1 U79 ( .IN1(n6), .IN2(n130), .IN3(n140), .IN4(n34), .Q(n31) );
  OA21X1 U80 ( .IN1(n33), .IN2(n7), .IN3(n37), .Q(n38) );
  AOI22X1 U81 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n38), .QN(n36) );
  OA22X1 U82 ( .IN1(n67), .IN2(n7), .IN3(n141), .IN4(n34), .Q(n35) );
  NOR2X0 U83 ( .IN1(in2[5]), .IN2(n37), .QN(n41) );
  AO21X1 U84 ( .IN1(in2[5]), .IN2(n37), .IN3(n41), .Q(n42) );
  OA22X1 U85 ( .IN1(n7), .IN2(n130), .IN3(n140), .IN4(n42), .Q(n40) );
  AOI22X1 U86 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n38), .QN(n39) );
  OA21X1 U87 ( .IN1(n41), .IN2(n8), .IN3(n45), .Q(n46) );
  AOI22X1 U88 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n46), .QN(n44) );
  OA22X1 U89 ( .IN1(n67), .IN2(n8), .IN3(n141), .IN4(n42), .Q(n43) );
  NOR2X0 U90 ( .IN1(in2[7]), .IN2(n45), .QN(n49) );
  AO21X1 U91 ( .IN1(in2[7]), .IN2(n45), .IN3(n49), .Q(n50) );
  OA22X1 U92 ( .IN1(n8), .IN2(n130), .IN3(n140), .IN4(n50), .Q(n48) );
  AOI22X1 U93 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n46), .QN(n47) );
  OA21X1 U94 ( .IN1(n49), .IN2(n9), .IN3(n53), .Q(n54) );
  AOI22X1 U95 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n54), .QN(n52) );
  OA22X1 U96 ( .IN1(n67), .IN2(n9), .IN3(n141), .IN4(n50), .Q(n51) );
  NOR2X0 U97 ( .IN1(in2[9]), .IN2(n53), .QN(n57) );
  AO21X1 U98 ( .IN1(in2[9]), .IN2(n53), .IN3(n57), .Q(n58) );
  OA22X1 U99 ( .IN1(n9), .IN2(n130), .IN3(n140), .IN4(n58), .Q(n56) );
  AOI22X1 U100 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n54), .QN(n55) );
  OA21X1 U101 ( .IN1(n57), .IN2(n10), .IN3(n61), .Q(n62) );
  AOI22X1 U102 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n62), .QN(n60) );
  OA22X1 U103 ( .IN1(n67), .IN2(n10), .IN3(n141), .IN4(n58), .Q(n59) );
  NOR2X0 U104 ( .IN1(in2[11]), .IN2(n61), .QN(n65) );
  AO21X1 U105 ( .IN1(in2[11]), .IN2(n61), .IN3(n65), .Q(n66) );
  OA22X1 U106 ( .IN1(n10), .IN2(n130), .IN3(n140), .IN4(n66), .Q(n64) );
  AOI22X1 U107 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n62), .QN(n63) );
  OA21X1 U108 ( .IN1(n65), .IN2(n11), .IN3(n77), .Q(n70) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n70), .QN(n69) );
  OA22X1 U110 ( .IN1(n67), .IN2(n11), .IN3(n141), .IN4(n66), .Q(n68) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n12), .S(n71), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n11), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n13), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n12), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n12), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n14), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n13), .IN4(n85), .IN5(n84), 
        .Q(out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n15), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n14), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n14), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n16), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n15), .IN4(n97), .IN5(n96), 
        .Q(out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n17), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n16), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n16), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n18), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n17), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n19), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n18), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n18), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n20), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n19), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n21), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n20), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n20), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n21), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_21 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n57), .IN2(n10), .QN(n61) );
  NAND2X0 U4 ( .IN1(n25), .IN2(n6), .QN(n30) );
  NAND2X0 U5 ( .IN1(n33), .IN2(n7), .QN(n37) );
  NAND2X0 U6 ( .IN1(n49), .IN2(n9), .QN(n53) );
  NAND2X0 U7 ( .IN1(n41), .IN2(n8), .QN(n45) );
  NAND2X0 U8 ( .IN1(n65), .IN2(n11), .QN(n77) );
  NAND2X0 U9 ( .IN1(n81), .IN2(n13), .QN(n89) );
  NAND2X0 U10 ( .IN1(n93), .IN2(n15), .QN(n101) );
  NAND2X0 U11 ( .IN1(n105), .IN2(n17), .QN(n114) );
  NAND2X0 U12 ( .IN1(in1[2]), .IN2(n77), .QN(n71) );
  NAND2X0 U13 ( .IN1(n70), .IN2(n132), .QN(n74) );
  NAND2X0 U14 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U15 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U16 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U17 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U18 ( .IN1(n118), .IN2(n19), .QN(n125) );
  NAND2X0 U19 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U20 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U21 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U22 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U23 ( .IN1(n141), .IN2(n130), .QN(n24) );
  NAND2X0 U24 ( .IN1(n27), .IN2(n132), .QN(n4) );
  NAND2X0 U25 ( .IN1(n56), .IN2(n55), .QN(out1[9]) );
  NAND2X0 U26 ( .IN1(n60), .IN2(n59), .QN(out1[10]) );
  NAND2X0 U27 ( .IN1(n64), .IN2(n63), .QN(out1[11]) );
  NAND2X0 U28 ( .IN1(n69), .IN2(n68), .QN(out1[12]) );
  NAND2X0 U29 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U30 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U31 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NAND2X0 U32 ( .IN1(n32), .IN2(n31), .QN(out1[3]) );
  NAND2X0 U33 ( .IN1(n36), .IN2(n35), .QN(out1[4]) );
  NAND2X0 U34 ( .IN1(n40), .IN2(n39), .QN(out1[5]) );
  NAND2X0 U35 ( .IN1(n44), .IN2(n43), .QN(out1[6]) );
  NAND2X0 U36 ( .IN1(n48), .IN2(n47), .QN(out1[7]) );
  NAND2X0 U37 ( .IN1(n52), .IN2(n51), .QN(out1[8]) );
  NAND2X0 U38 ( .IN1(n23), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U39 ( .IN1(in1[2]), .IN2(n22), .QN(n23) );
  NOR2X0 U40 ( .IN1(n28), .IN2(n26), .QN(n3) );
  NOR2X0 U41 ( .IN1(n142), .IN2(n21), .QN(n1) );
  INVX0 U42 ( .INP(n132), .ZN(n141) );
  INVX0 U43 ( .INP(n130), .ZN(n137) );
  NAND3X0 U44 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  NOR3X0 U45 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  NOR2X0 U46 ( .IN1(n142), .IN2(n111), .QN(n138) );
  MUX21X1 U47 ( .IN1(n22), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  INVX0 U48 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U49 ( .INP(in2[2]), .ZN(n6) );
  INVX0 U50 ( .INP(in2[4]), .ZN(n7) );
  INVX0 U51 ( .INP(in2[6]), .ZN(n8) );
  INVX0 U52 ( .INP(in2[8]), .ZN(n9) );
  INVX0 U53 ( .INP(in2[10]), .ZN(n10) );
  INVX0 U54 ( .INP(in2[12]), .ZN(n11) );
  INVX0 U55 ( .INP(in2[13]), .ZN(n12) );
  INVX0 U56 ( .INP(in2[14]), .ZN(n13) );
  INVX0 U57 ( .INP(in2[15]), .ZN(n14) );
  INVX0 U58 ( .INP(in2[16]), .ZN(n15) );
  INVX0 U59 ( .INP(in2[17]), .ZN(n16) );
  INVX0 U60 ( .INP(in2[18]), .ZN(n17) );
  INVX0 U61 ( .INP(in2[19]), .ZN(n18) );
  INVX0 U62 ( .INP(in2[20]), .ZN(n19) );
  INVX0 U63 ( .INP(in2[21]), .ZN(n20) );
  INVX0 U64 ( .INP(in2[22]), .ZN(n21) );
  INVX0 U65 ( .INP(in1[1]), .ZN(n22) );
  INVX0 U66 ( .INP(in1[2]), .ZN(n111) );
  INVX0 U67 ( .INP(n138), .ZN(n140) );
  NOR2X0 U68 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n25) );
  AOI21X1 U69 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n25), .QN(n27) );
  NOR2X0 U70 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U71 ( .IN1(n24), .IN2(in2[0]), .IN3(n138), .IN4(n27), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U72 ( .INP(n133), .ZN(n67) );
  NOR2X0 U73 ( .IN1(n67), .IN2(n6), .QN(n28) );
  OA21X1 U74 ( .IN1(n25), .IN2(n6), .IN3(n30), .Q(n29) );
  AO22X1 U75 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n29), .Q(n26) );
  AOI22X1 U76 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n29), .QN(n32) );
  NOR2X0 U77 ( .IN1(in2[3]), .IN2(n30), .QN(n33) );
  AO21X1 U78 ( .IN1(in2[3]), .IN2(n30), .IN3(n33), .Q(n34) );
  OA22X1 U79 ( .IN1(n6), .IN2(n130), .IN3(n140), .IN4(n34), .Q(n31) );
  OA21X1 U80 ( .IN1(n33), .IN2(n7), .IN3(n37), .Q(n38) );
  AOI22X1 U81 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n38), .QN(n36) );
  OA22X1 U82 ( .IN1(n67), .IN2(n7), .IN3(n141), .IN4(n34), .Q(n35) );
  NOR2X0 U83 ( .IN1(in2[5]), .IN2(n37), .QN(n41) );
  AO21X1 U84 ( .IN1(in2[5]), .IN2(n37), .IN3(n41), .Q(n42) );
  OA22X1 U85 ( .IN1(n7), .IN2(n130), .IN3(n140), .IN4(n42), .Q(n40) );
  AOI22X1 U86 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n38), .QN(n39) );
  OA21X1 U87 ( .IN1(n41), .IN2(n8), .IN3(n45), .Q(n46) );
  AOI22X1 U88 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n46), .QN(n44) );
  OA22X1 U89 ( .IN1(n67), .IN2(n8), .IN3(n141), .IN4(n42), .Q(n43) );
  NOR2X0 U90 ( .IN1(in2[7]), .IN2(n45), .QN(n49) );
  AO21X1 U91 ( .IN1(in2[7]), .IN2(n45), .IN3(n49), .Q(n50) );
  OA22X1 U92 ( .IN1(n8), .IN2(n130), .IN3(n140), .IN4(n50), .Q(n48) );
  AOI22X1 U93 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n46), .QN(n47) );
  OA21X1 U94 ( .IN1(n49), .IN2(n9), .IN3(n53), .Q(n54) );
  AOI22X1 U95 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n54), .QN(n52) );
  OA22X1 U96 ( .IN1(n67), .IN2(n9), .IN3(n141), .IN4(n50), .Q(n51) );
  NOR2X0 U97 ( .IN1(in2[9]), .IN2(n53), .QN(n57) );
  AO21X1 U98 ( .IN1(in2[9]), .IN2(n53), .IN3(n57), .Q(n58) );
  OA22X1 U99 ( .IN1(n9), .IN2(n130), .IN3(n140), .IN4(n58), .Q(n56) );
  AOI22X1 U100 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n54), .QN(n55) );
  OA21X1 U101 ( .IN1(n57), .IN2(n10), .IN3(n61), .Q(n62) );
  AOI22X1 U102 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n62), .QN(n60) );
  OA22X1 U103 ( .IN1(n67), .IN2(n10), .IN3(n141), .IN4(n58), .Q(n59) );
  NOR2X0 U104 ( .IN1(in2[11]), .IN2(n61), .QN(n65) );
  AO21X1 U105 ( .IN1(in2[11]), .IN2(n61), .IN3(n65), .Q(n66) );
  OA22X1 U106 ( .IN1(n10), .IN2(n130), .IN3(n140), .IN4(n66), .Q(n64) );
  AOI22X1 U107 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n62), .QN(n63) );
  OA21X1 U108 ( .IN1(n65), .IN2(n11), .IN3(n77), .Q(n70) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n70), .QN(n69) );
  OA22X1 U110 ( .IN1(n67), .IN2(n11), .IN3(n141), .IN4(n66), .Q(n68) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n12), .S(n71), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n11), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n13), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n12), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n12), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n14), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n13), .IN4(n85), .IN5(n84), 
        .Q(out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n15), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n14), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n14), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n16), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n15), .IN4(n97), .IN5(n96), 
        .Q(out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n17), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n16), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n16), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n18), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n17), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n19), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n18), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n18), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n20), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n19), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n21), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n20), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n20), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n21), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_22 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n25), .IN2(n6), .QN(n30) );
  NAND2X0 U4 ( .IN1(n33), .IN2(n7), .QN(n37) );
  NAND2X0 U5 ( .IN1(n41), .IN2(n8), .QN(n45) );
  NAND2X0 U6 ( .IN1(n57), .IN2(n10), .QN(n61) );
  NAND2X0 U7 ( .IN1(n49), .IN2(n9), .QN(n53) );
  NAND2X0 U8 ( .IN1(n65), .IN2(n11), .QN(n77) );
  NAND2X0 U9 ( .IN1(n81), .IN2(n13), .QN(n89) );
  NAND2X0 U10 ( .IN1(n93), .IN2(n15), .QN(n101) );
  NAND2X0 U11 ( .IN1(n105), .IN2(n17), .QN(n114) );
  NAND2X0 U12 ( .IN1(n118), .IN2(n19), .QN(n125) );
  NAND2X0 U13 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U14 ( .IN1(in1[2]), .IN2(n77), .QN(n71) );
  NAND2X0 U15 ( .IN1(n70), .IN2(n132), .QN(n74) );
  NAND2X0 U16 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U17 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U18 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U19 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U20 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U21 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U22 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U23 ( .IN1(n141), .IN2(n130), .QN(n24) );
  NAND2X0 U24 ( .IN1(n27), .IN2(n132), .QN(n4) );
  NAND2X0 U25 ( .IN1(n64), .IN2(n63), .QN(out1[11]) );
  NAND2X0 U26 ( .IN1(n69), .IN2(n68), .QN(out1[12]) );
  NAND2X0 U27 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U28 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U29 ( .IN1(n23), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U30 ( .IN1(in1[2]), .IN2(n22), .QN(n23) );
  NAND2X0 U31 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NAND2X0 U32 ( .IN1(n32), .IN2(n31), .QN(out1[3]) );
  NAND2X0 U33 ( .IN1(n36), .IN2(n35), .QN(out1[4]) );
  NAND2X0 U34 ( .IN1(n40), .IN2(n39), .QN(out1[5]) );
  NAND2X0 U35 ( .IN1(n44), .IN2(n43), .QN(out1[6]) );
  NAND2X0 U36 ( .IN1(n48), .IN2(n47), .QN(out1[7]) );
  NAND2X0 U37 ( .IN1(n52), .IN2(n51), .QN(out1[8]) );
  NAND2X0 U38 ( .IN1(n56), .IN2(n55), .QN(out1[9]) );
  NAND2X0 U39 ( .IN1(n60), .IN2(n59), .QN(out1[10]) );
  NOR2X0 U40 ( .IN1(n28), .IN2(n26), .QN(n3) );
  NOR2X0 U41 ( .IN1(n142), .IN2(n21), .QN(n1) );
  INVX0 U42 ( .INP(n132), .ZN(n141) );
  INVX0 U43 ( .INP(n130), .ZN(n137) );
  NAND3X0 U44 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  NOR3X0 U45 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  NOR2X0 U46 ( .IN1(n142), .IN2(n111), .QN(n138) );
  MUX21X1 U47 ( .IN1(n22), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  INVX0 U48 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U49 ( .INP(in2[2]), .ZN(n6) );
  INVX0 U50 ( .INP(in2[4]), .ZN(n7) );
  INVX0 U51 ( .INP(in2[6]), .ZN(n8) );
  INVX0 U52 ( .INP(in2[8]), .ZN(n9) );
  INVX0 U53 ( .INP(in2[10]), .ZN(n10) );
  INVX0 U54 ( .INP(in2[12]), .ZN(n11) );
  INVX0 U55 ( .INP(in2[13]), .ZN(n12) );
  INVX0 U56 ( .INP(in2[14]), .ZN(n13) );
  INVX0 U57 ( .INP(in2[15]), .ZN(n14) );
  INVX0 U58 ( .INP(in2[16]), .ZN(n15) );
  INVX0 U59 ( .INP(in2[17]), .ZN(n16) );
  INVX0 U60 ( .INP(in2[18]), .ZN(n17) );
  INVX0 U61 ( .INP(in2[19]), .ZN(n18) );
  INVX0 U62 ( .INP(in2[20]), .ZN(n19) );
  INVX0 U63 ( .INP(in2[21]), .ZN(n20) );
  INVX0 U64 ( .INP(in2[22]), .ZN(n21) );
  INVX0 U65 ( .INP(in1[1]), .ZN(n22) );
  INVX0 U66 ( .INP(in1[2]), .ZN(n111) );
  INVX0 U67 ( .INP(n138), .ZN(n140) );
  NOR2X0 U68 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n25) );
  AOI21X1 U69 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n25), .QN(n27) );
  NOR2X0 U70 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U71 ( .IN1(n24), .IN2(in2[0]), .IN3(n138), .IN4(n27), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U72 ( .INP(n133), .ZN(n67) );
  NOR2X0 U73 ( .IN1(n67), .IN2(n6), .QN(n28) );
  OA21X1 U74 ( .IN1(n25), .IN2(n6), .IN3(n30), .Q(n29) );
  AO22X1 U75 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n29), .Q(n26) );
  AOI22X1 U76 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n29), .QN(n32) );
  NOR2X0 U77 ( .IN1(in2[3]), .IN2(n30), .QN(n33) );
  AO21X1 U78 ( .IN1(in2[3]), .IN2(n30), .IN3(n33), .Q(n34) );
  OA22X1 U79 ( .IN1(n6), .IN2(n130), .IN3(n140), .IN4(n34), .Q(n31) );
  OA21X1 U80 ( .IN1(n33), .IN2(n7), .IN3(n37), .Q(n38) );
  AOI22X1 U81 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n38), .QN(n36) );
  OA22X1 U82 ( .IN1(n67), .IN2(n7), .IN3(n141), .IN4(n34), .Q(n35) );
  NOR2X0 U83 ( .IN1(in2[5]), .IN2(n37), .QN(n41) );
  AO21X1 U84 ( .IN1(in2[5]), .IN2(n37), .IN3(n41), .Q(n42) );
  OA22X1 U85 ( .IN1(n7), .IN2(n130), .IN3(n140), .IN4(n42), .Q(n40) );
  AOI22X1 U86 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n38), .QN(n39) );
  OA21X1 U87 ( .IN1(n41), .IN2(n8), .IN3(n45), .Q(n46) );
  AOI22X1 U88 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n46), .QN(n44) );
  OA22X1 U89 ( .IN1(n67), .IN2(n8), .IN3(n141), .IN4(n42), .Q(n43) );
  NOR2X0 U90 ( .IN1(in2[7]), .IN2(n45), .QN(n49) );
  AO21X1 U91 ( .IN1(in2[7]), .IN2(n45), .IN3(n49), .Q(n50) );
  OA22X1 U92 ( .IN1(n8), .IN2(n130), .IN3(n140), .IN4(n50), .Q(n48) );
  AOI22X1 U93 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n46), .QN(n47) );
  OA21X1 U94 ( .IN1(n49), .IN2(n9), .IN3(n53), .Q(n54) );
  AOI22X1 U95 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n54), .QN(n52) );
  OA22X1 U96 ( .IN1(n67), .IN2(n9), .IN3(n141), .IN4(n50), .Q(n51) );
  NOR2X0 U97 ( .IN1(in2[9]), .IN2(n53), .QN(n57) );
  AO21X1 U98 ( .IN1(in2[9]), .IN2(n53), .IN3(n57), .Q(n58) );
  OA22X1 U99 ( .IN1(n9), .IN2(n130), .IN3(n140), .IN4(n58), .Q(n56) );
  AOI22X1 U100 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n54), .QN(n55) );
  OA21X1 U101 ( .IN1(n57), .IN2(n10), .IN3(n61), .Q(n62) );
  AOI22X1 U102 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n62), .QN(n60) );
  OA22X1 U103 ( .IN1(n67), .IN2(n10), .IN3(n141), .IN4(n58), .Q(n59) );
  NOR2X0 U104 ( .IN1(in2[11]), .IN2(n61), .QN(n65) );
  AO21X1 U105 ( .IN1(in2[11]), .IN2(n61), .IN3(n65), .Q(n66) );
  OA22X1 U106 ( .IN1(n10), .IN2(n130), .IN3(n140), .IN4(n66), .Q(n64) );
  AOI22X1 U107 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n62), .QN(n63) );
  OA21X1 U108 ( .IN1(n65), .IN2(n11), .IN3(n77), .Q(n70) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n70), .QN(n69) );
  OA22X1 U110 ( .IN1(n67), .IN2(n11), .IN3(n141), .IN4(n66), .Q(n68) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n12), .S(n71), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n11), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n13), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n12), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n12), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n14), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n13), .IN4(n85), .IN5(n84), 
        .Q(out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n15), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n14), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n14), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n16), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n15), .IN4(n97), .IN5(n96), 
        .Q(out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n17), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n16), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n16), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n18), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n17), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n19), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n18), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n18), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n20), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n19), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n21), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n20), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n20), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n21), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_23 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n25), .IN2(n6), .QN(n30) );
  NAND2X0 U4 ( .IN1(n33), .IN2(n7), .QN(n37) );
  NAND2X0 U5 ( .IN1(n41), .IN2(n8), .QN(n45) );
  NAND2X0 U6 ( .IN1(n49), .IN2(n9), .QN(n53) );
  NAND2X0 U7 ( .IN1(n57), .IN2(n10), .QN(n61) );
  NAND2X0 U8 ( .IN1(n65), .IN2(n11), .QN(n77) );
  NAND2X0 U9 ( .IN1(n81), .IN2(n13), .QN(n89) );
  NAND2X0 U10 ( .IN1(n93), .IN2(n15), .QN(n101) );
  NAND2X0 U11 ( .IN1(n105), .IN2(n17), .QN(n114) );
  NAND2X0 U12 ( .IN1(n118), .IN2(n19), .QN(n125) );
  NAND2X0 U13 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U14 ( .IN1(in1[2]), .IN2(n77), .QN(n71) );
  NAND2X0 U15 ( .IN1(n70), .IN2(n132), .QN(n74) );
  NAND2X0 U16 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U17 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U18 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U19 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U20 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U21 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U22 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U23 ( .IN1(n23), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U24 ( .IN1(in1[2]), .IN2(n22), .QN(n23) );
  NAND2X0 U25 ( .IN1(n32), .IN2(n31), .QN(out1[3]) );
  NAND2X0 U26 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U27 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U28 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NAND2X0 U29 ( .IN1(n27), .IN2(n132), .QN(n4) );
  NAND2X0 U30 ( .IN1(n36), .IN2(n35), .QN(out1[4]) );
  NAND2X0 U31 ( .IN1(n40), .IN2(n39), .QN(out1[5]) );
  NAND2X0 U32 ( .IN1(n44), .IN2(n43), .QN(out1[6]) );
  NAND2X0 U33 ( .IN1(n48), .IN2(n47), .QN(out1[7]) );
  NAND2X0 U34 ( .IN1(n52), .IN2(n51), .QN(out1[8]) );
  NAND2X0 U35 ( .IN1(n56), .IN2(n55), .QN(out1[9]) );
  NAND2X0 U36 ( .IN1(n60), .IN2(n59), .QN(out1[10]) );
  NAND2X0 U37 ( .IN1(n64), .IN2(n63), .QN(out1[11]) );
  NAND2X0 U38 ( .IN1(n69), .IN2(n68), .QN(out1[12]) );
  NAND2X0 U39 ( .IN1(n141), .IN2(n130), .QN(n24) );
  NOR2X0 U40 ( .IN1(n28), .IN2(n26), .QN(n3) );
  NOR2X0 U41 ( .IN1(n142), .IN2(n21), .QN(n1) );
  INVX0 U42 ( .INP(n132), .ZN(n141) );
  INVX0 U43 ( .INP(n130), .ZN(n137) );
  NAND3X0 U44 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  NOR3X0 U45 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  NOR2X0 U46 ( .IN1(n142), .IN2(n111), .QN(n138) );
  MUX21X1 U47 ( .IN1(n22), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  INVX0 U48 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U49 ( .INP(in2[2]), .ZN(n6) );
  INVX0 U50 ( .INP(in2[4]), .ZN(n7) );
  INVX0 U51 ( .INP(in2[6]), .ZN(n8) );
  INVX0 U52 ( .INP(in2[8]), .ZN(n9) );
  INVX0 U53 ( .INP(in2[10]), .ZN(n10) );
  INVX0 U54 ( .INP(in2[12]), .ZN(n11) );
  INVX0 U55 ( .INP(in2[13]), .ZN(n12) );
  INVX0 U56 ( .INP(in2[14]), .ZN(n13) );
  INVX0 U57 ( .INP(in2[15]), .ZN(n14) );
  INVX0 U58 ( .INP(in2[16]), .ZN(n15) );
  INVX0 U59 ( .INP(in2[17]), .ZN(n16) );
  INVX0 U60 ( .INP(in2[18]), .ZN(n17) );
  INVX0 U61 ( .INP(in2[19]), .ZN(n18) );
  INVX0 U62 ( .INP(in2[20]), .ZN(n19) );
  INVX0 U63 ( .INP(in2[21]), .ZN(n20) );
  INVX0 U64 ( .INP(in2[22]), .ZN(n21) );
  INVX0 U65 ( .INP(in1[1]), .ZN(n22) );
  INVX0 U66 ( .INP(in1[2]), .ZN(n111) );
  INVX0 U67 ( .INP(n138), .ZN(n140) );
  NOR2X0 U68 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n25) );
  AOI21X1 U69 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n25), .QN(n27) );
  NOR2X0 U70 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U71 ( .IN1(n24), .IN2(in2[0]), .IN3(n138), .IN4(n27), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U72 ( .INP(n133), .ZN(n67) );
  NOR2X0 U73 ( .IN1(n67), .IN2(n6), .QN(n28) );
  OA21X1 U74 ( .IN1(n25), .IN2(n6), .IN3(n30), .Q(n29) );
  AO22X1 U75 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n29), .Q(n26) );
  AOI22X1 U76 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n29), .QN(n32) );
  NOR2X0 U77 ( .IN1(in2[3]), .IN2(n30), .QN(n33) );
  AO21X1 U78 ( .IN1(in2[3]), .IN2(n30), .IN3(n33), .Q(n34) );
  OA22X1 U79 ( .IN1(n6), .IN2(n130), .IN3(n140), .IN4(n34), .Q(n31) );
  OA21X1 U80 ( .IN1(n33), .IN2(n7), .IN3(n37), .Q(n38) );
  AOI22X1 U81 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n38), .QN(n36) );
  OA22X1 U82 ( .IN1(n67), .IN2(n7), .IN3(n141), .IN4(n34), .Q(n35) );
  NOR2X0 U83 ( .IN1(in2[5]), .IN2(n37), .QN(n41) );
  AO21X1 U84 ( .IN1(in2[5]), .IN2(n37), .IN3(n41), .Q(n42) );
  OA22X1 U85 ( .IN1(n7), .IN2(n130), .IN3(n140), .IN4(n42), .Q(n40) );
  AOI22X1 U86 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n38), .QN(n39) );
  OA21X1 U87 ( .IN1(n41), .IN2(n8), .IN3(n45), .Q(n46) );
  AOI22X1 U88 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n46), .QN(n44) );
  OA22X1 U89 ( .IN1(n67), .IN2(n8), .IN3(n141), .IN4(n42), .Q(n43) );
  NOR2X0 U90 ( .IN1(in2[7]), .IN2(n45), .QN(n49) );
  AO21X1 U91 ( .IN1(in2[7]), .IN2(n45), .IN3(n49), .Q(n50) );
  OA22X1 U92 ( .IN1(n8), .IN2(n130), .IN3(n140), .IN4(n50), .Q(n48) );
  AOI22X1 U93 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n46), .QN(n47) );
  OA21X1 U94 ( .IN1(n49), .IN2(n9), .IN3(n53), .Q(n54) );
  AOI22X1 U95 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n54), .QN(n52) );
  OA22X1 U96 ( .IN1(n67), .IN2(n9), .IN3(n141), .IN4(n50), .Q(n51) );
  NOR2X0 U97 ( .IN1(in2[9]), .IN2(n53), .QN(n57) );
  AO21X1 U98 ( .IN1(in2[9]), .IN2(n53), .IN3(n57), .Q(n58) );
  OA22X1 U99 ( .IN1(n9), .IN2(n130), .IN3(n140), .IN4(n58), .Q(n56) );
  AOI22X1 U100 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n54), .QN(n55) );
  OA21X1 U101 ( .IN1(n57), .IN2(n10), .IN3(n61), .Q(n62) );
  AOI22X1 U102 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n62), .QN(n60) );
  OA22X1 U103 ( .IN1(n67), .IN2(n10), .IN3(n141), .IN4(n58), .Q(n59) );
  NOR2X0 U104 ( .IN1(in2[11]), .IN2(n61), .QN(n65) );
  AO21X1 U105 ( .IN1(in2[11]), .IN2(n61), .IN3(n65), .Q(n66) );
  OA22X1 U106 ( .IN1(n10), .IN2(n130), .IN3(n140), .IN4(n66), .Q(n64) );
  AOI22X1 U107 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n62), .QN(n63) );
  OA21X1 U108 ( .IN1(n65), .IN2(n11), .IN3(n77), .Q(n70) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n70), .QN(n69) );
  OA22X1 U110 ( .IN1(n67), .IN2(n11), .IN3(n141), .IN4(n66), .Q(n68) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n12), .S(n71), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n11), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n13), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n12), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n12), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n14), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n13), .IN4(n85), .IN5(n84), 
        .Q(out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n15), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n14), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n14), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n16), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n15), .IN4(n97), .IN5(n96), 
        .Q(out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n17), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n16), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n16), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n18), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n17), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n19), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n18), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n18), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n20), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n19), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n21), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n20), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n20), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n21), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_24 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n25), .IN2(n6), .QN(n30) );
  NAND2X0 U4 ( .IN1(n33), .IN2(n7), .QN(n37) );
  NAND2X0 U5 ( .IN1(n41), .IN2(n8), .QN(n45) );
  NAND2X0 U6 ( .IN1(n49), .IN2(n9), .QN(n53) );
  NAND2X0 U7 ( .IN1(n57), .IN2(n10), .QN(n61) );
  NAND2X0 U8 ( .IN1(n65), .IN2(n11), .QN(n77) );
  NAND2X0 U9 ( .IN1(n81), .IN2(n13), .QN(n89) );
  NAND2X0 U10 ( .IN1(n105), .IN2(n17), .QN(n114) );
  NAND2X0 U11 ( .IN1(n93), .IN2(n15), .QN(n101) );
  NAND2X0 U12 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U13 ( .IN1(n118), .IN2(n19), .QN(n125) );
  NAND2X0 U14 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U15 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U16 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U17 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U18 ( .IN1(n27), .IN2(n132), .QN(n4) );
  NAND2X0 U19 ( .IN1(n141), .IN2(n130), .QN(n24) );
  NAND2X0 U20 ( .IN1(n32), .IN2(n31), .QN(out1[3]) );
  NAND2X0 U21 ( .IN1(n36), .IN2(n35), .QN(out1[4]) );
  NAND2X0 U22 ( .IN1(in1[2]), .IN2(n77), .QN(n71) );
  NAND2X0 U23 ( .IN1(n70), .IN2(n132), .QN(n74) );
  NAND2X0 U24 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U25 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U26 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U27 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U28 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NAND2X0 U29 ( .IN1(n40), .IN2(n39), .QN(out1[5]) );
  NAND2X0 U30 ( .IN1(n44), .IN2(n43), .QN(out1[6]) );
  NAND2X0 U31 ( .IN1(n48), .IN2(n47), .QN(out1[7]) );
  NAND2X0 U32 ( .IN1(n52), .IN2(n51), .QN(out1[8]) );
  NAND2X0 U33 ( .IN1(n56), .IN2(n55), .QN(out1[9]) );
  NAND2X0 U34 ( .IN1(n60), .IN2(n59), .QN(out1[10]) );
  NAND2X0 U35 ( .IN1(n64), .IN2(n63), .QN(out1[11]) );
  NAND2X0 U36 ( .IN1(n69), .IN2(n68), .QN(out1[12]) );
  NAND2X0 U37 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U38 ( .IN1(n23), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U39 ( .IN1(in1[2]), .IN2(n22), .QN(n23) );
  INVX0 U40 ( .INP(in1[2]), .ZN(n111) );
  NOR2X0 U41 ( .IN1(n28), .IN2(n26), .QN(n3) );
  INVX0 U42 ( .INP(n130), .ZN(n137) );
  INVX0 U43 ( .INP(n132), .ZN(n141) );
  NOR3X0 U44 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  NAND3X0 U45 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  NOR2X0 U46 ( .IN1(n142), .IN2(n21), .QN(n1) );
  NOR2X0 U47 ( .IN1(n142), .IN2(n111), .QN(n138) );
  MUX21X1 U48 ( .IN1(n22), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  INVX0 U49 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U50 ( .INP(in2[2]), .ZN(n6) );
  INVX0 U51 ( .INP(in2[4]), .ZN(n7) );
  INVX0 U52 ( .INP(in2[6]), .ZN(n8) );
  INVX0 U53 ( .INP(in2[8]), .ZN(n9) );
  INVX0 U54 ( .INP(in2[10]), .ZN(n10) );
  INVX0 U55 ( .INP(in2[12]), .ZN(n11) );
  INVX0 U56 ( .INP(in2[13]), .ZN(n12) );
  INVX0 U57 ( .INP(in2[14]), .ZN(n13) );
  INVX0 U58 ( .INP(in2[15]), .ZN(n14) );
  INVX0 U59 ( .INP(in2[16]), .ZN(n15) );
  INVX0 U60 ( .INP(in2[17]), .ZN(n16) );
  INVX0 U61 ( .INP(in2[18]), .ZN(n17) );
  INVX0 U62 ( .INP(in2[19]), .ZN(n18) );
  INVX0 U63 ( .INP(in2[20]), .ZN(n19) );
  INVX0 U64 ( .INP(in2[21]), .ZN(n20) );
  INVX0 U65 ( .INP(in2[22]), .ZN(n21) );
  INVX0 U66 ( .INP(in1[1]), .ZN(n22) );
  INVX0 U67 ( .INP(n138), .ZN(n140) );
  NOR2X0 U68 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n25) );
  AOI21X1 U69 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n25), .QN(n27) );
  NOR2X0 U70 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U71 ( .IN1(n24), .IN2(in2[0]), .IN3(n138), .IN4(n27), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U72 ( .INP(n133), .ZN(n67) );
  NOR2X0 U73 ( .IN1(n67), .IN2(n6), .QN(n28) );
  OA21X1 U74 ( .IN1(n25), .IN2(n6), .IN3(n30), .Q(n29) );
  AO22X1 U75 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n29), .Q(n26) );
  AOI22X1 U76 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n29), .QN(n32) );
  NOR2X0 U77 ( .IN1(in2[3]), .IN2(n30), .QN(n33) );
  AO21X1 U78 ( .IN1(in2[3]), .IN2(n30), .IN3(n33), .Q(n34) );
  OA22X1 U79 ( .IN1(n6), .IN2(n130), .IN3(n140), .IN4(n34), .Q(n31) );
  OA21X1 U80 ( .IN1(n33), .IN2(n7), .IN3(n37), .Q(n38) );
  AOI22X1 U81 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n38), .QN(n36) );
  OA22X1 U82 ( .IN1(n67), .IN2(n7), .IN3(n141), .IN4(n34), .Q(n35) );
  NOR2X0 U83 ( .IN1(in2[5]), .IN2(n37), .QN(n41) );
  AO21X1 U84 ( .IN1(in2[5]), .IN2(n37), .IN3(n41), .Q(n42) );
  OA22X1 U85 ( .IN1(n7), .IN2(n130), .IN3(n140), .IN4(n42), .Q(n40) );
  AOI22X1 U86 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n38), .QN(n39) );
  OA21X1 U87 ( .IN1(n41), .IN2(n8), .IN3(n45), .Q(n46) );
  AOI22X1 U88 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n46), .QN(n44) );
  OA22X1 U89 ( .IN1(n67), .IN2(n8), .IN3(n141), .IN4(n42), .Q(n43) );
  NOR2X0 U90 ( .IN1(in2[7]), .IN2(n45), .QN(n49) );
  AO21X1 U91 ( .IN1(in2[7]), .IN2(n45), .IN3(n49), .Q(n50) );
  OA22X1 U92 ( .IN1(n8), .IN2(n130), .IN3(n140), .IN4(n50), .Q(n48) );
  AOI22X1 U93 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n46), .QN(n47) );
  OA21X1 U94 ( .IN1(n49), .IN2(n9), .IN3(n53), .Q(n54) );
  AOI22X1 U95 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n54), .QN(n52) );
  OA22X1 U96 ( .IN1(n67), .IN2(n9), .IN3(n141), .IN4(n50), .Q(n51) );
  NOR2X0 U97 ( .IN1(in2[9]), .IN2(n53), .QN(n57) );
  AO21X1 U98 ( .IN1(in2[9]), .IN2(n53), .IN3(n57), .Q(n58) );
  OA22X1 U99 ( .IN1(n9), .IN2(n130), .IN3(n140), .IN4(n58), .Q(n56) );
  AOI22X1 U100 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n54), .QN(n55) );
  OA21X1 U101 ( .IN1(n57), .IN2(n10), .IN3(n61), .Q(n62) );
  AOI22X1 U102 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n62), .QN(n60) );
  OA22X1 U103 ( .IN1(n67), .IN2(n10), .IN3(n141), .IN4(n58), .Q(n59) );
  NOR2X0 U104 ( .IN1(in2[11]), .IN2(n61), .QN(n65) );
  AO21X1 U105 ( .IN1(in2[11]), .IN2(n61), .IN3(n65), .Q(n66) );
  OA22X1 U106 ( .IN1(n10), .IN2(n130), .IN3(n140), .IN4(n66), .Q(n64) );
  AOI22X1 U107 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n62), .QN(n63) );
  OA21X1 U108 ( .IN1(n65), .IN2(n11), .IN3(n77), .Q(n70) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n70), .QN(n69) );
  OA22X1 U110 ( .IN1(n67), .IN2(n11), .IN3(n141), .IN4(n66), .Q(n68) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n12), .S(n71), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n11), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n13), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n12), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n12), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n14), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n13), .IN4(n85), .IN5(n84), 
        .Q(out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n15), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n14), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n14), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n16), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n15), .IN4(n97), .IN5(n96), 
        .Q(out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n17), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n16), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n16), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n18), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n17), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n19), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n18), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n18), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n20), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n19), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n21), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n20), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n20), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n21), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_25 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n33), .IN2(n7), .QN(n37) );
  NAND2X0 U4 ( .IN1(n41), .IN2(n8), .QN(n45) );
  NAND2X0 U5 ( .IN1(n49), .IN2(n9), .QN(n53) );
  NAND2X0 U6 ( .IN1(n57), .IN2(n10), .QN(n61) );
  NAND2X0 U7 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U8 ( .IN1(n25), .IN2(n6), .QN(n30) );
  NAND2X0 U9 ( .IN1(n65), .IN2(n11), .QN(n77) );
  NAND2X0 U10 ( .IN1(n81), .IN2(n13), .QN(n89) );
  NAND2X0 U11 ( .IN1(n93), .IN2(n15), .QN(n101) );
  NAND2X0 U12 ( .IN1(n118), .IN2(n19), .QN(n125) );
  NAND2X0 U13 ( .IN1(n105), .IN2(n17), .QN(n114) );
  NAND2X0 U14 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U15 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U16 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U17 ( .IN1(n40), .IN2(n39), .QN(out1[5]) );
  NAND2X0 U18 ( .IN1(n44), .IN2(n43), .QN(out1[6]) );
  NAND2X0 U19 ( .IN1(in1[2]), .IN2(n77), .QN(n71) );
  NAND2X0 U20 ( .IN1(n70), .IN2(n132), .QN(n74) );
  NAND2X0 U21 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U22 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U23 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U24 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U25 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U26 ( .IN1(n23), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U27 ( .IN1(in1[2]), .IN2(n22), .QN(n23) );
  NAND2X0 U28 ( .IN1(n36), .IN2(n35), .QN(out1[4]) );
  NAND2X0 U29 ( .IN1(n32), .IN2(n31), .QN(out1[3]) );
  NAND2X0 U30 ( .IN1(n27), .IN2(n132), .QN(n4) );
  NAND2X0 U31 ( .IN1(n48), .IN2(n47), .QN(out1[7]) );
  NAND2X0 U32 ( .IN1(n52), .IN2(n51), .QN(out1[8]) );
  NAND2X0 U33 ( .IN1(n56), .IN2(n55), .QN(out1[9]) );
  NAND2X0 U34 ( .IN1(n60), .IN2(n59), .QN(out1[10]) );
  NAND2X0 U35 ( .IN1(n64), .IN2(n63), .QN(out1[11]) );
  NAND2X0 U36 ( .IN1(n69), .IN2(n68), .QN(out1[12]) );
  NAND2X0 U37 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U38 ( .IN1(n141), .IN2(n130), .QN(n24) );
  NAND2X0 U39 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NOR2X0 U40 ( .IN1(n28), .IN2(n26), .QN(n3) );
  NOR2X0 U41 ( .IN1(n142), .IN2(n21), .QN(n1) );
  INVX0 U42 ( .INP(n132), .ZN(n141) );
  INVX0 U43 ( .INP(n130), .ZN(n137) );
  NAND3X0 U44 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  NOR2X0 U45 ( .IN1(n142), .IN2(n111), .QN(n138) );
  MUX21X1 U46 ( .IN1(n22), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  NOR3X0 U47 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  INVX0 U48 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U49 ( .INP(in2[2]), .ZN(n6) );
  INVX0 U50 ( .INP(in2[4]), .ZN(n7) );
  INVX0 U51 ( .INP(in2[6]), .ZN(n8) );
  INVX0 U52 ( .INP(in2[8]), .ZN(n9) );
  INVX0 U53 ( .INP(in2[10]), .ZN(n10) );
  INVX0 U54 ( .INP(in2[12]), .ZN(n11) );
  INVX0 U55 ( .INP(in2[13]), .ZN(n12) );
  INVX0 U56 ( .INP(in2[14]), .ZN(n13) );
  INVX0 U57 ( .INP(in2[15]), .ZN(n14) );
  INVX0 U58 ( .INP(in2[16]), .ZN(n15) );
  INVX0 U59 ( .INP(in2[17]), .ZN(n16) );
  INVX0 U60 ( .INP(in2[18]), .ZN(n17) );
  INVX0 U61 ( .INP(in2[19]), .ZN(n18) );
  INVX0 U62 ( .INP(in2[20]), .ZN(n19) );
  INVX0 U63 ( .INP(in2[21]), .ZN(n20) );
  INVX0 U64 ( .INP(in2[22]), .ZN(n21) );
  INVX0 U65 ( .INP(in1[1]), .ZN(n22) );
  INVX0 U66 ( .INP(in1[2]), .ZN(n111) );
  INVX0 U67 ( .INP(n138), .ZN(n140) );
  NOR2X0 U68 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n25) );
  AOI21X1 U69 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n25), .QN(n27) );
  NOR2X0 U70 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U71 ( .IN1(n24), .IN2(in2[0]), .IN3(n138), .IN4(n27), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U72 ( .INP(n133), .ZN(n67) );
  NOR2X0 U73 ( .IN1(n67), .IN2(n6), .QN(n28) );
  OA21X1 U74 ( .IN1(n25), .IN2(n6), .IN3(n30), .Q(n29) );
  AO22X1 U75 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n29), .Q(n26) );
  AOI22X1 U76 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n29), .QN(n32) );
  NOR2X0 U77 ( .IN1(in2[3]), .IN2(n30), .QN(n33) );
  AO21X1 U78 ( .IN1(in2[3]), .IN2(n30), .IN3(n33), .Q(n34) );
  OA22X1 U79 ( .IN1(n6), .IN2(n130), .IN3(n140), .IN4(n34), .Q(n31) );
  OA21X1 U80 ( .IN1(n33), .IN2(n7), .IN3(n37), .Q(n38) );
  AOI22X1 U81 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n38), .QN(n36) );
  OA22X1 U82 ( .IN1(n67), .IN2(n7), .IN3(n141), .IN4(n34), .Q(n35) );
  NOR2X0 U83 ( .IN1(in2[5]), .IN2(n37), .QN(n41) );
  AO21X1 U84 ( .IN1(in2[5]), .IN2(n37), .IN3(n41), .Q(n42) );
  OA22X1 U85 ( .IN1(n7), .IN2(n130), .IN3(n140), .IN4(n42), .Q(n40) );
  AOI22X1 U86 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n38), .QN(n39) );
  OA21X1 U87 ( .IN1(n41), .IN2(n8), .IN3(n45), .Q(n46) );
  AOI22X1 U88 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n46), .QN(n44) );
  OA22X1 U89 ( .IN1(n67), .IN2(n8), .IN3(n141), .IN4(n42), .Q(n43) );
  NOR2X0 U90 ( .IN1(in2[7]), .IN2(n45), .QN(n49) );
  AO21X1 U91 ( .IN1(in2[7]), .IN2(n45), .IN3(n49), .Q(n50) );
  OA22X1 U92 ( .IN1(n8), .IN2(n130), .IN3(n140), .IN4(n50), .Q(n48) );
  AOI22X1 U93 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n46), .QN(n47) );
  OA21X1 U94 ( .IN1(n49), .IN2(n9), .IN3(n53), .Q(n54) );
  AOI22X1 U95 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n54), .QN(n52) );
  OA22X1 U96 ( .IN1(n67), .IN2(n9), .IN3(n141), .IN4(n50), .Q(n51) );
  NOR2X0 U97 ( .IN1(in2[9]), .IN2(n53), .QN(n57) );
  AO21X1 U98 ( .IN1(in2[9]), .IN2(n53), .IN3(n57), .Q(n58) );
  OA22X1 U99 ( .IN1(n9), .IN2(n130), .IN3(n140), .IN4(n58), .Q(n56) );
  AOI22X1 U100 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n54), .QN(n55) );
  OA21X1 U101 ( .IN1(n57), .IN2(n10), .IN3(n61), .Q(n62) );
  AOI22X1 U102 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n62), .QN(n60) );
  OA22X1 U103 ( .IN1(n67), .IN2(n10), .IN3(n141), .IN4(n58), .Q(n59) );
  NOR2X0 U104 ( .IN1(in2[11]), .IN2(n61), .QN(n65) );
  AO21X1 U105 ( .IN1(in2[11]), .IN2(n61), .IN3(n65), .Q(n66) );
  OA22X1 U106 ( .IN1(n10), .IN2(n130), .IN3(n140), .IN4(n66), .Q(n64) );
  AOI22X1 U107 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n62), .QN(n63) );
  OA21X1 U108 ( .IN1(n65), .IN2(n11), .IN3(n77), .Q(n70) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n70), .QN(n69) );
  OA22X1 U110 ( .IN1(n67), .IN2(n11), .IN3(n141), .IN4(n66), .Q(n68) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n12), .S(n71), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n11), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n13), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n12), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n12), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n14), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n13), .IN4(n85), .IN5(n84), 
        .Q(out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n15), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n14), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n14), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n16), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n15), .IN4(n97), .IN5(n96), 
        .Q(out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n17), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n16), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n16), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n18), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n17), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n19), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n18), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n18), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n20), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n19), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n21), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n20), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n20), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n21), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_26 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93;

  NAND2X0 U3 ( .IN1(n30), .IN2(n7), .QN(n32) );
  NAND2X0 U4 ( .IN1(n34), .IN2(n8), .QN(n36) );
  NAND2X0 U5 ( .IN1(n38), .IN2(n9), .QN(n40) );
  NAND2X0 U6 ( .IN1(n42), .IN2(n10), .QN(n47) );
  NAND2X0 U7 ( .IN1(n78), .IN2(n18), .QN(n82) );
  NAND2X0 U8 ( .IN1(n26), .IN2(n6), .QN(n28) );
  NAND2X0 U9 ( .IN1(in1[2]), .IN2(n47), .QN(n44) );
  NAND2X0 U10 ( .IN1(n52), .IN2(n12), .QN(n55) );
  NAND2X0 U11 ( .IN1(in1[2]), .IN2(n55), .QN(n51) );
  NAND2X0 U12 ( .IN1(n60), .IN2(n14), .QN(n63) );
  NAND2X0 U13 ( .IN1(in1[2]), .IN2(n63), .QN(n59) );
  NAND2X0 U14 ( .IN1(n68), .IN2(n16), .QN(n71) );
  NAND2X0 U15 ( .IN1(in1[2]), .IN2(n71), .QN(n67) );
  NAND2X0 U16 ( .IN1(in1[2]), .IN2(n82), .QN(n77) );
  NAND2X0 U17 ( .IN1(in2[21]), .IN2(n82), .QN(n83) );
  NAND2X0 U18 ( .IN1(n75), .IN2(in1[2]), .QN(n86) );
  NAND2X0 U19 ( .IN1(n3), .IN2(n4), .QN(n22) );
  NAND2X0 U20 ( .IN1(n23), .IN2(n22), .QN(out1[2]) );
  INVX0 U21 ( .INP(n86), .ZN(n89) );
  NAND2X0 U22 ( .IN1(in2[1]), .IN2(in2[0]), .QN(n4) );
  NOR2X0 U23 ( .IN1(n21), .IN2(n86), .QN(n3) );
  NOR2X0 U24 ( .IN1(in1[2]), .IN2(n75), .QN(n90) );
  NBUFFX2 U25 ( .INP(in1[2]), .Z(out1[25]) );
  NOR2X0 U26 ( .IN1(n75), .IN2(n72), .QN(n92) );
  NBUFFX2 U27 ( .INP(in1[2]), .Z(out1[26]) );
  INVX0 U28 ( .INP(in2[2]), .ZN(n5) );
  INVX0 U29 ( .INP(in2[4]), .ZN(n6) );
  INVX0 U30 ( .INP(in2[6]), .ZN(n7) );
  INVX0 U31 ( .INP(in2[8]), .ZN(n8) );
  INVX0 U32 ( .INP(in2[10]), .ZN(n9) );
  INVX0 U33 ( .INP(in2[12]), .ZN(n10) );
  INVX0 U34 ( .INP(in2[13]), .ZN(n11) );
  INVX0 U35 ( .INP(in2[14]), .ZN(n12) );
  INVX0 U36 ( .INP(in2[15]), .ZN(n13) );
  INVX0 U37 ( .INP(in2[16]), .ZN(n14) );
  INVX0 U38 ( .INP(in2[17]), .ZN(n15) );
  INVX0 U39 ( .INP(in2[18]), .ZN(n16) );
  INVX0 U40 ( .INP(in2[19]), .ZN(n17) );
  INVX0 U41 ( .INP(in2[20]), .ZN(n18) );
  INVX0 U42 ( .INP(in2[21]), .ZN(n19) );
  INVX0 U43 ( .INP(in2[22]), .ZN(n20) );
  INVX0 U44 ( .INP(in1[1]), .ZN(n75) );
  INVX0 U45 ( .INP(in1[2]), .ZN(n72) );
  NOR2X0 U46 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n21) );
  OR3X1 U47 ( .IN1(in2[2]), .IN2(in2[0]), .IN3(in2[1]), .Q(n24) );
  OA21X1 U48 ( .IN1(n21), .IN2(n5), .IN3(n24), .Q(n25) );
  AOI22X1 U49 ( .IN1(in2[2]), .IN2(n90), .IN3(n92), .IN4(n25), .QN(n23) );
  NOR2X0 U50 ( .IN1(in2[3]), .IN2(n24), .QN(n26) );
  AOI21X1 U51 ( .IN1(in2[3]), .IN2(n24), .IN3(n26), .QN(n27) );
  AO222X1 U52 ( .IN1(in2[3]), .IN2(n90), .IN3(n92), .IN4(n27), .IN5(n89), 
        .IN6(n25), .Q(out1[3]) );
  OA21X1 U53 ( .IN1(n26), .IN2(n6), .IN3(n28), .Q(n29) );
  AO222X1 U54 ( .IN1(in2[4]), .IN2(n90), .IN3(n92), .IN4(n29), .IN5(n89), 
        .IN6(n27), .Q(out1[4]) );
  NOR2X0 U55 ( .IN1(in2[5]), .IN2(n28), .QN(n30) );
  AOI21X1 U56 ( .IN1(in2[5]), .IN2(n28), .IN3(n30), .QN(n31) );
  AO222X1 U57 ( .IN1(in2[5]), .IN2(n90), .IN3(n92), .IN4(n31), .IN5(n89), 
        .IN6(n29), .Q(out1[5]) );
  OA21X1 U58 ( .IN1(n30), .IN2(n7), .IN3(n32), .Q(n33) );
  AO222X1 U59 ( .IN1(in2[6]), .IN2(n90), .IN3(n92), .IN4(n33), .IN5(n89), 
        .IN6(n31), .Q(out1[6]) );
  NOR2X0 U60 ( .IN1(in2[7]), .IN2(n32), .QN(n34) );
  AOI21X1 U61 ( .IN1(in2[7]), .IN2(n32), .IN3(n34), .QN(n35) );
  AO222X1 U62 ( .IN1(in2[7]), .IN2(n90), .IN3(n92), .IN4(n35), .IN5(n89), 
        .IN6(n33), .Q(out1[7]) );
  OA21X1 U63 ( .IN1(n34), .IN2(n8), .IN3(n36), .Q(n37) );
  AO222X1 U64 ( .IN1(in2[8]), .IN2(n90), .IN3(n92), .IN4(n37), .IN5(n89), 
        .IN6(n35), .Q(out1[8]) );
  NOR2X0 U65 ( .IN1(in2[9]), .IN2(n36), .QN(n38) );
  AOI21X1 U66 ( .IN1(in2[9]), .IN2(n36), .IN3(n38), .QN(n39) );
  AO222X1 U67 ( .IN1(in2[9]), .IN2(n90), .IN3(n92), .IN4(n39), .IN5(n89), 
        .IN6(n37), .Q(out1[9]) );
  OA21X1 U68 ( .IN1(n38), .IN2(n9), .IN3(n40), .Q(n41) );
  AO222X1 U69 ( .IN1(in2[10]), .IN2(n90), .IN3(n92), .IN4(n41), .IN5(n89), 
        .IN6(n39), .Q(out1[10]) );
  NOR2X0 U70 ( .IN1(in2[11]), .IN2(n40), .QN(n42) );
  AOI21X1 U71 ( .IN1(in2[11]), .IN2(n40), .IN3(n42), .QN(n43) );
  AO222X1 U72 ( .IN1(in2[11]), .IN2(n90), .IN3(n92), .IN4(n43), .IN5(n89), 
        .IN6(n41), .Q(out1[11]) );
  OA21X1 U73 ( .IN1(n42), .IN2(n10), .IN3(n47), .Q(n45) );
  AO222X1 U74 ( .IN1(in2[12]), .IN2(n90), .IN3(n92), .IN4(n45), .IN5(n89), 
        .IN6(n43), .Q(out1[12]) );
  MUX21X1 U75 ( .IN1(n11), .IN2(in2[13]), .S(n44), .Q(n46) );
  AO22X1 U76 ( .IN1(in1[1]), .IN2(n46), .IN3(n89), .IN4(n45), .Q(out1[13]) );
  NOR2X0 U77 ( .IN1(in2[13]), .IN2(n47), .QN(n52) );
  AO21X1 U78 ( .IN1(in2[13]), .IN2(n47), .IN3(n86), .Q(n50) );
  NOR2X0 U79 ( .IN1(n52), .IN2(n72), .QN(n48) );
  MUX21X1 U80 ( .IN1(n12), .IN2(in2[14]), .S(n48), .Q(n49) );
  OAI22X1 U81 ( .IN1(n52), .IN2(n50), .IN3(n75), .IN4(n49), .QN(out1[14]) );
  MUX21X1 U82 ( .IN1(n13), .IN2(in2[15]), .S(n51), .Q(n54) );
  OA21X1 U83 ( .IN1(n52), .IN2(n12), .IN3(n89), .Q(n53) );
  AO22X1 U84 ( .IN1(in1[1]), .IN2(n54), .IN3(n53), .IN4(n55), .Q(out1[15]) );
  NOR2X0 U85 ( .IN1(in2[15]), .IN2(n55), .QN(n60) );
  AO21X1 U86 ( .IN1(in2[15]), .IN2(n55), .IN3(n86), .Q(n58) );
  NOR2X0 U87 ( .IN1(n60), .IN2(n72), .QN(n56) );
  MUX21X1 U88 ( .IN1(n14), .IN2(in2[16]), .S(n56), .Q(n57) );
  OAI22X1 U89 ( .IN1(n60), .IN2(n58), .IN3(n75), .IN4(n57), .QN(out1[16]) );
  MUX21X1 U90 ( .IN1(n15), .IN2(in2[17]), .S(n59), .Q(n62) );
  OA21X1 U91 ( .IN1(n60), .IN2(n14), .IN3(n89), .Q(n61) );
  AO22X1 U92 ( .IN1(in1[1]), .IN2(n62), .IN3(n61), .IN4(n63), .Q(out1[17]) );
  NOR2X0 U93 ( .IN1(in2[17]), .IN2(n63), .QN(n68) );
  AO21X1 U94 ( .IN1(in2[17]), .IN2(n63), .IN3(n86), .Q(n66) );
  NOR2X0 U95 ( .IN1(n68), .IN2(n72), .QN(n64) );
  MUX21X1 U96 ( .IN1(n16), .IN2(in2[18]), .S(n64), .Q(n65) );
  OAI22X1 U97 ( .IN1(n68), .IN2(n66), .IN3(n75), .IN4(n65), .QN(out1[18]) );
  MUX21X1 U98 ( .IN1(n17), .IN2(in2[19]), .S(n67), .Q(n70) );
  OA21X1 U99 ( .IN1(n68), .IN2(n16), .IN3(n89), .Q(n69) );
  AO22X1 U100 ( .IN1(in1[1]), .IN2(n70), .IN3(n69), .IN4(n71), .Q(out1[19]) );
  NOR2X0 U101 ( .IN1(in2[19]), .IN2(n71), .QN(n78) );
  AO21X1 U102 ( .IN1(in2[19]), .IN2(n71), .IN3(n86), .Q(n76) );
  NOR2X0 U103 ( .IN1(n78), .IN2(n72), .QN(n73) );
  MUX21X1 U104 ( .IN1(n18), .IN2(in2[20]), .S(n73), .Q(n74) );
  OAI22X1 U105 ( .IN1(n78), .IN2(n76), .IN3(n75), .IN4(n74), .QN(out1[20]) );
  MUX21X1 U106 ( .IN1(n19), .IN2(in2[21]), .S(n77), .Q(n80) );
  MUX21X1 U107 ( .IN1(n18), .IN2(in2[20]), .S(n78), .Q(n79) );
  AO22X1 U108 ( .IN1(in1[1]), .IN2(n80), .IN3(n89), .IN4(n79), .Q(out1[21]) );
  INVX0 U109 ( .INP(n92), .ZN(n81) );
  OR2X1 U110 ( .IN1(n82), .IN2(in2[21]), .Q(n88) );
  NOR2X0 U111 ( .IN1(n81), .IN2(n88), .QN(n87) );
  NOR2X0 U112 ( .IN1(in2[22]), .IN2(n81), .QN(n84) );
  OA221X1 U113 ( .IN1(n84), .IN2(n89), .IN3(n84), .IN4(n83), .IN5(n88), .Q(n85) );
  AO221X1 U114 ( .IN1(in2[22]), .IN2(n87), .IN3(in2[22]), .IN4(n90), .IN5(n85), 
        .Q(out1[22]) );
  NOR2X0 U115 ( .IN1(n86), .IN2(n88), .QN(n93) );
  AO21X1 U116 ( .IN1(n89), .IN2(n88), .IN3(n87), .Q(n91) );
  AO221X1 U117 ( .IN1(in2[22]), .IN2(n93), .IN3(n20), .IN4(n91), .IN5(n90), 
        .Q(out1[23]) );
  AO21X1 U118 ( .IN1(n93), .IN2(n20), .IN3(n92), .Q(out1[24]) );
endmodule


module mul26_2 ( clk, rst_n, in1, in2, en, mulout );
  input [25:0] in1;
  input [25:0] in2;
  output [50:0] mulout;
  input clk, rst_n, en;
  wire   N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24,
         N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38,
         N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N62, N63,
         N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77,
         N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91,
         N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n130, n131, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22,
         SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24,
         SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26,
         SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28,
         SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30,
         SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32,
         SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34,
         SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36,
         SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38,
         SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40,
         SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42,
         SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44,
         SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46,
         SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48,
         SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50,
         SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52,
         SYNOPSYS_UNCONNECTED_53, SYNOPSYS_UNCONNECTED_54,
         SYNOPSYS_UNCONNECTED_55, SYNOPSYS_UNCONNECTED_56,
         SYNOPSYS_UNCONNECTED_57, SYNOPSYS_UNCONNECTED_58,
         SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_60,
         SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_62,
         SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_64,
         SYNOPSYS_UNCONNECTED_65, SYNOPSYS_UNCONNECTED_66,
         SYNOPSYS_UNCONNECTED_67, SYNOPSYS_UNCONNECTED_68,
         SYNOPSYS_UNCONNECTED_69, SYNOPSYS_UNCONNECTED_70,
         SYNOPSYS_UNCONNECTED_71, SYNOPSYS_UNCONNECTED_72,
         SYNOPSYS_UNCONNECTED_73, SYNOPSYS_UNCONNECTED_74,
         SYNOPSYS_UNCONNECTED_75, SYNOPSYS_UNCONNECTED_76,
         SYNOPSYS_UNCONNECTED_77, SYNOPSYS_UNCONNECTED_78,
         SYNOPSYS_UNCONNECTED_79, SYNOPSYS_UNCONNECTED_80,
         SYNOPSYS_UNCONNECTED_81, SYNOPSYS_UNCONNECTED_82,
         SYNOPSYS_UNCONNECTED_83, SYNOPSYS_UNCONNECTED_84,
         SYNOPSYS_UNCONNECTED_85, SYNOPSYS_UNCONNECTED_86,
         SYNOPSYS_UNCONNECTED_87, SYNOPSYS_UNCONNECTED_88,
         SYNOPSYS_UNCONNECTED_89, SYNOPSYS_UNCONNECTED_90,
         SYNOPSYS_UNCONNECTED_91, SYNOPSYS_UNCONNECTED_92,
         SYNOPSYS_UNCONNECTED_93, SYNOPSYS_UNCONNECTED_94,
         SYNOPSYS_UNCONNECTED_95, SYNOPSYS_UNCONNECTED_96,
         SYNOPSYS_UNCONNECTED_97, SYNOPSYS_UNCONNECTED_98,
         SYNOPSYS_UNCONNECTED_99, SYNOPSYS_UNCONNECTED_100,
         SYNOPSYS_UNCONNECTED_101, SYNOPSYS_UNCONNECTED_102,
         SYNOPSYS_UNCONNECTED_103, SYNOPSYS_UNCONNECTED_104,
         SYNOPSYS_UNCONNECTED_105, SYNOPSYS_UNCONNECTED_106,
         SYNOPSYS_UNCONNECTED_107, SYNOPSYS_UNCONNECTED_108,
         SYNOPSYS_UNCONNECTED_109, SYNOPSYS_UNCONNECTED_110,
         SYNOPSYS_UNCONNECTED_111, SYNOPSYS_UNCONNECTED_112,
         SYNOPSYS_UNCONNECTED_113, SYNOPSYS_UNCONNECTED_114,
         SYNOPSYS_UNCONNECTED_115, SYNOPSYS_UNCONNECTED_116,
         SYNOPSYS_UNCONNECTED_117, SYNOPSYS_UNCONNECTED_118,
         SYNOPSYS_UNCONNECTED_119, SYNOPSYS_UNCONNECTED_120,
         SYNOPSYS_UNCONNECTED_121, SYNOPSYS_UNCONNECTED_122,
         SYNOPSYS_UNCONNECTED_123, SYNOPSYS_UNCONNECTED_124,
         SYNOPSYS_UNCONNECTED_125, SYNOPSYS_UNCONNECTED_126,
         SYNOPSYS_UNCONNECTED_127, SYNOPSYS_UNCONNECTED_128,
         SYNOPSYS_UNCONNECTED_129, SYNOPSYS_UNCONNECTED_130,
         SYNOPSYS_UNCONNECTED_131, SYNOPSYS_UNCONNECTED_132,
         SYNOPSYS_UNCONNECTED_133, SYNOPSYS_UNCONNECTED_134,
         SYNOPSYS_UNCONNECTED_135, SYNOPSYS_UNCONNECTED_136,
         SYNOPSYS_UNCONNECTED_137, SYNOPSYS_UNCONNECTED_138,
         SYNOPSYS_UNCONNECTED_139, SYNOPSYS_UNCONNECTED_140,
         SYNOPSYS_UNCONNECTED_141, SYNOPSYS_UNCONNECTED_142,
         SYNOPSYS_UNCONNECTED_143, SYNOPSYS_UNCONNECTED_144,
         SYNOPSYS_UNCONNECTED_145, SYNOPSYS_UNCONNECTED_146,
         SYNOPSYS_UNCONNECTED_147, SYNOPSYS_UNCONNECTED_148,
         SYNOPSYS_UNCONNECTED_149, SYNOPSYS_UNCONNECTED_150,
         SYNOPSYS_UNCONNECTED_151, SYNOPSYS_UNCONNECTED_152,
         SYNOPSYS_UNCONNECTED_153, SYNOPSYS_UNCONNECTED_154,
         SYNOPSYS_UNCONNECTED_155, SYNOPSYS_UNCONNECTED_156,
         SYNOPSYS_UNCONNECTED_157, SYNOPSYS_UNCONNECTED_158,
         SYNOPSYS_UNCONNECTED_159, SYNOPSYS_UNCONNECTED_160,
         SYNOPSYS_UNCONNECTED_161, SYNOPSYS_UNCONNECTED_162,
         SYNOPSYS_UNCONNECTED_163, SYNOPSYS_UNCONNECTED_164,
         SYNOPSYS_UNCONNECTED_165, SYNOPSYS_UNCONNECTED_166,
         SYNOPSYS_UNCONNECTED_167, SYNOPSYS_UNCONNECTED_168,
         SYNOPSYS_UNCONNECTED_169, SYNOPSYS_UNCONNECTED_170,
         SYNOPSYS_UNCONNECTED_171, SYNOPSYS_UNCONNECTED_172,
         SYNOPSYS_UNCONNECTED_173, SYNOPSYS_UNCONNECTED_174,
         SYNOPSYS_UNCONNECTED_175, SYNOPSYS_UNCONNECTED_176,
         SYNOPSYS_UNCONNECTED_177, SYNOPSYS_UNCONNECTED_178,
         SYNOPSYS_UNCONNECTED_179, SYNOPSYS_UNCONNECTED_180,
         SYNOPSYS_UNCONNECTED_181, SYNOPSYS_UNCONNECTED_182,
         SYNOPSYS_UNCONNECTED_183, SYNOPSYS_UNCONNECTED_184,
         SYNOPSYS_UNCONNECTED_185, SYNOPSYS_UNCONNECTED_186,
         SYNOPSYS_UNCONNECTED_187, SYNOPSYS_UNCONNECTED_188,
         SYNOPSYS_UNCONNECTED_189, SYNOPSYS_UNCONNECTED_190,
         SYNOPSYS_UNCONNECTED_191, SYNOPSYS_UNCONNECTED_192,
         SYNOPSYS_UNCONNECTED_193, SYNOPSYS_UNCONNECTED_194,
         SYNOPSYS_UNCONNECTED_195, SYNOPSYS_UNCONNECTED_196,
         SYNOPSYS_UNCONNECTED_197, SYNOPSYS_UNCONNECTED_198,
         SYNOPSYS_UNCONNECTED_199, SYNOPSYS_UNCONNECTED_200,
         SYNOPSYS_UNCONNECTED_201, SYNOPSYS_UNCONNECTED_202,
         SYNOPSYS_UNCONNECTED_203, SYNOPSYS_UNCONNECTED_204,
         SYNOPSYS_UNCONNECTED_205, SYNOPSYS_UNCONNECTED_206,
         SYNOPSYS_UNCONNECTED_207, SYNOPSYS_UNCONNECTED_208,
         SYNOPSYS_UNCONNECTED_209, SYNOPSYS_UNCONNECTED_210,
         SYNOPSYS_UNCONNECTED_211, SYNOPSYS_UNCONNECTED_212,
         SYNOPSYS_UNCONNECTED_213, SYNOPSYS_UNCONNECTED_214,
         SYNOPSYS_UNCONNECTED_215, SYNOPSYS_UNCONNECTED_216,
         SYNOPSYS_UNCONNECTED_217, SYNOPSYS_UNCONNECTED_218,
         SYNOPSYS_UNCONNECTED_219, SYNOPSYS_UNCONNECTED_220,
         SYNOPSYS_UNCONNECTED_221, SYNOPSYS_UNCONNECTED_222,
         SYNOPSYS_UNCONNECTED_223, SYNOPSYS_UNCONNECTED_224,
         SYNOPSYS_UNCONNECTED_225, SYNOPSYS_UNCONNECTED_226,
         SYNOPSYS_UNCONNECTED_227, SYNOPSYS_UNCONNECTED_228,
         SYNOPSYS_UNCONNECTED_229, SYNOPSYS_UNCONNECTED_230,
         SYNOPSYS_UNCONNECTED_231, SYNOPSYS_UNCONNECTED_232,
         SYNOPSYS_UNCONNECTED_233, SYNOPSYS_UNCONNECTED_234,
         SYNOPSYS_UNCONNECTED_235, SYNOPSYS_UNCONNECTED_236,
         SYNOPSYS_UNCONNECTED_237, SYNOPSYS_UNCONNECTED_238,
         SYNOPSYS_UNCONNECTED_239, SYNOPSYS_UNCONNECTED_240,
         SYNOPSYS_UNCONNECTED_241, SYNOPSYS_UNCONNECTED_242,
         SYNOPSYS_UNCONNECTED_243, SYNOPSYS_UNCONNECTED_244,
         SYNOPSYS_UNCONNECTED_245, SYNOPSYS_UNCONNECTED_246,
         SYNOPSYS_UNCONNECTED_247, SYNOPSYS_UNCONNECTED_248,
         SYNOPSYS_UNCONNECTED_249, SYNOPSYS_UNCONNECTED_250,
         SYNOPSYS_UNCONNECTED_251, SYNOPSYS_UNCONNECTED_252,
         SYNOPSYS_UNCONNECTED_253, SYNOPSYS_UNCONNECTED_254,
         SYNOPSYS_UNCONNECTED_255, SYNOPSYS_UNCONNECTED_256,
         SYNOPSYS_UNCONNECTED_257, SYNOPSYS_UNCONNECTED_258,
         SYNOPSYS_UNCONNECTED_259, SYNOPSYS_UNCONNECTED_260,
         SYNOPSYS_UNCONNECTED_261, SYNOPSYS_UNCONNECTED_262,
         SYNOPSYS_UNCONNECTED_263, SYNOPSYS_UNCONNECTED_264,
         SYNOPSYS_UNCONNECTED_265, SYNOPSYS_UNCONNECTED_266,
         SYNOPSYS_UNCONNECTED_267, SYNOPSYS_UNCONNECTED_268,
         SYNOPSYS_UNCONNECTED_269, SYNOPSYS_UNCONNECTED_270,
         SYNOPSYS_UNCONNECTED_271, SYNOPSYS_UNCONNECTED_272,
         SYNOPSYS_UNCONNECTED_273, SYNOPSYS_UNCONNECTED_274,
         SYNOPSYS_UNCONNECTED_275, SYNOPSYS_UNCONNECTED_276,
         SYNOPSYS_UNCONNECTED_277, SYNOPSYS_UNCONNECTED_278,
         SYNOPSYS_UNCONNECTED_279, SYNOPSYS_UNCONNECTED_280,
         SYNOPSYS_UNCONNECTED_281, SYNOPSYS_UNCONNECTED_282,
         SYNOPSYS_UNCONNECTED_283, SYNOPSYS_UNCONNECTED_284,
         SYNOPSYS_UNCONNECTED_285, SYNOPSYS_UNCONNECTED_286,
         SYNOPSYS_UNCONNECTED_287, SYNOPSYS_UNCONNECTED_288,
         SYNOPSYS_UNCONNECTED_289, SYNOPSYS_UNCONNECTED_290,
         SYNOPSYS_UNCONNECTED_291, SYNOPSYS_UNCONNECTED_292,
         SYNOPSYS_UNCONNECTED_293, SYNOPSYS_UNCONNECTED_294,
         SYNOPSYS_UNCONNECTED_295, SYNOPSYS_UNCONNECTED_296,
         SYNOPSYS_UNCONNECTED_297, SYNOPSYS_UNCONNECTED_298,
         SYNOPSYS_UNCONNECTED_299, SYNOPSYS_UNCONNECTED_300,
         SYNOPSYS_UNCONNECTED_301, SYNOPSYS_UNCONNECTED_302,
         SYNOPSYS_UNCONNECTED_303, SYNOPSYS_UNCONNECTED_304,
         SYNOPSYS_UNCONNECTED_305, SYNOPSYS_UNCONNECTED_306,
         SYNOPSYS_UNCONNECTED_307, SYNOPSYS_UNCONNECTED_308,
         SYNOPSYS_UNCONNECTED_309, SYNOPSYS_UNCONNECTED_310,
         SYNOPSYS_UNCONNECTED_311, SYNOPSYS_UNCONNECTED_312,
         SYNOPSYS_UNCONNECTED_313, SYNOPSYS_UNCONNECTED_314,
         SYNOPSYS_UNCONNECTED_315, SYNOPSYS_UNCONNECTED_316,
         SYNOPSYS_UNCONNECTED_317, SYNOPSYS_UNCONNECTED_318,
         SYNOPSYS_UNCONNECTED_319, SYNOPSYS_UNCONNECTED_320,
         SYNOPSYS_UNCONNECTED_321, SYNOPSYS_UNCONNECTED_322,
         SYNOPSYS_UNCONNECTED_323, SYNOPSYS_UNCONNECTED_324,
         SYNOPSYS_UNCONNECTED_325, SYNOPSYS_UNCONNECTED_326,
         SYNOPSYS_UNCONNECTED_327, SYNOPSYS_UNCONNECTED_328,
         SYNOPSYS_UNCONNECTED_329, SYNOPSYS_UNCONNECTED_330,
         SYNOPSYS_UNCONNECTED_331, SYNOPSYS_UNCONNECTED_332,
         SYNOPSYS_UNCONNECTED_333, SYNOPSYS_UNCONNECTED_334,
         SYNOPSYS_UNCONNECTED_335, SYNOPSYS_UNCONNECTED_336,
         SYNOPSYS_UNCONNECTED_337, SYNOPSYS_UNCONNECTED_338,
         SYNOPSYS_UNCONNECTED_339, SYNOPSYS_UNCONNECTED_340,
         SYNOPSYS_UNCONNECTED_341, SYNOPSYS_UNCONNECTED_342,
         SYNOPSYS_UNCONNECTED_343, SYNOPSYS_UNCONNECTED_344,
         SYNOPSYS_UNCONNECTED_345, SYNOPSYS_UNCONNECTED_346,
         SYNOPSYS_UNCONNECTED_347, SYNOPSYS_UNCONNECTED_348,
         SYNOPSYS_UNCONNECTED_349, SYNOPSYS_UNCONNECTED_350,
         SYNOPSYS_UNCONNECTED_351, SYNOPSYS_UNCONNECTED_352,
         SYNOPSYS_UNCONNECTED_353, SYNOPSYS_UNCONNECTED_354,
         SYNOPSYS_UNCONNECTED_355, SYNOPSYS_UNCONNECTED_356,
         SYNOPSYS_UNCONNECTED_357, SYNOPSYS_UNCONNECTED_358,
         SYNOPSYS_UNCONNECTED_359, SYNOPSYS_UNCONNECTED_360,
         SYNOPSYS_UNCONNECTED_361, SYNOPSYS_UNCONNECTED_362,
         SYNOPSYS_UNCONNECTED_363, SYNOPSYS_UNCONNECTED_364,
         SYNOPSYS_UNCONNECTED_365, SYNOPSYS_UNCONNECTED_366,
         SYNOPSYS_UNCONNECTED_367, SYNOPSYS_UNCONNECTED_368,
         SYNOPSYS_UNCONNECTED_369, SYNOPSYS_UNCONNECTED_370,
         SYNOPSYS_UNCONNECTED_371, SYNOPSYS_UNCONNECTED_372,
         SYNOPSYS_UNCONNECTED_373, SYNOPSYS_UNCONNECTED_374,
         SYNOPSYS_UNCONNECTED_375, SYNOPSYS_UNCONNECTED_376,
         SYNOPSYS_UNCONNECTED_377, SYNOPSYS_UNCONNECTED_378,
         SYNOPSYS_UNCONNECTED_379, SYNOPSYS_UNCONNECTED_380,
         SYNOPSYS_UNCONNECTED_381, SYNOPSYS_UNCONNECTED_382,
         SYNOPSYS_UNCONNECTED_383, SYNOPSYS_UNCONNECTED_384,
         SYNOPSYS_UNCONNECTED_385, SYNOPSYS_UNCONNECTED_386,
         SYNOPSYS_UNCONNECTED_387, SYNOPSYS_UNCONNECTED_388,
         SYNOPSYS_UNCONNECTED_389, SYNOPSYS_UNCONNECTED_390,
         SYNOPSYS_UNCONNECTED_391, SYNOPSYS_UNCONNECTED_392,
         SYNOPSYS_UNCONNECTED_393, SYNOPSYS_UNCONNECTED_394,
         SYNOPSYS_UNCONNECTED_395, SYNOPSYS_UNCONNECTED_396,
         SYNOPSYS_UNCONNECTED_397, SYNOPSYS_UNCONNECTED_398,
         SYNOPSYS_UNCONNECTED_399, SYNOPSYS_UNCONNECTED_400,
         SYNOPSYS_UNCONNECTED_401, SYNOPSYS_UNCONNECTED_402,
         SYNOPSYS_UNCONNECTED_403, SYNOPSYS_UNCONNECTED_404,
         SYNOPSYS_UNCONNECTED_405, SYNOPSYS_UNCONNECTED_406,
         SYNOPSYS_UNCONNECTED_407, SYNOPSYS_UNCONNECTED_408,
         SYNOPSYS_UNCONNECTED_409, SYNOPSYS_UNCONNECTED_410,
         SYNOPSYS_UNCONNECTED_411, SYNOPSYS_UNCONNECTED_412;
  wire   [26:2] boothout1;
  wire   [26:0] boothout2;
  wire   [26:0] boothout3;
  wire   [26:0] boothout4;
  wire   [26:0] boothout5;
  wire   [26:0] boothout6;
  wire   [26:0] boothout7;
  wire   [26:0] boothout8;
  wire   [26:0] boothout9;
  wire   [26:0] boothout10;
  wire   [26:0] boothout11;
  wire   [25:0] boothout12;
  wire   [22:0] boothout13;
  wire   [29:2] cout1;
  wire   [31:3] mulout1;
  wire   [35:8] cout2;
  wire   [37:6] mulout2;
  wire   [41:14] cout3;
  wire   [42:12] mulout3;
  wire   [46:20] cout4;
  wire   [47:18] mulout4;
  wire   [31:3] cout5;
  wire   [46:4] mulout5;
  wire   [37:9] cout6;
  wire   [42:6] mulout6;
  wire   [46:18] cout7;
  wire   [47:12] mulout7;
  wire   [38:4] cout8;
  wire   [46:5] mulout8;
  wire   [46:12] cout9;
  wire   [47:6] mulout9;
  wire   [46:5] cout10;
  wire   [47:6] mulout10;
  wire   [46:6] cout11;
  wire   [47:7] mulout11;
  wire   [47:0] a;
  wire   [47:8] b;

  booth27_26 booth1 ( .out1({boothout1, SYNOPSYS_UNCONNECTED_1, 
        SYNOPSYS_UNCONNECTED_2}), .in1({in1[1:0], 1'b0}), .in2({1'b0, 1'b0, 
        1'b1, n33, n32, n31, n30, n29, n28, n27, n26, n25, n24, in2[12], n23, 
        in2[10], n22, in2[8], n20, in2[6], n19, in2[4], n18, in2[2], n17, 
        in2[0]}) );
  booth27_25 booth2 ( .out1(boothout2), .in1(in1[3:1]), .in2({1'b0, 1'b0, 1'b1, 
        n33, n32, n31, n30, n29, n28, n27, n26, n25, n24, in2[12], n23, 
        in2[10], n22, in2[8], n20, in2[6], n19, in2[4], n18, in2[2], n17, 
        in2[0]}) );
  booth27_24 booth3 ( .out1(boothout3), .in1(in1[5:3]), .in2({1'b0, 1'b0, 1'b1, 
        n33, n32, n31, n30, n29, n28, n27, n26, n25, n24, in2[12], n23, 
        in2[10], n22, in2[8], n20, in2[6], n19, in2[4], n18, in2[2], n17, 
        in2[0]}) );
  booth27_23 booth4 ( .out1(boothout4), .in1(in1[7:5]), .in2({1'b0, 1'b0, 1'b1, 
        n33, n32, n31, n30, n29, n28, n27, n26, n25, n24, in2[12], n23, 
        in2[10], n22, in2[8], n20, in2[6], n19, in2[4], n18, in2[2], n17, 
        in2[0]}) );
  booth27_22 booth5 ( .out1(boothout5), .in1(in1[9:7]), .in2({1'b0, 1'b0, 1'b1, 
        n33, n32, n31, n30, n29, n28, n27, n26, n25, n24, in2[12], n23, 
        in2[10], n22, in2[8], n20, in2[6], n19, in2[4], n18, in2[2], n17, 
        in2[0]}) );
  booth27_21 booth6 ( .out1(boothout6), .in1(in1[11:9]), .in2({1'b0, 1'b0, 
        1'b1, n33, n32, n31, n30, n29, n28, n27, n26, n25, n24, in2[12], n23, 
        in2[10], n22, in2[8], n20, in2[6], n19, in2[4], n18, in2[2], n17, 
        in2[0]}) );
  booth27_20 booth7 ( .out1(boothout7), .in1(in1[13:11]), .in2({1'b0, 1'b0, 
        1'b1, n33, n32, n31, n30, n29, n28, n27, n26, n25, n24, in2[12], n23, 
        in2[10], n22, in2[8], n20, in2[6], n19, in2[4], n18, in2[2], n17, 
        in2[0]}) );
  booth27_19 booth8 ( .out1(boothout8), .in1(in1[15:13]), .in2({1'b0, 1'b0, 
        1'b1, n33, n32, n31, n30, n29, n28, n27, n26, n25, n24, in2[12], n23, 
        in2[10], n22, in2[8], n20, in2[6], n19, in2[4], n18, in2[2], n17, 
        in2[0]}) );
  booth27_18 booth9 ( .out1(boothout9), .in1(in1[17:15]), .in2({1'b0, 1'b0, 
        1'b1, n33, n32, n31, n30, n29, n28, n27, n26, n25, n24, in2[12], n23, 
        in2[10], n22, in2[8], n20, in2[6], n19, in2[4], n18, in2[2], n17, 
        in2[0]}) );
  booth27_17 booth10 ( .out1(boothout10), .in1(in1[19:17]), .in2({1'b0, 1'b0, 
        1'b1, n33, n32, n31, n30, n29, n28, n27, n26, n25, n24, in2[12], n23, 
        in2[10], n22, in2[8], n20, in2[6], n19, in2[4], n18, in2[2], n17, 
        in2[0]}) );
  booth27_16 booth11 ( .out1(boothout11), .in1(in1[21:19]), .in2({1'b0, 1'b0, 
        1'b1, n33, n32, n31, n30, n29, n28, n27, n26, n25, n24, in2[12], n23, 
        in2[10], n22, in2[8], n20, in2[6], n19, in2[4], n18, in2[2], n17, 
        in2[0]}) );
  booth27_15 booth12 ( .out1({SYNOPSYS_UNCONNECTED_3, boothout12}), .in1({1'b1, 
        in1[22:21]}), .in2({1'b0, 1'b0, 1'b1, n33, n32, n31, n30, n29, n28, 
        n27, n26, n25, n24, in2[12], n23, in2[10], n22, in2[8], n20, in2[6], 
        n19, in2[4], n18, in2[2], n17, in2[0]}) );
  booth27_14 booth13 ( .out1({SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, 
        SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, boothout13}), .in1({
        1'b0, 1'b0, 1'b1}), .in2({1'b0, 1'b0, 1'b1, n33, n32, n31, n30, n29, 
        n28, n27, n26, n25, n24, in2[12], n23, in2[10], n22, in2[8], n20, 
        in2[6], n19, in2[4], n18, in2[2], n17, in2[0]}) );
  csa51squ_24 csa51squ1 ( .cout({SYNOPSYS_UNCONNECTED_8, 
        SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10, 
        SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12, 
        SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14, 
        SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16, 
        SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18, 
        SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20, 
        SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22, 
        SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24, 
        SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26, 
        SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28, cout1, 
        SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30}), .sumout({
        SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32, 
        SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34, 
        SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36, 
        SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38, 
        SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40, 
        SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42, 
        SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44, 
        SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46, 
        SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48, 
        SYNOPSYS_UNCONNECTED_49, mulout1[31], SYNOPSYS_UNCONNECTED_50, 
        mulout1[29:3], SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52, 
        SYNOPSYS_UNCONNECTED_53}), .in1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, boothout1, 1'b0, 1'b0}), .in2({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, boothout2, 
        1'b0, 1'b0}), .in3({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n131, 
        1'b0, boothout3[25:0], 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_23 csa51squ2 ( .cout({SYNOPSYS_UNCONNECTED_54, 
        SYNOPSYS_UNCONNECTED_55, SYNOPSYS_UNCONNECTED_56, 
        SYNOPSYS_UNCONNECTED_57, SYNOPSYS_UNCONNECTED_58, 
        SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_60, 
        SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_62, 
        SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_64, 
        SYNOPSYS_UNCONNECTED_65, SYNOPSYS_UNCONNECTED_66, 
        SYNOPSYS_UNCONNECTED_67, SYNOPSYS_UNCONNECTED_68, cout2, 
        SYNOPSYS_UNCONNECTED_69, SYNOPSYS_UNCONNECTED_70, 
        SYNOPSYS_UNCONNECTED_71, SYNOPSYS_UNCONNECTED_72, 
        SYNOPSYS_UNCONNECTED_73, SYNOPSYS_UNCONNECTED_74, 
        SYNOPSYS_UNCONNECTED_75, SYNOPSYS_UNCONNECTED_76}), .sumout({
        SYNOPSYS_UNCONNECTED_77, SYNOPSYS_UNCONNECTED_78, 
        SYNOPSYS_UNCONNECTED_79, SYNOPSYS_UNCONNECTED_80, 
        SYNOPSYS_UNCONNECTED_81, SYNOPSYS_UNCONNECTED_82, 
        SYNOPSYS_UNCONNECTED_83, SYNOPSYS_UNCONNECTED_84, 
        SYNOPSYS_UNCONNECTED_85, SYNOPSYS_UNCONNECTED_86, 
        SYNOPSYS_UNCONNECTED_87, SYNOPSYS_UNCONNECTED_88, 
        SYNOPSYS_UNCONNECTED_89, mulout2[37], SYNOPSYS_UNCONNECTED_90, 
        mulout2[35:6], SYNOPSYS_UNCONNECTED_91, SYNOPSYS_UNCONNECTED_92, 
        SYNOPSYS_UNCONNECTED_93, SYNOPSYS_UNCONNECTED_94, 
        SYNOPSYS_UNCONNECTED_95, SYNOPSYS_UNCONNECTED_96}), .in1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, boothout4, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, boothout5, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .in3({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n130, 1'b0, boothout6[25:0], 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_22 csa51squ3 ( .cout({SYNOPSYS_UNCONNECTED_97, 
        SYNOPSYS_UNCONNECTED_98, SYNOPSYS_UNCONNECTED_99, 
        SYNOPSYS_UNCONNECTED_100, SYNOPSYS_UNCONNECTED_101, 
        SYNOPSYS_UNCONNECTED_102, SYNOPSYS_UNCONNECTED_103, 
        SYNOPSYS_UNCONNECTED_104, SYNOPSYS_UNCONNECTED_105, cout3, 
        SYNOPSYS_UNCONNECTED_106, SYNOPSYS_UNCONNECTED_107, 
        SYNOPSYS_UNCONNECTED_108, SYNOPSYS_UNCONNECTED_109, 
        SYNOPSYS_UNCONNECTED_110, SYNOPSYS_UNCONNECTED_111, 
        SYNOPSYS_UNCONNECTED_112, SYNOPSYS_UNCONNECTED_113, 
        SYNOPSYS_UNCONNECTED_114, SYNOPSYS_UNCONNECTED_115, 
        SYNOPSYS_UNCONNECTED_116, SYNOPSYS_UNCONNECTED_117, 
        SYNOPSYS_UNCONNECTED_118, SYNOPSYS_UNCONNECTED_119}), .sumout({
        SYNOPSYS_UNCONNECTED_120, SYNOPSYS_UNCONNECTED_121, 
        SYNOPSYS_UNCONNECTED_122, SYNOPSYS_UNCONNECTED_123, 
        SYNOPSYS_UNCONNECTED_124, SYNOPSYS_UNCONNECTED_125, 
        SYNOPSYS_UNCONNECTED_126, SYNOPSYS_UNCONNECTED_127, mulout3, 
        SYNOPSYS_UNCONNECTED_128, SYNOPSYS_UNCONNECTED_129, 
        SYNOPSYS_UNCONNECTED_130, SYNOPSYS_UNCONNECTED_131, 
        SYNOPSYS_UNCONNECTED_132, SYNOPSYS_UNCONNECTED_133, 
        SYNOPSYS_UNCONNECTED_134, SYNOPSYS_UNCONNECTED_135, 
        SYNOPSYS_UNCONNECTED_136, SYNOPSYS_UNCONNECTED_137, 
        SYNOPSYS_UNCONNECTED_138, SYNOPSYS_UNCONNECTED_139}), .in1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, boothout7, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, boothout8, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .in3({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        boothout9, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_21 csa51squ4 ( .cout({SYNOPSYS_UNCONNECTED_140, 
        SYNOPSYS_UNCONNECTED_141, SYNOPSYS_UNCONNECTED_142, 
        SYNOPSYS_UNCONNECTED_143, cout4, SYNOPSYS_UNCONNECTED_144, 
        SYNOPSYS_UNCONNECTED_145, SYNOPSYS_UNCONNECTED_146, 
        SYNOPSYS_UNCONNECTED_147, SYNOPSYS_UNCONNECTED_148, 
        SYNOPSYS_UNCONNECTED_149, SYNOPSYS_UNCONNECTED_150, 
        SYNOPSYS_UNCONNECTED_151, SYNOPSYS_UNCONNECTED_152, 
        SYNOPSYS_UNCONNECTED_153, SYNOPSYS_UNCONNECTED_154, 
        SYNOPSYS_UNCONNECTED_155, SYNOPSYS_UNCONNECTED_156, 
        SYNOPSYS_UNCONNECTED_157, SYNOPSYS_UNCONNECTED_158, 
        SYNOPSYS_UNCONNECTED_159, SYNOPSYS_UNCONNECTED_160, 
        SYNOPSYS_UNCONNECTED_161, SYNOPSYS_UNCONNECTED_162, 
        SYNOPSYS_UNCONNECTED_163}), .sumout({SYNOPSYS_UNCONNECTED_164, 
        SYNOPSYS_UNCONNECTED_165, SYNOPSYS_UNCONNECTED_166, mulout4, 
        SYNOPSYS_UNCONNECTED_167, SYNOPSYS_UNCONNECTED_168, 
        SYNOPSYS_UNCONNECTED_169, SYNOPSYS_UNCONNECTED_170, 
        SYNOPSYS_UNCONNECTED_171, SYNOPSYS_UNCONNECTED_172, 
        SYNOPSYS_UNCONNECTED_173, SYNOPSYS_UNCONNECTED_174, 
        SYNOPSYS_UNCONNECTED_175, SYNOPSYS_UNCONNECTED_176, 
        SYNOPSYS_UNCONNECTED_177, SYNOPSYS_UNCONNECTED_178, 
        SYNOPSYS_UNCONNECTED_179, SYNOPSYS_UNCONNECTED_180, 
        SYNOPSYS_UNCONNECTED_181, SYNOPSYS_UNCONNECTED_182, 
        SYNOPSYS_UNCONNECTED_183, SYNOPSYS_UNCONNECTED_184}), .in1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, boothout10, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 1'b0, 1'b0, 1'b0, boothout11, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .in3({1'b0, 1'b0, 1'b0, boothout12, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_20 csa51squ5 ( .cout({SYNOPSYS_UNCONNECTED_185, 
        SYNOPSYS_UNCONNECTED_186, SYNOPSYS_UNCONNECTED_187, 
        SYNOPSYS_UNCONNECTED_188, SYNOPSYS_UNCONNECTED_189, 
        SYNOPSYS_UNCONNECTED_190, SYNOPSYS_UNCONNECTED_191, 
        SYNOPSYS_UNCONNECTED_192, SYNOPSYS_UNCONNECTED_193, 
        SYNOPSYS_UNCONNECTED_194, SYNOPSYS_UNCONNECTED_195, 
        SYNOPSYS_UNCONNECTED_196, SYNOPSYS_UNCONNECTED_197, 
        SYNOPSYS_UNCONNECTED_198, SYNOPSYS_UNCONNECTED_199, 
        SYNOPSYS_UNCONNECTED_200, SYNOPSYS_UNCONNECTED_201, 
        SYNOPSYS_UNCONNECTED_202, SYNOPSYS_UNCONNECTED_203, cout5, 
        SYNOPSYS_UNCONNECTED_204, SYNOPSYS_UNCONNECTED_205, 
        SYNOPSYS_UNCONNECTED_206}), .sumout({SYNOPSYS_UNCONNECTED_207, 
        SYNOPSYS_UNCONNECTED_208, SYNOPSYS_UNCONNECTED_209, 
        SYNOPSYS_UNCONNECTED_210, mulout5, SYNOPSYS_UNCONNECTED_211, 
        SYNOPSYS_UNCONNECTED_212, SYNOPSYS_UNCONNECTED_213, 
        SYNOPSYS_UNCONNECTED_214}), .in1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, cout1, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, mulout1[31], 1'b0, mulout1[29:3], 1'b0, 1'b0, 1'b0}), 
        .in3({1'b0, 1'b0, 1'b0, 1'b1, boothout13, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_19 csa51squ6 ( .cout({SYNOPSYS_UNCONNECTED_215, 
        SYNOPSYS_UNCONNECTED_216, SYNOPSYS_UNCONNECTED_217, 
        SYNOPSYS_UNCONNECTED_218, SYNOPSYS_UNCONNECTED_219, 
        SYNOPSYS_UNCONNECTED_220, SYNOPSYS_UNCONNECTED_221, 
        SYNOPSYS_UNCONNECTED_222, SYNOPSYS_UNCONNECTED_223, 
        SYNOPSYS_UNCONNECTED_224, SYNOPSYS_UNCONNECTED_225, 
        SYNOPSYS_UNCONNECTED_226, SYNOPSYS_UNCONNECTED_227, cout6, 
        SYNOPSYS_UNCONNECTED_228, SYNOPSYS_UNCONNECTED_229, 
        SYNOPSYS_UNCONNECTED_230, SYNOPSYS_UNCONNECTED_231, 
        SYNOPSYS_UNCONNECTED_232, SYNOPSYS_UNCONNECTED_233, 
        SYNOPSYS_UNCONNECTED_234, SYNOPSYS_UNCONNECTED_235, 
        SYNOPSYS_UNCONNECTED_236}), .sumout({SYNOPSYS_UNCONNECTED_237, 
        SYNOPSYS_UNCONNECTED_238, SYNOPSYS_UNCONNECTED_239, 
        SYNOPSYS_UNCONNECTED_240, SYNOPSYS_UNCONNECTED_241, 
        SYNOPSYS_UNCONNECTED_242, SYNOPSYS_UNCONNECTED_243, 
        SYNOPSYS_UNCONNECTED_244, mulout6, SYNOPSYS_UNCONNECTED_245, 
        SYNOPSYS_UNCONNECTED_246, SYNOPSYS_UNCONNECTED_247, 
        SYNOPSYS_UNCONNECTED_248, SYNOPSYS_UNCONNECTED_249, 
        SYNOPSYS_UNCONNECTED_250}), .in1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, cout2, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        mulout2[37], 1'b0, mulout2[35:6], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .in3({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, cout3, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  csa51squ_18 csa51squ7 ( .cout({SYNOPSYS_UNCONNECTED_251, 
        SYNOPSYS_UNCONNECTED_252, SYNOPSYS_UNCONNECTED_253, 
        SYNOPSYS_UNCONNECTED_254, cout7, SYNOPSYS_UNCONNECTED_255, 
        SYNOPSYS_UNCONNECTED_256, SYNOPSYS_UNCONNECTED_257, 
        SYNOPSYS_UNCONNECTED_258, SYNOPSYS_UNCONNECTED_259, 
        SYNOPSYS_UNCONNECTED_260, SYNOPSYS_UNCONNECTED_261, 
        SYNOPSYS_UNCONNECTED_262, SYNOPSYS_UNCONNECTED_263, 
        SYNOPSYS_UNCONNECTED_264, SYNOPSYS_UNCONNECTED_265, 
        SYNOPSYS_UNCONNECTED_266, SYNOPSYS_UNCONNECTED_267, 
        SYNOPSYS_UNCONNECTED_268, SYNOPSYS_UNCONNECTED_269, 
        SYNOPSYS_UNCONNECTED_270, SYNOPSYS_UNCONNECTED_271, 
        SYNOPSYS_UNCONNECTED_272}), .sumout({SYNOPSYS_UNCONNECTED_273, 
        SYNOPSYS_UNCONNECTED_274, SYNOPSYS_UNCONNECTED_275, mulout7, 
        SYNOPSYS_UNCONNECTED_276, SYNOPSYS_UNCONNECTED_277, 
        SYNOPSYS_UNCONNECTED_278, SYNOPSYS_UNCONNECTED_279, 
        SYNOPSYS_UNCONNECTED_280, SYNOPSYS_UNCONNECTED_281, 
        SYNOPSYS_UNCONNECTED_282, SYNOPSYS_UNCONNECTED_283, 
        SYNOPSYS_UNCONNECTED_284, SYNOPSYS_UNCONNECTED_285, 
        SYNOPSYS_UNCONNECTED_286, SYNOPSYS_UNCONNECTED_287}), .in1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mulout3, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 1'b0, 
        1'b0, cout4, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in3({1'b0, 1'b0, 1'b0, mulout4, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_17 csa51squ8 ( .cout({SYNOPSYS_UNCONNECTED_288, 
        SYNOPSYS_UNCONNECTED_289, SYNOPSYS_UNCONNECTED_290, 
        SYNOPSYS_UNCONNECTED_291, SYNOPSYS_UNCONNECTED_292, 
        SYNOPSYS_UNCONNECTED_293, SYNOPSYS_UNCONNECTED_294, 
        SYNOPSYS_UNCONNECTED_295, SYNOPSYS_UNCONNECTED_296, 
        SYNOPSYS_UNCONNECTED_297, SYNOPSYS_UNCONNECTED_298, 
        SYNOPSYS_UNCONNECTED_299, cout8, SYNOPSYS_UNCONNECTED_300, 
        SYNOPSYS_UNCONNECTED_301, SYNOPSYS_UNCONNECTED_302, 
        SYNOPSYS_UNCONNECTED_303}), .sumout({SYNOPSYS_UNCONNECTED_304, 
        SYNOPSYS_UNCONNECTED_305, SYNOPSYS_UNCONNECTED_306, 
        SYNOPSYS_UNCONNECTED_307, mulout8, SYNOPSYS_UNCONNECTED_308, 
        SYNOPSYS_UNCONNECTED_309, SYNOPSYS_UNCONNECTED_310, 
        SYNOPSYS_UNCONNECTED_311, SYNOPSYS_UNCONNECTED_312}), .in1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, cout5, 1'b0, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 
        1'b0, 1'b0, 1'b1, mulout5, 1'b0, 1'b0, 1'b0, 1'b0}), .in3({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, cout6, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_16 csa51squ9 ( .cout({SYNOPSYS_UNCONNECTED_313, 
        SYNOPSYS_UNCONNECTED_314, SYNOPSYS_UNCONNECTED_315, 
        SYNOPSYS_UNCONNECTED_316, cout9, SYNOPSYS_UNCONNECTED_317, 
        SYNOPSYS_UNCONNECTED_318, SYNOPSYS_UNCONNECTED_319, 
        SYNOPSYS_UNCONNECTED_320, SYNOPSYS_UNCONNECTED_321, 
        SYNOPSYS_UNCONNECTED_322, SYNOPSYS_UNCONNECTED_323, 
        SYNOPSYS_UNCONNECTED_324, SYNOPSYS_UNCONNECTED_325, 
        SYNOPSYS_UNCONNECTED_326, SYNOPSYS_UNCONNECTED_327, 
        SYNOPSYS_UNCONNECTED_328}), .sumout({SYNOPSYS_UNCONNECTED_329, 
        SYNOPSYS_UNCONNECTED_330, SYNOPSYS_UNCONNECTED_331, mulout9, 
        SYNOPSYS_UNCONNECTED_332, SYNOPSYS_UNCONNECTED_333, 
        SYNOPSYS_UNCONNECTED_334, SYNOPSYS_UNCONNECTED_335, 
        SYNOPSYS_UNCONNECTED_336, SYNOPSYS_UNCONNECTED_337}), .in1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mulout6, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .in2({1'b0, 1'b0, 1'b0, cout7, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .in3({1'b0, 1'b0, 1'b0, mulout7, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_15 csa51squ10 ( .cout({SYNOPSYS_UNCONNECTED_338, 
        SYNOPSYS_UNCONNECTED_339, SYNOPSYS_UNCONNECTED_340, 
        SYNOPSYS_UNCONNECTED_341, cout10, SYNOPSYS_UNCONNECTED_342, 
        SYNOPSYS_UNCONNECTED_343, SYNOPSYS_UNCONNECTED_344, 
        SYNOPSYS_UNCONNECTED_345, SYNOPSYS_UNCONNECTED_346}), .sumout({
        SYNOPSYS_UNCONNECTED_347, SYNOPSYS_UNCONNECTED_348, 
        SYNOPSYS_UNCONNECTED_349, mulout10, SYNOPSYS_UNCONNECTED_350, 
        SYNOPSYS_UNCONNECTED_351, SYNOPSYS_UNCONNECTED_352, 
        SYNOPSYS_UNCONNECTED_353, SYNOPSYS_UNCONNECTED_354, 
        SYNOPSYS_UNCONNECTED_355}), .in1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, cout8, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .in2({1'b0, 1'b0, 1'b0, 1'b1, mulout8, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .in3({1'b0, 1'b0, 1'b0, cout9, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_14 csa51squ11 ( .cout({SYNOPSYS_UNCONNECTED_356, 
        SYNOPSYS_UNCONNECTED_357, SYNOPSYS_UNCONNECTED_358, 
        SYNOPSYS_UNCONNECTED_359, cout11, SYNOPSYS_UNCONNECTED_360, 
        SYNOPSYS_UNCONNECTED_361, SYNOPSYS_UNCONNECTED_362, 
        SYNOPSYS_UNCONNECTED_363, SYNOPSYS_UNCONNECTED_364, 
        SYNOPSYS_UNCONNECTED_365}), .sumout({SYNOPSYS_UNCONNECTED_366, 
        SYNOPSYS_UNCONNECTED_367, SYNOPSYS_UNCONNECTED_368, mulout11, 
        SYNOPSYS_UNCONNECTED_369, SYNOPSYS_UNCONNECTED_370, 
        SYNOPSYS_UNCONNECTED_371, SYNOPSYS_UNCONNECTED_372, 
        SYNOPSYS_UNCONNECTED_373, SYNOPSYS_UNCONNECTED_374, 
        SYNOPSYS_UNCONNECTED_375}), .in1({1'b0, 1'b0, 1'b0, mulout9, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 1'b0, 1'b0, cout10, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in3({1'b0, 1'b0, 1'b0, mulout10, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_13 csa51squ12 ( .sumout({SYNOPSYS_UNCONNECTED_376, 
        SYNOPSYS_UNCONNECTED_377, SYNOPSYS_UNCONNECTED_378, N101, N100, N99, 
        N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, 
        N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, 
        N70, N69, N68, N67, N66, N65, N64, N63, N62, SYNOPSYS_UNCONNECTED_379, 
        SYNOPSYS_UNCONNECTED_380, SYNOPSYS_UNCONNECTED_381, 
        SYNOPSYS_UNCONNECTED_382, SYNOPSYS_UNCONNECTED_383, 
        SYNOPSYS_UNCONNECTED_384, SYNOPSYS_UNCONNECTED_385, 
        SYNOPSYS_UNCONNECTED_386}), .in1({1'b0, 1'b0, 1'b0, mulout11, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 1'b0, 1'b0, cout11, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in3({1'b1, 1'b0, 1'b1, 
        1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 
        1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .cout_46_(N50), .cout_44_(N48), .cout_42_(N46), .cout_40_(N44), .cout_38_(
        N42), .cout_36_(N40), .cout_34_(N38), .cout_32_(N36), .cout_30_(N34), 
        .cout_28_(N32), .cout_27_(N31), .cout_7__BAR(N11), .cout_8__BAR(N12), 
        .cout_9__BAR(N13), .cout_10__BAR(N14), .cout_11__BAR(N15), 
        .cout_12__BAR(N16), .cout_13__BAR(N17), .cout_14__BAR(N18), 
        .cout_15__BAR(N19), .cout_16__BAR(N20), .cout_17__BAR(N21), 
        .cout_18__BAR(N22), .cout_19__BAR(N23), .cout_20__BAR(N24), 
        .cout_21__BAR(N25), .cout_22__BAR(N26), .cout_23__BAR(N27), 
        .cout_24__BAR(N28), .cout_25__BAR(N29), .cout_26__BAR(N30), 
        .cout_29__BAR(N33), .cout_31__BAR(N35), .cout_33__BAR(N37), 
        .cout_35__BAR(N39), .cout_37__BAR(N41), .cout_39__BAR(N43), 
        .cout_41__BAR(N45), .cout_43__BAR(N47), .cout_45__BAR(N49) );
  cla51squ_2 cla51squ ( .out({SYNOPSYS_UNCONNECTED_387, 
        SYNOPSYS_UNCONNECTED_388, SYNOPSYS_UNCONNECTED_389, mulout[47:23], 
        SYNOPSYS_UNCONNECTED_390, SYNOPSYS_UNCONNECTED_391, 
        SYNOPSYS_UNCONNECTED_392, SYNOPSYS_UNCONNECTED_393, 
        SYNOPSYS_UNCONNECTED_394, SYNOPSYS_UNCONNECTED_395, 
        SYNOPSYS_UNCONNECTED_396, SYNOPSYS_UNCONNECTED_397, 
        SYNOPSYS_UNCONNECTED_398, SYNOPSYS_UNCONNECTED_399, 
        SYNOPSYS_UNCONNECTED_400, SYNOPSYS_UNCONNECTED_401, 
        SYNOPSYS_UNCONNECTED_402, SYNOPSYS_UNCONNECTED_403, 
        SYNOPSYS_UNCONNECTED_404, SYNOPSYS_UNCONNECTED_405, 
        SYNOPSYS_UNCONNECTED_406, SYNOPSYS_UNCONNECTED_407, 
        SYNOPSYS_UNCONNECTED_408, SYNOPSYS_UNCONNECTED_409, 
        SYNOPSYS_UNCONNECTED_410, SYNOPSYS_UNCONNECTED_411, 
        SYNOPSYS_UNCONNECTED_412}), .a({1'b0, 1'b0, 1'b0, a[47:8], 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({1'b0, 1'b0, 1'b0, b, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  DFFARX1 b_reg_47_ ( .D(N101), .CLK(clk), .RSTB(rst_n), .Q(b[47]) );
  DFFARX1 b_reg_46_ ( .D(N100), .CLK(clk), .RSTB(rst_n), .Q(b[46]) );
  DFFARX1 b_reg_45_ ( .D(N99), .CLK(clk), .RSTB(rst_n), .Q(b[45]) );
  DFFARX1 b_reg_44_ ( .D(N98), .CLK(clk), .RSTB(rst_n), .Q(b[44]) );
  DFFARX1 b_reg_43_ ( .D(N97), .CLK(clk), .RSTB(rst_n), .Q(b[43]) );
  DFFARX1 b_reg_42_ ( .D(N96), .CLK(clk), .RSTB(rst_n), .Q(b[42]) );
  DFFARX1 b_reg_41_ ( .D(N95), .CLK(clk), .RSTB(rst_n), .Q(b[41]) );
  DFFARX1 b_reg_40_ ( .D(N94), .CLK(clk), .RSTB(rst_n), .Q(b[40]) );
  DFFARX1 b_reg_39_ ( .D(N93), .CLK(clk), .RSTB(rst_n), .Q(b[39]) );
  DFFARX1 b_reg_38_ ( .D(N92), .CLK(clk), .RSTB(rst_n), .Q(b[38]) );
  DFFARX1 b_reg_37_ ( .D(N91), .CLK(clk), .RSTB(rst_n), .Q(b[37]) );
  DFFARX1 b_reg_36_ ( .D(N90), .CLK(clk), .RSTB(rst_n), .Q(b[36]) );
  DFFARX1 b_reg_35_ ( .D(N89), .CLK(clk), .RSTB(rst_n), .Q(b[35]) );
  DFFARX1 b_reg_34_ ( .D(N88), .CLK(clk), .RSTB(rst_n), .Q(b[34]) );
  DFFARX1 b_reg_33_ ( .D(N87), .CLK(clk), .RSTB(rst_n), .Q(b[33]) );
  DFFARX1 b_reg_32_ ( .D(N86), .CLK(clk), .RSTB(rst_n), .Q(b[32]) );
  DFFARX1 b_reg_31_ ( .D(N85), .CLK(clk), .RSTB(rst_n), .Q(b[31]) );
  DFFARX1 b_reg_30_ ( .D(N84), .CLK(clk), .RSTB(rst_n), .Q(b[30]) );
  DFFARX1 b_reg_29_ ( .D(N83), .CLK(clk), .RSTB(rst_n), .Q(b[29]) );
  DFFARX1 b_reg_28_ ( .D(N82), .CLK(clk), .RSTB(rst_n), .Q(b[28]) );
  DFFARX1 b_reg_27_ ( .D(N81), .CLK(clk), .RSTB(rst_n), .Q(b[27]) );
  DFFARX1 b_reg_26_ ( .D(N80), .CLK(clk), .RSTB(rst_n), .Q(b[26]) );
  DFFARX1 b_reg_25_ ( .D(N79), .CLK(clk), .RSTB(rst_n), .Q(b[25]) );
  DFFARX1 b_reg_24_ ( .D(N78), .CLK(clk), .RSTB(rst_n), .Q(b[24]) );
  DFFARX1 b_reg_23_ ( .D(N77), .CLK(clk), .RSTB(rst_n), .Q(b[23]) );
  DFFARX1 b_reg_22_ ( .D(N76), .CLK(clk), .RSTB(rst_n), .Q(b[22]) );
  DFFARX1 b_reg_21_ ( .D(N75), .CLK(clk), .RSTB(rst_n), .Q(b[21]) );
  DFFARX1 b_reg_20_ ( .D(N74), .CLK(clk), .RSTB(rst_n), .Q(b[20]) );
  DFFARX1 b_reg_19_ ( .D(N73), .CLK(clk), .RSTB(rst_n), .Q(b[19]) );
  DFFARX1 b_reg_18_ ( .D(N72), .CLK(clk), .RSTB(rst_n), .Q(b[18]) );
  DFFARX1 b_reg_17_ ( .D(N71), .CLK(clk), .RSTB(rst_n), .Q(b[17]) );
  DFFARX1 b_reg_16_ ( .D(N70), .CLK(clk), .RSTB(rst_n), .Q(b[16]) );
  DFFARX1 b_reg_15_ ( .D(N69), .CLK(clk), .RSTB(rst_n), .Q(b[15]) );
  DFFARX1 b_reg_14_ ( .D(N68), .CLK(clk), .RSTB(rst_n), .Q(b[14]) );
  DFFARX1 b_reg_13_ ( .D(N67), .CLK(clk), .RSTB(rst_n), .Q(b[13]) );
  DFFARX1 b_reg_12_ ( .D(N66), .CLK(clk), .RSTB(rst_n), .Q(b[12]) );
  DFFARX1 b_reg_11_ ( .D(N65), .CLK(clk), .RSTB(rst_n), .Q(b[11]) );
  DFFARX1 b_reg_10_ ( .D(N64), .CLK(clk), .RSTB(rst_n), .Q(b[10]) );
  DFFARX1 b_reg_9_ ( .D(N63), .CLK(clk), .RSTB(rst_n), .Q(b[9]) );
  DFFARX1 b_reg_8_ ( .D(N62), .CLK(clk), .RSTB(rst_n), .Q(b[8]) );
  DFFARX1 a_reg_47_ ( .D(N50), .CLK(clk), .RSTB(rst_n), .Q(a[47]) );
  DFFARX1 a_reg_46_ ( .D(n62), .CLK(clk), .RSTB(rst_n), .Q(a[46]) );
  DFFARX1 a_reg_45_ ( .D(N48), .CLK(clk), .RSTB(rst_n), .Q(a[45]) );
  DFFARX1 a_reg_44_ ( .D(n63), .CLK(clk), .RSTB(rst_n), .Q(a[44]) );
  DFFARX1 a_reg_43_ ( .D(N46), .CLK(clk), .RSTB(rst_n), .Q(a[43]) );
  DFFARX1 a_reg_42_ ( .D(n64), .CLK(clk), .RSTB(rst_n), .Q(a[42]) );
  DFFARX1 a_reg_41_ ( .D(N44), .CLK(clk), .RSTB(rst_n), .Q(a[41]) );
  DFFARX1 a_reg_40_ ( .D(n65), .CLK(clk), .RSTB(rst_n), .Q(a[40]) );
  DFFARX1 a_reg_39_ ( .D(N42), .CLK(clk), .RSTB(rst_n), .Q(a[39]) );
  DFFARX1 a_reg_38_ ( .D(n66), .CLK(clk), .RSTB(rst_n), .Q(a[38]) );
  DFFARX1 a_reg_37_ ( .D(N40), .CLK(clk), .RSTB(rst_n), .Q(a[37]) );
  DFFARX1 a_reg_36_ ( .D(n67), .CLK(clk), .RSTB(rst_n), .Q(a[36]) );
  DFFARX1 a_reg_35_ ( .D(N38), .CLK(clk), .RSTB(rst_n), .Q(a[35]) );
  DFFARX1 a_reg_34_ ( .D(n68), .CLK(clk), .RSTB(rst_n), .Q(a[34]) );
  DFFARX1 a_reg_33_ ( .D(N36), .CLK(clk), .RSTB(rst_n), .Q(a[33]) );
  DFFARX1 a_reg_32_ ( .D(n69), .CLK(clk), .RSTB(rst_n), .Q(a[32]) );
  DFFARX1 a_reg_31_ ( .D(N34), .CLK(clk), .RSTB(rst_n), .Q(a[31]) );
  DFFARX1 a_reg_30_ ( .D(n70), .CLK(clk), .RSTB(rst_n), .Q(a[30]) );
  DFFARX1 a_reg_29_ ( .D(N32), .CLK(clk), .RSTB(rst_n), .Q(a[29]) );
  DFFARX1 a_reg_28_ ( .D(N31), .CLK(clk), .RSTB(rst_n), .Q(a[28]) );
  DFFARX1 a_reg_27_ ( .D(n71), .CLK(clk), .RSTB(rst_n), .Q(a[27]) );
  DFFARX1 a_reg_26_ ( .D(n72), .CLK(clk), .RSTB(rst_n), .Q(a[26]) );
  DFFARX1 a_reg_25_ ( .D(n73), .CLK(clk), .RSTB(rst_n), .Q(a[25]) );
  DFFARX1 a_reg_24_ ( .D(n74), .CLK(clk), .RSTB(rst_n), .Q(a[24]) );
  DFFARX1 a_reg_23_ ( .D(n75), .CLK(clk), .RSTB(rst_n), .Q(a[23]) );
  DFFARX1 a_reg_22_ ( .D(n76), .CLK(clk), .RSTB(rst_n), .Q(a[22]) );
  DFFARX1 a_reg_21_ ( .D(n77), .CLK(clk), .RSTB(rst_n), .Q(a[21]) );
  DFFARX1 a_reg_20_ ( .D(n78), .CLK(clk), .RSTB(rst_n), .Q(a[20]) );
  DFFARX1 a_reg_19_ ( .D(n79), .CLK(clk), .RSTB(rst_n), .Q(a[19]) );
  DFFARX1 a_reg_18_ ( .D(n80), .CLK(clk), .RSTB(rst_n), .Q(a[18]) );
  DFFARX1 a_reg_17_ ( .D(n81), .CLK(clk), .RSTB(rst_n), .Q(a[17]) );
  DFFARX1 a_reg_16_ ( .D(n82), .CLK(clk), .RSTB(rst_n), .Q(a[16]) );
  DFFARX1 a_reg_15_ ( .D(n83), .CLK(clk), .RSTB(rst_n), .Q(a[15]) );
  DFFARX1 a_reg_14_ ( .D(n84), .CLK(clk), .RSTB(rst_n), .Q(a[14]) );
  DFFARX1 a_reg_13_ ( .D(n85), .CLK(clk), .RSTB(rst_n), .Q(a[13]) );
  DFFARX1 a_reg_12_ ( .D(n86), .CLK(clk), .RSTB(rst_n), .Q(a[12]) );
  DFFARX1 a_reg_11_ ( .D(n87), .CLK(clk), .RSTB(rst_n), .Q(a[11]) );
  DFFARX1 a_reg_10_ ( .D(n88), .CLK(clk), .RSTB(rst_n), .Q(a[10]) );
  DFFARX1 a_reg_9_ ( .D(n89), .CLK(clk), .RSTB(rst_n), .Q(a[9]) );
  DFFARX1 a_reg_8_ ( .D(n90), .CLK(clk), .RSTB(rst_n), .Q(a[8]) );
  INVX0 U5 ( .INP(boothout3[26]), .ZN(n131) );
  INVX0 U8 ( .INP(boothout6[26]), .ZN(n130) );
  NBUFFX8 U3 ( .INP(in2[18]), .Z(n29) );
  NBUFFX8 U4 ( .INP(in2[16]), .Z(n27) );
  NBUFFX8 U6 ( .INP(in2[14]), .Z(n25) );
  NBUFFX8 U7 ( .INP(in2[20]), .Z(n31) );
  NBUFFX8 U9 ( .INP(in2[19]), .Z(n30) );
  NBUFFX8 U10 ( .INP(in2[15]), .Z(n26) );
  NBUFFX8 U11 ( .INP(in2[17]), .Z(n28) );
  NBUFFX8 U12 ( .INP(in2[13]), .Z(n24) );
  NBUFFX8 U13 ( .INP(in2[21]), .Z(n32) );
  NBUFFX8 U14 ( .INP(in2[22]), .Z(n33) );
  NBUFFX8 U15 ( .INP(in2[3]), .Z(n18) );
  NBUFFX8 U16 ( .INP(in2[9]), .Z(n22) );
  NBUFFX8 U17 ( .INP(in2[11]), .Z(n23) );
  NBUFFX8 U18 ( .INP(in2[5]), .Z(n19) );
  INVX0 U19 ( .INP(n21), .ZN(n20) );
  NBUFFX8 U20 ( .INP(in2[1]), .Z(n17) );
  INVX0 U35 ( .INP(in2[7]), .ZN(n21) );
  INVX0 U71 ( .INP(N49), .ZN(n62) );
  INVX0 U72 ( .INP(N47), .ZN(n63) );
  INVX0 U73 ( .INP(N45), .ZN(n64) );
  INVX0 U74 ( .INP(N43), .ZN(n65) );
  INVX0 U75 ( .INP(N41), .ZN(n66) );
  INVX0 U76 ( .INP(N39), .ZN(n67) );
  INVX0 U77 ( .INP(N37), .ZN(n68) );
  INVX0 U78 ( .INP(N35), .ZN(n69) );
  INVX0 U79 ( .INP(N33), .ZN(n70) );
  INVX0 U80 ( .INP(N30), .ZN(n71) );
  INVX0 U81 ( .INP(N29), .ZN(n72) );
  INVX0 U82 ( .INP(N28), .ZN(n73) );
  INVX0 U83 ( .INP(N27), .ZN(n74) );
  INVX0 U84 ( .INP(N26), .ZN(n75) );
  INVX0 U85 ( .INP(N25), .ZN(n76) );
  INVX0 U86 ( .INP(N24), .ZN(n77) );
  INVX0 U87 ( .INP(N23), .ZN(n78) );
  INVX0 U88 ( .INP(N22), .ZN(n79) );
  INVX0 U89 ( .INP(N21), .ZN(n80) );
  INVX0 U90 ( .INP(N20), .ZN(n81) );
  INVX0 U91 ( .INP(N19), .ZN(n82) );
  INVX0 U92 ( .INP(N18), .ZN(n83) );
  INVX0 U93 ( .INP(N17), .ZN(n84) );
  INVX0 U94 ( .INP(N16), .ZN(n85) );
  INVX0 U95 ( .INP(N15), .ZN(n86) );
  INVX0 U96 ( .INP(N14), .ZN(n87) );
  INVX0 U97 ( .INP(N13), .ZN(n88) );
  INVX0 U98 ( .INP(N12), .ZN(n89) );
  INVX0 U99 ( .INP(N11), .ZN(n90) );
endmodule


module add_209 ( s, a, b, co, ci_BAR );
  input a, b, ci_BAR;
  output s, co;


  XOR2X1 U1 ( .IN1(a), .IN2(ci_BAR), .Q(s) );
endmodule


module add_210 ( s, a, b, ci, co_BAR );
  input a, b, ci;
  output s, co_BAR;


  NAND2X0 U1 ( .IN1(ci), .IN2(a), .QN(co_BAR) );
  OA21X1 U2 ( .IN1(ci), .IN2(a), .IN3(co_BAR), .Q(s) );
endmodule


module add_211 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_212 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_213 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_214 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_215 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  INVX0 U1 ( .INP(a), .ZN(s) );
  NBUFFX2 U2 ( .INP(a), .Z(co) );
endmodule


module add_216 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  NBUFFX2 U1 ( .INP(a), .Z(s) );
endmodule


module adder8_15 ( out, a, b, cin );
  output [7:0] out;
  input [7:0] a;
  input [7:0] b;
  input cin;

  wire   [6:1] c;

  add_216 add_01 ( .s(out[0]), .a(a[0]), .b(1'b1), .ci(1'b1) );
  add_215 add_02 ( .s(out[1]), .a(a[1]), .b(1'b0), .ci(1'b1), .co(c[1]) );
  add_214 add_03 ( .s(out[2]), .a(a[2]), .b(1'b0), .ci(c[1]), .co(c[2]) );
  add_213 add_04 ( .s(out[3]), .a(a[3]), .b(1'b0), .ci(c[2]), .co(c[3]) );
  add_212 add_05 ( .s(out[4]), .a(a[4]), .b(1'b0), .ci(c[3]), .co(c[4]) );
  add_211 add_06 ( .s(out[5]), .a(a[5]), .b(1'b0), .ci(c[4]), .co(c[5]) );
  add_210 add_07 ( .s(out[6]), .a(a[6]), .b(1'b0), .ci(c[5]), .co_BAR(c[6]) );
  add_209 add_08 ( .s(out[7]), .a(a[7]), .b(1'b1), .ci_BAR(c[6]) );
endmodule


module add_217 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  XOR3X1 U1 ( .IN1(b), .IN2(ci), .IN3(a), .Q(s) );
endmodule


module add_218 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_219 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_220 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_221 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_222 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_223 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_224 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(b), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(b), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module adder8_16 ( out, a, b, cin );
  output [7:0] out;
  input [7:0] a;
  input [7:0] b;
  input cin;

  wire   [6:0] c;

  add_224 add_01 ( .s(out[0]), .a(a[0]), .b(b[0]), .ci(1'b0), .co(c[0]) );
  add_223 add_02 ( .s(out[1]), .a(a[1]), .b(b[1]), .ci(c[0]), .co(c[1]) );
  add_222 add_03 ( .s(out[2]), .a(a[2]), .b(b[2]), .ci(c[1]), .co(c[2]) );
  add_221 add_04 ( .s(out[3]), .a(a[3]), .b(b[3]), .ci(c[2]), .co(c[3]) );
  add_220 add_05 ( .s(out[4]), .a(a[4]), .b(b[4]), .ci(c[3]), .co(c[4]) );
  add_219 add_06 ( .s(out[5]), .a(a[5]), .b(b[5]), .ci(c[4]), .co(c[5]) );
  add_218 add_07 ( .s(out[6]), .a(a[6]), .b(b[6]), .ci(c[5]), .co(c[6]) );
  add_217 add_08 ( .s(out[7]), .a(a[7]), .b(b[7]), .ci(c[6]) );
endmodule


module floating_point_multiple_2 ( clk, rst_n, input_factor_01, 
        input_factor_02, output_multiply );
  input [31:0] input_factor_01;
  input [31:0] input_factor_02;
  output [31:0] output_multiply;
  input clk, rst_n;
  wire   N5, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22,
         N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N48, N49, N50, N51,
         N52, N53, N54, N55, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22,
         SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24,
         SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26;
  wire   [47:23] base_multiply_result;
  wire   [47:23] mulout;
  wire   [7:0] exponent_factor_12;
  wire   [7:0] pre_mul_output_exponent;

  mul26_2 mul26_01 ( .clk(clk), .rst_n(rst_n), .in1({1'b0, 1'b0, 1'b1, 
        input_factor_01[22:0]}), .in2({1'b0, 1'b0, 1'b1, input_factor_02[22:0]}), .en(1'b1), .mulout({SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, 
        SYNOPSYS_UNCONNECTED_3, mulout, SYNOPSYS_UNCONNECTED_4, 
        SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, 
        SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, 
        SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11, 
        SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13, 
        SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, 
        SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17, 
        SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19, 
        SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21, 
        SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_23, 
        SYNOPSYS_UNCONNECTED_24, SYNOPSYS_UNCONNECTED_25, 
        SYNOPSYS_UNCONNECTED_26}) );
  adder8_16 adder8_01 ( .out(exponent_factor_12), .a(input_factor_01[30:23]), 
        .b(input_factor_02[30:23]), .cin(1'b0) );
  adder8_15 adder8_02 ( .out(pre_mul_output_exponent), .a(exponent_factor_12), 
        .b({1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0}), .cin(1'b1) );
  DFFARX1 mul_output_sign_reg ( .D(N5), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[31]) );
  DFFARX1 base_multiply_result_reg_47_ ( .D(mulout[47]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[47]) );
  DFFARX1 base_multiply_result_reg_46_ ( .D(mulout[46]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[46]) );
  DFFARX1 base_multiply_result_reg_45_ ( .D(mulout[45]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[45]) );
  DFFARX1 base_multiply_result_reg_44_ ( .D(mulout[44]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[44]) );
  DFFARX1 base_multiply_result_reg_43_ ( .D(mulout[43]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[43]) );
  DFFARX1 base_multiply_result_reg_42_ ( .D(mulout[42]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[42]) );
  DFFARX1 base_multiply_result_reg_41_ ( .D(mulout[41]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[41]) );
  DFFARX1 base_multiply_result_reg_40_ ( .D(mulout[40]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[40]) );
  DFFARX1 base_multiply_result_reg_39_ ( .D(mulout[39]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[39]) );
  DFFARX1 base_multiply_result_reg_38_ ( .D(mulout[38]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[38]) );
  DFFARX1 base_multiply_result_reg_37_ ( .D(mulout[37]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[37]) );
  DFFARX1 base_multiply_result_reg_36_ ( .D(mulout[36]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[36]) );
  DFFARX1 base_multiply_result_reg_35_ ( .D(mulout[35]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[35]) );
  DFFARX1 base_multiply_result_reg_34_ ( .D(mulout[34]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[34]) );
  DFFARX1 base_multiply_result_reg_33_ ( .D(mulout[33]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[33]) );
  DFFARX1 base_multiply_result_reg_32_ ( .D(mulout[32]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[32]) );
  DFFARX1 base_multiply_result_reg_31_ ( .D(mulout[31]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[31]) );
  DFFARX1 base_multiply_result_reg_30_ ( .D(mulout[30]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[30]) );
  DFFARX1 base_multiply_result_reg_29_ ( .D(mulout[29]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[29]) );
  DFFARX1 base_multiply_result_reg_28_ ( .D(mulout[28]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[28]) );
  DFFARX1 base_multiply_result_reg_27_ ( .D(mulout[27]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[27]) );
  DFFARX1 base_multiply_result_reg_26_ ( .D(mulout[26]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[26]) );
  DFFARX1 base_multiply_result_reg_25_ ( .D(mulout[25]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[25]) );
  DFFARX1 base_multiply_result_reg_24_ ( .D(mulout[24]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[24]) );
  DFFARX1 base_multiply_result_reg_23_ ( .D(mulout[23]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[23]) );
  DFFARX1 mul_output_significand_reg_22_ ( .D(N32), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[22]) );
  DFFARX1 mul_output_significand_reg_21_ ( .D(N31), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[21]) );
  DFFARX1 mul_output_significand_reg_20_ ( .D(N30), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[20]) );
  DFFARX1 mul_output_significand_reg_19_ ( .D(N29), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[19]) );
  DFFARX1 mul_output_significand_reg_18_ ( .D(N28), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[18]) );
  DFFARX1 mul_output_significand_reg_17_ ( .D(N27), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[17]) );
  DFFARX1 mul_output_significand_reg_16_ ( .D(N26), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[16]) );
  DFFARX1 mul_output_significand_reg_15_ ( .D(N25), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[15]) );
  DFFARX1 mul_output_significand_reg_14_ ( .D(N24), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[14]) );
  DFFARX1 mul_output_significand_reg_13_ ( .D(N23), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[13]) );
  DFFARX1 mul_output_significand_reg_12_ ( .D(N22), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[12]) );
  DFFARX1 mul_output_significand_reg_11_ ( .D(N21), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[11]) );
  DFFARX1 mul_output_significand_reg_10_ ( .D(N20), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[10]) );
  DFFARX1 mul_output_significand_reg_9_ ( .D(N19), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[9]) );
  DFFARX1 mul_output_significand_reg_8_ ( .D(N18), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[8]) );
  DFFARX1 mul_output_significand_reg_7_ ( .D(N17), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[7]) );
  DFFARX1 mul_output_significand_reg_6_ ( .D(N16), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[6]) );
  DFFARX1 mul_output_significand_reg_5_ ( .D(N15), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[5]) );
  DFFARX1 mul_output_significand_reg_4_ ( .D(N14), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[4]) );
  DFFARX1 mul_output_significand_reg_3_ ( .D(N13), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[3]) );
  DFFARX1 mul_output_significand_reg_2_ ( .D(N12), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[2]) );
  DFFARX1 mul_output_significand_reg_1_ ( .D(N11), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[1]) );
  DFFARX1 mul_output_significand_reg_0_ ( .D(N10), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[0]) );
  DFFARX1 mul_output_exponent_reg_7_ ( .D(N55), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[30]) );
  DFFARX1 mul_output_exponent_reg_6_ ( .D(N54), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[29]) );
  DFFARX1 mul_output_exponent_reg_5_ ( .D(N53), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[28]) );
  DFFARX1 mul_output_exponent_reg_4_ ( .D(N52), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[27]) );
  DFFARX1 mul_output_exponent_reg_3_ ( .D(N51), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[26]) );
  DFFARX1 mul_output_exponent_reg_2_ ( .D(N50), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[25]) );
  DFFARX1 mul_output_exponent_reg_1_ ( .D(N49), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[24]) );
  DFFARX1 mul_output_exponent_reg_0_ ( .D(N48), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[23]) );
  AND2X1 U3 ( .IN1(base_multiply_result[47]), .IN2(n35), .Q(n32) );
  INVX0 U4 ( .INP(n1), .ZN(n2) );
  OR2X1 U5 ( .IN1(base_multiply_result[47]), .IN2(n24), .Q(n1) );
  INVX0 U6 ( .INP(input_factor_02[31]), .ZN(n3) );
  NOR4X0 U7 ( .IN1(input_factor_01[0]), .IN2(input_factor_01[10]), .IN3(
        input_factor_01[11]), .IN4(input_factor_01[12]), .QN(n7) );
  NOR4X0 U8 ( .IN1(input_factor_01[13]), .IN2(input_factor_01[14]), .IN3(
        input_factor_01[15]), .IN4(input_factor_01[16]), .QN(n6) );
  NOR4X0 U9 ( .IN1(input_factor_01[17]), .IN2(input_factor_01[18]), .IN3(
        input_factor_01[19]), .IN4(input_factor_01[1]), .QN(n5) );
  NOR4X0 U10 ( .IN1(input_factor_01[20]), .IN2(input_factor_01[21]), .IN3(
        input_factor_01[22]), .IN4(input_factor_01[23]), .QN(n4) );
  NAND4X0 U11 ( .IN1(n7), .IN2(n6), .IN3(n5), .IN4(n4), .QN(n23) );
  NOR4X0 U12 ( .IN1(input_factor_01[24]), .IN2(input_factor_01[25]), .IN3(
        input_factor_01[26]), .IN4(input_factor_01[27]), .QN(n11) );
  NOR4X0 U13 ( .IN1(input_factor_01[28]), .IN2(input_factor_01[29]), .IN3(
        input_factor_01[2]), .IN4(input_factor_01[30]), .QN(n10) );
  NOR4X0 U14 ( .IN1(input_factor_01[31]), .IN2(input_factor_01[3]), .IN3(
        input_factor_01[4]), .IN4(input_factor_01[5]), .QN(n9) );
  NOR4X0 U15 ( .IN1(input_factor_01[6]), .IN2(input_factor_01[7]), .IN3(
        input_factor_01[8]), .IN4(input_factor_01[9]), .QN(n8) );
  NAND4X0 U16 ( .IN1(n11), .IN2(n10), .IN3(n9), .IN4(n8), .QN(n22) );
  NOR4X0 U17 ( .IN1(input_factor_02[0]), .IN2(input_factor_02[10]), .IN3(
        input_factor_02[11]), .IN4(input_factor_02[12]), .QN(n15) );
  NOR4X0 U18 ( .IN1(input_factor_02[13]), .IN2(input_factor_02[14]), .IN3(
        input_factor_02[15]), .IN4(input_factor_02[16]), .QN(n14) );
  NOR4X0 U19 ( .IN1(input_factor_02[17]), .IN2(input_factor_02[18]), .IN3(
        input_factor_02[19]), .IN4(input_factor_02[1]), .QN(n13) );
  NOR4X0 U20 ( .IN1(input_factor_02[20]), .IN2(input_factor_02[21]), .IN3(
        input_factor_02[22]), .IN4(input_factor_02[23]), .QN(n12) );
  NAND4X0 U21 ( .IN1(n15), .IN2(n14), .IN3(n13), .IN4(n12), .QN(n21) );
  NOR4X0 U22 ( .IN1(input_factor_02[24]), .IN2(input_factor_02[25]), .IN3(
        input_factor_02[26]), .IN4(input_factor_02[27]), .QN(n19) );
  NOR4X0 U23 ( .IN1(input_factor_02[28]), .IN2(input_factor_02[29]), .IN3(
        input_factor_02[2]), .IN4(input_factor_02[30]), .QN(n18) );
  NOR4X0 U24 ( .IN1(input_factor_02[31]), .IN2(input_factor_02[3]), .IN3(
        input_factor_02[4]), .IN4(input_factor_02[5]), .QN(n17) );
  NOR4X0 U25 ( .IN1(input_factor_02[6]), .IN2(input_factor_02[7]), .IN3(
        input_factor_02[8]), .IN4(input_factor_02[9]), .QN(n16) );
  NAND4X0 U26 ( .IN1(n19), .IN2(n18), .IN3(n17), .IN4(n16), .QN(n20) );
  OA22X1 U27 ( .IN1(n23), .IN2(n22), .IN3(n21), .IN4(n20), .Q(n35) );
  INVX0 U28 ( .INP(n35), .ZN(n24) );
  AO22X1 U29 ( .IN1(n2), .IN2(base_multiply_result[23]), .IN3(n32), .IN4(
        base_multiply_result[24]), .Q(N10) );
  AO22X1 U30 ( .IN1(n2), .IN2(base_multiply_result[24]), .IN3(n32), .IN4(
        base_multiply_result[25]), .Q(N11) );
  AO22X1 U31 ( .IN1(n2), .IN2(base_multiply_result[25]), .IN3(n32), .IN4(
        base_multiply_result[26]), .Q(N12) );
  AO22X1 U32 ( .IN1(n2), .IN2(base_multiply_result[26]), .IN3(n32), .IN4(
        base_multiply_result[27]), .Q(N13) );
  AO22X1 U33 ( .IN1(n2), .IN2(base_multiply_result[27]), .IN3(n32), .IN4(
        base_multiply_result[28]), .Q(N14) );
  AO22X1 U34 ( .IN1(n2), .IN2(base_multiply_result[28]), .IN3(n32), .IN4(
        base_multiply_result[29]), .Q(N15) );
  AO22X1 U35 ( .IN1(n2), .IN2(base_multiply_result[29]), .IN3(n32), .IN4(
        base_multiply_result[30]), .Q(N16) );
  AO22X1 U36 ( .IN1(n2), .IN2(base_multiply_result[30]), .IN3(n32), .IN4(
        base_multiply_result[31]), .Q(N17) );
  AO22X1 U37 ( .IN1(n2), .IN2(base_multiply_result[31]), .IN3(n32), .IN4(
        base_multiply_result[32]), .Q(N18) );
  AO22X1 U38 ( .IN1(n2), .IN2(base_multiply_result[32]), .IN3(n32), .IN4(
        base_multiply_result[33]), .Q(N19) );
  AO22X1 U39 ( .IN1(n2), .IN2(base_multiply_result[33]), .IN3(n32), .IN4(
        base_multiply_result[34]), .Q(N20) );
  AO22X1 U40 ( .IN1(n2), .IN2(base_multiply_result[34]), .IN3(n32), .IN4(
        base_multiply_result[35]), .Q(N21) );
  AO22X1 U41 ( .IN1(n2), .IN2(base_multiply_result[35]), .IN3(n32), .IN4(
        base_multiply_result[36]), .Q(N22) );
  AO22X1 U42 ( .IN1(n2), .IN2(base_multiply_result[36]), .IN3(n32), .IN4(
        base_multiply_result[37]), .Q(N23) );
  AO22X1 U43 ( .IN1(n2), .IN2(base_multiply_result[37]), .IN3(n32), .IN4(
        base_multiply_result[38]), .Q(N24) );
  AO22X1 U44 ( .IN1(n2), .IN2(base_multiply_result[38]), .IN3(n32), .IN4(
        base_multiply_result[39]), .Q(N25) );
  AO22X1 U45 ( .IN1(n2), .IN2(base_multiply_result[39]), .IN3(n32), .IN4(
        base_multiply_result[40]), .Q(N26) );
  AO22X1 U46 ( .IN1(n2), .IN2(base_multiply_result[40]), .IN3(n32), .IN4(
        base_multiply_result[41]), .Q(N27) );
  AO22X1 U47 ( .IN1(n2), .IN2(base_multiply_result[41]), .IN3(n32), .IN4(
        base_multiply_result[42]), .Q(N28) );
  AO22X1 U48 ( .IN1(n2), .IN2(base_multiply_result[42]), .IN3(n32), .IN4(
        base_multiply_result[43]), .Q(N29) );
  AO22X1 U49 ( .IN1(n2), .IN2(base_multiply_result[43]), .IN3(n32), .IN4(
        base_multiply_result[44]), .Q(N30) );
  AO22X1 U50 ( .IN1(n2), .IN2(base_multiply_result[44]), .IN3(n32), .IN4(
        base_multiply_result[45]), .Q(N31) );
  AO22X1 U51 ( .IN1(n2), .IN2(base_multiply_result[45]), .IN3(n32), .IN4(
        base_multiply_result[46]), .Q(N32) );
  MUX21X1 U52 ( .IN1(n2), .IN2(n32), .S(pre_mul_output_exponent[0]), .Q(N48)
         );
  AO21X1 U53 ( .IN1(pre_mul_output_exponent[0]), .IN2(n2), .IN3(n32), .Q(n25)
         );
  NOR3X0 U54 ( .IN1(pre_mul_output_exponent[1]), .IN2(
        pre_mul_output_exponent[0]), .IN3(n1), .QN(n27) );
  AO21X1 U55 ( .IN1(pre_mul_output_exponent[1]), .IN2(n25), .IN3(n27), .Q(N49)
         );
  INVX0 U56 ( .INP(input_factor_01[31]), .ZN(n26) );
  OA221X1 U57 ( .IN1(input_factor_01[31]), .IN2(input_factor_02[31]), .IN3(n26), .IN4(n3), .IN5(n35), .Q(N5) );
  AO221X1 U58 ( .IN1(n2), .IN2(pre_mul_output_exponent[1]), .IN3(n2), .IN4(
        pre_mul_output_exponent[0]), .IN5(n32), .Q(n28) );
  MUX21X1 U59 ( .IN1(n27), .IN2(n28), .S(pre_mul_output_exponent[2]), .Q(N50)
         );
  AND2X1 U60 ( .IN1(n2), .IN2(pre_mul_output_exponent[2]), .Q(n29) );
  OR4X1 U61 ( .IN1(pre_mul_output_exponent[1]), .IN2(
        pre_mul_output_exponent[0]), .IN3(pre_mul_output_exponent[3]), .IN4(
        pre_mul_output_exponent[2]), .Q(n34) );
  NOR2X0 U62 ( .IN1(n1), .IN2(n34), .QN(n31) );
  AO221X1 U63 ( .IN1(pre_mul_output_exponent[3]), .IN2(n29), .IN3(
        pre_mul_output_exponent[3]), .IN4(n28), .IN5(n31), .Q(N51) );
  OA21X1 U64 ( .IN1(base_multiply_result[47]), .IN2(n34), .IN3(n35), .Q(n30)
         );
  MUX21X1 U65 ( .IN1(n31), .IN2(n30), .S(pre_mul_output_exponent[4]), .Q(N52)
         );
  AO221X1 U66 ( .IN1(n2), .IN2(pre_mul_output_exponent[4]), .IN3(n2), .IN4(n34), .IN5(n32), .Q(n33) );
  NOR4X0 U67 ( .IN1(pre_mul_output_exponent[5]), .IN2(
        pre_mul_output_exponent[4]), .IN3(n34), .IN4(n1), .QN(n37) );
  AO21X1 U68 ( .IN1(pre_mul_output_exponent[5]), .IN2(n33), .IN3(n37), .Q(N53)
         );
  OR3X1 U69 ( .IN1(pre_mul_output_exponent[5]), .IN2(
        pre_mul_output_exponent[4]), .IN3(n34), .Q(n36) );
  OA21X1 U70 ( .IN1(base_multiply_result[47]), .IN2(n36), .IN3(n35), .Q(n39)
         );
  INVX0 U71 ( .INP(n37), .ZN(n38) );
  NOR2X0 U72 ( .IN1(pre_mul_output_exponent[6]), .IN2(n38), .QN(n41) );
  AO21X1 U73 ( .IN1(pre_mul_output_exponent[6]), .IN2(n39), .IN3(n41), .Q(N54)
         );
  AO21X1 U74 ( .IN1(n2), .IN2(pre_mul_output_exponent[6]), .IN3(n39), .Q(n40)
         );
  MUX21X1 U75 ( .IN1(n41), .IN2(n40), .S(pre_mul_output_exponent[7]), .Q(N55)
         );
endmodule


module cla51squ_3 ( out, a, b );
  output [50:0] out;
  input [50:0] a;
  input [50:0] b;
  wire   intadd_3_CI, intadd_3_n24, intadd_3_n23, intadd_3_n22, intadd_3_n21,
         intadd_3_n20, intadd_3_n19, intadd_3_n18, intadd_3_n17, intadd_3_n16,
         intadd_3_n15, intadd_3_n14, intadd_3_n13, intadd_3_n12, intadd_3_n11,
         intadd_3_n10, intadd_3_n9, intadd_3_n8, intadd_3_n7, intadd_3_n6,
         intadd_3_n5, intadd_3_n4, intadd_3_n3, intadd_3_n2, intadd_3_n1, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14;

  FADDX1 intadd_3_U25 ( .A(b[23]), .B(a[23]), .CI(intadd_3_CI), .CO(
        intadd_3_n24), .S(out[23]) );
  FADDX1 intadd_3_U24 ( .A(b[24]), .B(a[24]), .CI(intadd_3_n24), .CO(
        intadd_3_n23), .S(out[24]) );
  FADDX1 intadd_3_U23 ( .A(b[25]), .B(a[25]), .CI(intadd_3_n23), .CO(
        intadd_3_n22), .S(out[25]) );
  FADDX1 intadd_3_U22 ( .A(b[26]), .B(a[26]), .CI(intadd_3_n22), .CO(
        intadd_3_n21), .S(out[26]) );
  FADDX1 intadd_3_U21 ( .A(b[27]), .B(a[27]), .CI(intadd_3_n21), .CO(
        intadd_3_n20), .S(out[27]) );
  FADDX1 intadd_3_U20 ( .A(b[28]), .B(a[28]), .CI(intadd_3_n20), .CO(
        intadd_3_n19), .S(out[28]) );
  FADDX1 intadd_3_U19 ( .A(b[29]), .B(a[29]), .CI(intadd_3_n19), .CO(
        intadd_3_n18), .S(out[29]) );
  FADDX1 intadd_3_U18 ( .A(b[30]), .B(a[30]), .CI(intadd_3_n18), .CO(
        intadd_3_n17), .S(out[30]) );
  FADDX1 intadd_3_U17 ( .A(b[31]), .B(a[31]), .CI(intadd_3_n17), .CO(
        intadd_3_n16), .S(out[31]) );
  FADDX1 intadd_3_U16 ( .A(b[32]), .B(a[32]), .CI(intadd_3_n16), .CO(
        intadd_3_n15), .S(out[32]) );
  FADDX1 intadd_3_U15 ( .A(b[33]), .B(a[33]), .CI(intadd_3_n15), .CO(
        intadd_3_n14), .S(out[33]) );
  FADDX1 intadd_3_U14 ( .A(b[34]), .B(a[34]), .CI(intadd_3_n14), .CO(
        intadd_3_n13), .S(out[34]) );
  FADDX1 intadd_3_U13 ( .A(b[35]), .B(a[35]), .CI(intadd_3_n13), .CO(
        intadd_3_n12), .S(out[35]) );
  FADDX1 intadd_3_U12 ( .A(b[36]), .B(a[36]), .CI(intadd_3_n12), .CO(
        intadd_3_n11), .S(out[36]) );
  FADDX1 intadd_3_U11 ( .A(b[37]), .B(a[37]), .CI(intadd_3_n11), .CO(
        intadd_3_n10), .S(out[37]) );
  FADDX1 intadd_3_U10 ( .A(b[38]), .B(a[38]), .CI(intadd_3_n10), .CO(
        intadd_3_n9), .S(out[38]) );
  FADDX1 intadd_3_U9 ( .A(b[39]), .B(a[39]), .CI(intadd_3_n9), .CO(intadd_3_n8), .S(out[39]) );
  FADDX1 intadd_3_U8 ( .A(b[40]), .B(a[40]), .CI(intadd_3_n8), .CO(intadd_3_n7), .S(out[40]) );
  FADDX1 intadd_3_U7 ( .A(b[41]), .B(a[41]), .CI(intadd_3_n7), .CO(intadd_3_n6), .S(out[41]) );
  FADDX1 intadd_3_U6 ( .A(b[42]), .B(a[42]), .CI(intadd_3_n6), .CO(intadd_3_n5), .S(out[42]) );
  FADDX1 intadd_3_U5 ( .A(b[43]), .B(a[43]), .CI(intadd_3_n5), .CO(intadd_3_n4), .S(out[43]) );
  FADDX1 intadd_3_U4 ( .A(b[44]), .B(a[44]), .CI(intadd_3_n4), .CO(intadd_3_n3), .S(out[44]) );
  FADDX1 intadd_3_U3 ( .A(b[45]), .B(a[45]), .CI(intadd_3_n3), .CO(intadd_3_n2), .S(out[45]) );
  FADDX1 intadd_3_U2 ( .A(b[46]), .B(a[46]), .CI(intadd_3_n2), .CO(intadd_3_n1), .S(out[46]) );
  OA21X1 U2 ( .IN1(b[9]), .IN2(a[9]), .IN3(a[8]), .Q(n1) );
  AO22X1 U3 ( .IN1(b[9]), .IN2(a[9]), .IN3(b[8]), .IN4(n1), .Q(n2) );
  AO222X1 U4 ( .IN1(b[10]), .IN2(a[10]), .IN3(b[10]), .IN4(n2), .IN5(a[10]), 
        .IN6(n2), .Q(n3) );
  AO222X1 U5 ( .IN1(b[11]), .IN2(a[11]), .IN3(b[11]), .IN4(n3), .IN5(a[11]), 
        .IN6(n3), .Q(n4) );
  AO222X1 U6 ( .IN1(b[12]), .IN2(a[12]), .IN3(b[12]), .IN4(n4), .IN5(a[12]), 
        .IN6(n4), .Q(n5) );
  AO222X1 U7 ( .IN1(b[13]), .IN2(a[13]), .IN3(b[13]), .IN4(n5), .IN5(a[13]), 
        .IN6(n5), .Q(n6) );
  AO222X1 U8 ( .IN1(b[14]), .IN2(a[14]), .IN3(b[14]), .IN4(n6), .IN5(a[14]), 
        .IN6(n6), .Q(n7) );
  AO222X1 U9 ( .IN1(b[15]), .IN2(a[15]), .IN3(b[15]), .IN4(n7), .IN5(a[15]), 
        .IN6(n7), .Q(n8) );
  AO222X1 U10 ( .IN1(b[16]), .IN2(a[16]), .IN3(b[16]), .IN4(n8), .IN5(a[16]), 
        .IN6(n8), .Q(n9) );
  AO222X1 U11 ( .IN1(b[17]), .IN2(a[17]), .IN3(b[17]), .IN4(n9), .IN5(a[17]), 
        .IN6(n9), .Q(n10) );
  AO222X1 U12 ( .IN1(b[18]), .IN2(a[18]), .IN3(b[18]), .IN4(n10), .IN5(a[18]), 
        .IN6(n10), .Q(n11) );
  AO222X1 U13 ( .IN1(b[19]), .IN2(a[19]), .IN3(b[19]), .IN4(n11), .IN5(a[19]), 
        .IN6(n11), .Q(n12) );
  AO222X1 U14 ( .IN1(b[20]), .IN2(a[20]), .IN3(b[20]), .IN4(n12), .IN5(a[20]), 
        .IN6(n12), .Q(n13) );
  AO222X1 U15 ( .IN1(b[21]), .IN2(a[21]), .IN3(b[21]), .IN4(n13), .IN5(a[21]), 
        .IN6(n13), .Q(n14) );
  AO222X1 U16 ( .IN1(b[22]), .IN2(a[22]), .IN3(b[22]), .IN4(n14), .IN5(a[22]), 
        .IN6(n14), .Q(intadd_3_CI) );
  XOR3X1 U17 ( .IN1(intadd_3_n1), .IN2(a[47]), .IN3(b[47]), .Q(out[47]) );
endmodule


module csa51squ_25 ( sumout, in1, in2, in3, cout_50_, cout_49_, cout_48_, 
        cout_47_, cout_46_, cout_44_, cout_42_, cout_40_, cout_38_, cout_36_, 
        cout_34_, cout_32_, cout_30_, cout_28_, cout_27_, cout_7__BAR, cout_6_, 
        cout_5_, cout_4_, cout_3_, cout_2_, cout_1_, cout_0_, cout_8__BAR, 
        cout_9__BAR, cout_10__BAR, cout_11__BAR, cout_12__BAR, cout_13__BAR, 
        cout_14__BAR, cout_15__BAR, cout_16__BAR, cout_17__BAR, cout_18__BAR, 
        cout_19__BAR, cout_20__BAR, cout_21__BAR, cout_22__BAR, cout_23__BAR, 
        cout_24__BAR, cout_25__BAR, cout_26__BAR, cout_29__BAR, cout_31__BAR, 
        cout_33__BAR, cout_35__BAR, cout_37__BAR, cout_39__BAR, cout_41__BAR, 
        cout_43__BAR, cout_45__BAR );
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  output cout_50_, cout_49_, cout_48_, cout_47_, cout_46_, cout_44_, cout_42_,
         cout_40_, cout_38_, cout_36_, cout_34_, cout_32_, cout_30_, cout_28_,
         cout_27_, cout_7__BAR, cout_6_, cout_5_, cout_4_, cout_3_, cout_2_,
         cout_1_, cout_0_, cout_8__BAR, cout_9__BAR, cout_10__BAR,
         cout_11__BAR, cout_12__BAR, cout_13__BAR, cout_14__BAR, cout_15__BAR,
         cout_16__BAR, cout_17__BAR, cout_18__BAR, cout_19__BAR, cout_20__BAR,
         cout_21__BAR, cout_22__BAR, cout_23__BAR, cout_24__BAR, cout_25__BAR,
         cout_26__BAR, cout_29__BAR, cout_31__BAR, cout_33__BAR, cout_35__BAR,
         cout_37__BAR, cout_39__BAR, cout_41__BAR, cout_43__BAR, cout_45__BAR;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11;

  NAND2X0 U1 ( .IN1(in2[8]), .IN2(in1[8]), .QN(cout_8__BAR) );
  NAND2X0 U2 ( .IN1(in2[9]), .IN2(in1[9]), .QN(cout_9__BAR) );
  NAND2X0 U3 ( .IN1(in2[10]), .IN2(in1[10]), .QN(cout_10__BAR) );
  NAND2X0 U4 ( .IN1(in2[11]), .IN2(in1[11]), .QN(cout_11__BAR) );
  NAND2X0 U5 ( .IN1(in2[12]), .IN2(in1[12]), .QN(cout_12__BAR) );
  NAND2X0 U6 ( .IN1(in2[13]), .IN2(in1[13]), .QN(cout_13__BAR) );
  NAND2X0 U7 ( .IN1(in2[14]), .IN2(in1[14]), .QN(cout_14__BAR) );
  NAND2X0 U8 ( .IN1(in2[15]), .IN2(in1[15]), .QN(cout_15__BAR) );
  NAND2X0 U9 ( .IN1(in2[16]), .IN2(in1[16]), .QN(cout_16__BAR) );
  NAND2X0 U10 ( .IN1(in2[17]), .IN2(in1[17]), .QN(cout_17__BAR) );
  NAND2X0 U11 ( .IN1(in2[18]), .IN2(in1[18]), .QN(cout_18__BAR) );
  NAND2X0 U12 ( .IN1(in2[19]), .IN2(in1[19]), .QN(cout_19__BAR) );
  NAND2X0 U13 ( .IN1(in2[20]), .IN2(in1[20]), .QN(cout_20__BAR) );
  NAND2X0 U14 ( .IN1(in2[21]), .IN2(in1[21]), .QN(cout_21__BAR) );
  NAND2X0 U15 ( .IN1(in2[22]), .IN2(in1[22]), .QN(cout_22__BAR) );
  NAND2X0 U16 ( .IN1(in2[23]), .IN2(in1[23]), .QN(cout_23__BAR) );
  NAND2X0 U17 ( .IN1(in2[24]), .IN2(in1[24]), .QN(cout_24__BAR) );
  NAND2X0 U18 ( .IN1(in2[25]), .IN2(in1[25]), .QN(cout_25__BAR) );
  NAND2X0 U19 ( .IN1(in2[26]), .IN2(in1[26]), .QN(cout_26__BAR) );
  NAND2X0 U20 ( .IN1(in2[29]), .IN2(in1[29]), .QN(cout_29__BAR) );
  NAND2X0 U21 ( .IN1(in2[31]), .IN2(in1[31]), .QN(cout_31__BAR) );
  NAND2X0 U22 ( .IN1(in2[33]), .IN2(in1[33]), .QN(cout_33__BAR) );
  NAND2X0 U23 ( .IN1(in2[35]), .IN2(in1[35]), .QN(cout_35__BAR) );
  NAND2X0 U24 ( .IN1(in2[37]), .IN2(in1[37]), .QN(cout_37__BAR) );
  NAND2X0 U25 ( .IN1(in2[39]), .IN2(in1[39]), .QN(cout_39__BAR) );
  NAND2X0 U26 ( .IN1(in2[41]), .IN2(in1[41]), .QN(cout_41__BAR) );
  NAND2X0 U27 ( .IN1(in2[43]), .IN2(in1[43]), .QN(cout_43__BAR) );
  NAND2X0 U28 ( .IN1(in2[45]), .IN2(in1[45]), .QN(cout_45__BAR) );
  NAND2X0 U29 ( .IN1(in2[7]), .IN2(in1[7]), .QN(cout_7__BAR) );
  NAND2X0 U30 ( .IN1(n1), .IN2(cout_27_), .QN(sumout[27]) );
  NAND2X0 U31 ( .IN1(in1[27]), .IN2(in2[27]), .QN(n1) );
  NAND2X0 U32 ( .IN1(n2), .IN2(cout_28_), .QN(sumout[28]) );
  NAND2X0 U33 ( .IN1(in1[28]), .IN2(in2[28]), .QN(n2) );
  NAND2X0 U34 ( .IN1(n3), .IN2(cout_30_), .QN(sumout[30]) );
  NAND2X0 U35 ( .IN1(in1[30]), .IN2(in2[30]), .QN(n3) );
  NAND2X0 U36 ( .IN1(n4), .IN2(cout_32_), .QN(sumout[32]) );
  NAND2X0 U37 ( .IN1(in1[32]), .IN2(in2[32]), .QN(n4) );
  NAND2X0 U38 ( .IN1(n5), .IN2(cout_34_), .QN(sumout[34]) );
  NAND2X0 U39 ( .IN1(in1[34]), .IN2(in2[34]), .QN(n5) );
  NAND2X0 U40 ( .IN1(n6), .IN2(cout_36_), .QN(sumout[36]) );
  NAND2X0 U41 ( .IN1(in1[36]), .IN2(in2[36]), .QN(n6) );
  NAND2X0 U42 ( .IN1(n7), .IN2(cout_38_), .QN(sumout[38]) );
  NAND2X0 U43 ( .IN1(in1[38]), .IN2(in2[38]), .QN(n7) );
  NAND2X0 U44 ( .IN1(n8), .IN2(cout_40_), .QN(sumout[40]) );
  NAND2X0 U45 ( .IN1(in1[40]), .IN2(in2[40]), .QN(n8) );
  NAND2X0 U46 ( .IN1(n9), .IN2(cout_42_), .QN(sumout[42]) );
  NAND2X0 U47 ( .IN1(in1[42]), .IN2(in2[42]), .QN(n9) );
  NAND2X0 U48 ( .IN1(n10), .IN2(cout_44_), .QN(sumout[44]) );
  NAND2X0 U49 ( .IN1(in1[44]), .IN2(in2[44]), .QN(n10) );
  NAND2X0 U50 ( .IN1(n11), .IN2(cout_46_), .QN(sumout[46]) );
  NAND2X0 U51 ( .IN1(in1[46]), .IN2(in2[46]), .QN(n11) );
  OR2X1 U52 ( .IN1(in2[27]), .IN2(in1[27]), .Q(cout_27_) );
  OR2X1 U53 ( .IN1(in2[28]), .IN2(in1[28]), .Q(cout_28_) );
  OR2X1 U54 ( .IN1(in2[30]), .IN2(in1[30]), .Q(cout_30_) );
  OR2X1 U55 ( .IN1(in2[32]), .IN2(in1[32]), .Q(cout_32_) );
  OR2X1 U56 ( .IN1(in2[34]), .IN2(in1[34]), .Q(cout_34_) );
  OR2X1 U57 ( .IN1(in2[36]), .IN2(in1[36]), .Q(cout_36_) );
  OR2X1 U58 ( .IN1(in2[38]), .IN2(in1[38]), .Q(cout_38_) );
  OR2X1 U59 ( .IN1(in2[40]), .IN2(in1[40]), .Q(cout_40_) );
  OR2X1 U60 ( .IN1(in2[42]), .IN2(in1[42]), .Q(cout_42_) );
  OR2X1 U61 ( .IN1(in2[44]), .IN2(in1[44]), .Q(cout_44_) );
  OR2X1 U62 ( .IN1(in2[46]), .IN2(in1[46]), .Q(cout_46_) );
  OA21X1 U63 ( .IN1(in2[8]), .IN2(in1[8]), .IN3(cout_8__BAR), .Q(sumout[8]) );
  OA21X1 U64 ( .IN1(in2[9]), .IN2(in1[9]), .IN3(cout_9__BAR), .Q(sumout[9]) );
  OA21X1 U65 ( .IN1(in2[10]), .IN2(in1[10]), .IN3(cout_10__BAR), .Q(sumout[10]) );
  OA21X1 U66 ( .IN1(in2[11]), .IN2(in1[11]), .IN3(cout_11__BAR), .Q(sumout[11]) );
  OA21X1 U67 ( .IN1(in2[12]), .IN2(in1[12]), .IN3(cout_12__BAR), .Q(sumout[12]) );
  OA21X1 U68 ( .IN1(in2[13]), .IN2(in1[13]), .IN3(cout_13__BAR), .Q(sumout[13]) );
  OA21X1 U69 ( .IN1(in2[14]), .IN2(in1[14]), .IN3(cout_14__BAR), .Q(sumout[14]) );
  OA21X1 U70 ( .IN1(in2[15]), .IN2(in1[15]), .IN3(cout_15__BAR), .Q(sumout[15]) );
  OA21X1 U71 ( .IN1(in2[16]), .IN2(in1[16]), .IN3(cout_16__BAR), .Q(sumout[16]) );
  OA21X1 U72 ( .IN1(in2[17]), .IN2(in1[17]), .IN3(cout_17__BAR), .Q(sumout[17]) );
  OA21X1 U73 ( .IN1(in2[18]), .IN2(in1[18]), .IN3(cout_18__BAR), .Q(sumout[18]) );
  OA21X1 U74 ( .IN1(in2[19]), .IN2(in1[19]), .IN3(cout_19__BAR), .Q(sumout[19]) );
  OA21X1 U75 ( .IN1(in2[20]), .IN2(in1[20]), .IN3(cout_20__BAR), .Q(sumout[20]) );
  OA21X1 U76 ( .IN1(in2[21]), .IN2(in1[21]), .IN3(cout_21__BAR), .Q(sumout[21]) );
  OA21X1 U77 ( .IN1(in2[22]), .IN2(in1[22]), .IN3(cout_22__BAR), .Q(sumout[22]) );
  OA21X1 U78 ( .IN1(in2[23]), .IN2(in1[23]), .IN3(cout_23__BAR), .Q(sumout[23]) );
  OA21X1 U79 ( .IN1(in2[24]), .IN2(in1[24]), .IN3(cout_24__BAR), .Q(sumout[24]) );
  OA21X1 U80 ( .IN1(in2[25]), .IN2(in1[25]), .IN3(cout_25__BAR), .Q(sumout[25]) );
  OA21X1 U81 ( .IN1(in2[26]), .IN2(in1[26]), .IN3(cout_26__BAR), .Q(sumout[26]) );
  OA21X1 U82 ( .IN1(in2[29]), .IN2(in1[29]), .IN3(cout_29__BAR), .Q(sumout[29]) );
  OA21X1 U83 ( .IN1(in2[31]), .IN2(in1[31]), .IN3(cout_31__BAR), .Q(sumout[31]) );
  OA21X1 U84 ( .IN1(in2[33]), .IN2(in1[33]), .IN3(cout_33__BAR), .Q(sumout[33]) );
  OA21X1 U85 ( .IN1(in2[35]), .IN2(in1[35]), .IN3(cout_35__BAR), .Q(sumout[35]) );
  OA21X1 U86 ( .IN1(in2[37]), .IN2(in1[37]), .IN3(cout_37__BAR), .Q(sumout[37]) );
  OA21X1 U87 ( .IN1(in2[39]), .IN2(in1[39]), .IN3(cout_39__BAR), .Q(sumout[39]) );
  OA21X1 U88 ( .IN1(in2[41]), .IN2(in1[41]), .IN3(cout_41__BAR), .Q(sumout[41]) );
  OA21X1 U89 ( .IN1(in2[43]), .IN2(in1[43]), .IN3(cout_43__BAR), .Q(sumout[43]) );
  OA21X1 U90 ( .IN1(in2[45]), .IN2(in1[45]), .IN3(cout_45__BAR), .Q(sumout[45]) );
  XOR2X1 U91 ( .IN1(in1[47]), .IN2(in2[47]), .Q(sumout[47]) );
endmodule


module csa51squ_26 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;


  AO222X1 U1 ( .IN1(in2[6]), .IN2(in3[6]), .IN3(in2[6]), .IN4(in1[6]), .IN5(
        in3[6]), .IN6(in1[6]), .Q(cout[6]) );
  FADDX1 U2 ( .A(in1[10]), .B(in2[10]), .CI(in3[10]), .CO(cout[10]), .S(
        sumout[10]) );
  FADDX1 U3 ( .A(in1[11]), .B(in2[11]), .CI(in3[11]), .CO(cout[11]), .S(
        sumout[11]) );
  FADDX1 U4 ( .A(in1[12]), .B(in2[12]), .CI(in3[12]), .CO(cout[12]), .S(
        sumout[12]) );
  FADDX1 U5 ( .A(in1[13]), .B(in2[13]), .CI(in3[13]), .CO(cout[13]), .S(
        sumout[13]) );
  FADDX1 U6 ( .A(in1[14]), .B(in2[14]), .CI(in3[14]), .CO(cout[14]), .S(
        sumout[14]) );
  FADDX1 U7 ( .A(in1[15]), .B(in2[15]), .CI(in3[15]), .CO(cout[15]), .S(
        sumout[15]) );
  FADDX1 U8 ( .A(in1[16]), .B(in2[16]), .CI(in3[16]), .CO(cout[16]), .S(
        sumout[16]) );
  FADDX1 U9 ( .A(in1[17]), .B(in2[17]), .CI(in3[17]), .CO(cout[17]), .S(
        sumout[17]) );
  FADDX1 U10 ( .A(in1[18]), .B(in2[18]), .CI(in3[18]), .CO(cout[18]), .S(
        sumout[18]) );
  FADDX1 U11 ( .A(in1[19]), .B(in2[19]), .CI(in3[19]), .CO(cout[19]), .S(
        sumout[19]) );
  FADDX1 U12 ( .A(in1[20]), .B(in2[20]), .CI(in3[20]), .CO(cout[20]), .S(
        sumout[20]) );
  FADDX1 U13 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U14 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U15 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U16 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U17 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U18 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U19 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U20 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U21 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U22 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U23 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U24 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
  FADDX1 U25 ( .A(in1[33]), .B(in2[33]), .CI(in3[33]), .CO(cout[33]), .S(
        sumout[33]) );
  FADDX1 U26 ( .A(in1[34]), .B(in2[34]), .CI(in3[34]), .CO(cout[34]), .S(
        sumout[34]) );
  FADDX1 U27 ( .A(in1[35]), .B(in2[35]), .CI(in3[35]), .CO(cout[35]), .S(
        sumout[35]) );
  FADDX1 U28 ( .A(in1[36]), .B(in2[36]), .CI(in3[36]), .CO(cout[36]), .S(
        sumout[36]) );
  FADDX1 U29 ( .A(in1[37]), .B(in2[37]), .CI(in3[37]), .CO(cout[37]), .S(
        sumout[37]) );
  FADDX1 U30 ( .A(in1[38]), .B(in2[38]), .CI(in3[38]), .CO(cout[38]), .S(
        sumout[38]) );
  FADDX1 U31 ( .A(in1[39]), .B(in2[39]), .CI(in3[39]), .CO(cout[39]), .S(
        sumout[39]) );
  FADDX1 U32 ( .A(in1[40]), .B(in2[40]), .CI(in3[40]), .CO(cout[40]), .S(
        sumout[40]) );
  FADDX1 U33 ( .A(in1[41]), .B(in2[41]), .CI(in3[41]), .CO(cout[41]), .S(
        sumout[41]) );
  FADDX1 U34 ( .A(in1[42]), .B(in2[42]), .CI(in3[42]), .CO(cout[42]), .S(
        sumout[42]) );
  FADDX1 U35 ( .A(in1[43]), .B(in2[43]), .CI(in3[43]), .CO(cout[43]), .S(
        sumout[43]) );
  FADDX1 U36 ( .A(in1[44]), .B(in2[44]), .CI(in3[44]), .CO(cout[44]), .S(
        sumout[44]) );
  FADDX1 U37 ( .A(in1[45]), .B(in2[45]), .CI(in3[45]), .CO(cout[45]), .S(
        sumout[45]) );
  FADDX1 U38 ( .A(in1[46]), .B(in2[46]), .CI(in3[46]), .CO(cout[46]), .S(
        sumout[46]) );
  XOR3X1 U39 ( .IN1(in2[47]), .IN2(in3[47]), .IN3(in1[47]), .Q(sumout[47]) );
  FADDX1 U40 ( .A(in1[7]), .B(in2[7]), .CI(in3[7]), .CO(cout[7]), .S(sumout[7]) );
  FADDX1 U41 ( .A(in1[8]), .B(in2[8]), .CI(in3[8]), .CO(cout[8]), .S(sumout[8]) );
  FADDX1 U42 ( .A(in1[9]), .B(in2[9]), .CI(in3[9]), .CO(cout[9]), .S(sumout[9]) );
endmodule


module csa51squ_27 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14;

  AND2X1 U1 ( .IN1(in2[7]), .IN2(in1[7]), .Q(cout[7]) );
  NOR2X0 U2 ( .IN1(in2[7]), .IN2(in1[7]), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(cout[7]), .QN(sumout[7]) );
  AND2X1 U4 ( .IN1(in2[8]), .IN2(in1[8]), .Q(cout[8]) );
  NOR2X0 U5 ( .IN1(in2[8]), .IN2(in1[8]), .QN(n2) );
  NOR2X0 U6 ( .IN1(n2), .IN2(cout[8]), .QN(sumout[8]) );
  AND2X1 U7 ( .IN1(in2[9]), .IN2(in1[9]), .Q(cout[9]) );
  NOR2X0 U8 ( .IN1(in2[9]), .IN2(in1[9]), .QN(n3) );
  NOR2X0 U9 ( .IN1(n3), .IN2(cout[9]), .QN(sumout[9]) );
  AND2X1 U10 ( .IN1(in2[10]), .IN2(in1[10]), .Q(cout[10]) );
  NOR2X0 U11 ( .IN1(in2[10]), .IN2(in1[10]), .QN(n4) );
  NOR2X0 U12 ( .IN1(n4), .IN2(cout[10]), .QN(sumout[10]) );
  AND2X1 U13 ( .IN1(in2[11]), .IN2(in1[11]), .Q(cout[11]) );
  NOR2X0 U14 ( .IN1(in2[11]), .IN2(in1[11]), .QN(n5) );
  NOR2X0 U15 ( .IN1(n5), .IN2(cout[11]), .QN(sumout[11]) );
  AND2X1 U16 ( .IN1(in2[12]), .IN2(in1[12]), .Q(cout[12]) );
  NOR2X0 U17 ( .IN1(in2[12]), .IN2(in1[12]), .QN(n6) );
  NOR2X0 U18 ( .IN1(n6), .IN2(cout[12]), .QN(sumout[12]) );
  AND2X1 U19 ( .IN1(in3[40]), .IN2(in2[40]), .Q(cout[40]) );
  NOR2X0 U20 ( .IN1(in3[40]), .IN2(in2[40]), .QN(n7) );
  NOR2X0 U21 ( .IN1(n7), .IN2(cout[40]), .QN(sumout[40]) );
  AND2X1 U22 ( .IN1(in3[41]), .IN2(in2[41]), .Q(cout[41]) );
  NOR2X0 U23 ( .IN1(in3[41]), .IN2(in2[41]), .QN(n8) );
  NOR2X0 U24 ( .IN1(n8), .IN2(cout[41]), .QN(sumout[41]) );
  AND2X1 U25 ( .IN1(in3[42]), .IN2(in2[42]), .Q(cout[42]) );
  NOR2X0 U26 ( .IN1(in3[42]), .IN2(in2[42]), .QN(n9) );
  NOR2X0 U27 ( .IN1(n9), .IN2(cout[42]), .QN(sumout[42]) );
  AND2X1 U28 ( .IN1(in3[43]), .IN2(in2[43]), .Q(cout[43]) );
  NOR2X0 U29 ( .IN1(in3[43]), .IN2(in2[43]), .QN(n10) );
  NOR2X0 U30 ( .IN1(n10), .IN2(cout[43]), .QN(sumout[43]) );
  AND2X1 U31 ( .IN1(in3[44]), .IN2(in2[44]), .Q(cout[44]) );
  NOR2X0 U32 ( .IN1(in3[44]), .IN2(in2[44]), .QN(n11) );
  NOR2X0 U33 ( .IN1(n11), .IN2(cout[44]), .QN(sumout[44]) );
  AND2X1 U34 ( .IN1(in3[45]), .IN2(in2[45]), .Q(cout[45]) );
  NOR2X0 U35 ( .IN1(in3[45]), .IN2(in2[45]), .QN(n12) );
  NOR2X0 U36 ( .IN1(n12), .IN2(cout[45]), .QN(sumout[45]) );
  AND2X1 U37 ( .IN1(in3[46]), .IN2(in2[46]), .Q(cout[46]) );
  NOR2X0 U38 ( .IN1(in3[46]), .IN2(in2[46]), .QN(n13) );
  NOR2X0 U39 ( .IN1(n13), .IN2(cout[46]), .QN(sumout[46]) );
  INVX0 U40 ( .INP(in3[47]), .ZN(sumout[47]) );
  AND2X1 U41 ( .IN1(in2[5]), .IN2(in1[5]), .Q(cout[5]) );
  AND2X1 U42 ( .IN1(in2[6]), .IN2(in1[6]), .Q(cout[6]) );
  NOR2X0 U43 ( .IN1(in2[6]), .IN2(in1[6]), .QN(n14) );
  NOR2X0 U44 ( .IN1(n14), .IN2(cout[6]), .QN(sumout[6]) );
  FADDX1 U45 ( .A(in1[13]), .B(in2[13]), .CI(in3[13]), .CO(cout[13]), .S(
        sumout[13]) );
  FADDX1 U46 ( .A(in1[14]), .B(in2[14]), .CI(in3[14]), .CO(cout[14]), .S(
        sumout[14]) );
  FADDX1 U47 ( .A(in1[15]), .B(in2[15]), .CI(in3[15]), .CO(cout[15]), .S(
        sumout[15]) );
  FADDX1 U48 ( .A(in1[16]), .B(in2[16]), .CI(in3[16]), .CO(cout[16]), .S(
        sumout[16]) );
  FADDX1 U49 ( .A(in1[17]), .B(in2[17]), .CI(in3[17]), .CO(cout[17]), .S(
        sumout[17]) );
  FADDX1 U50 ( .A(in1[18]), .B(in2[18]), .CI(in3[18]), .CO(cout[18]), .S(
        sumout[18]) );
  FADDX1 U51 ( .A(in1[19]), .B(in2[19]), .CI(in3[19]), .CO(cout[19]), .S(
        sumout[19]) );
  FADDX1 U52 ( .A(in1[20]), .B(in2[20]), .CI(in3[20]), .CO(cout[20]), .S(
        sumout[20]) );
  FADDX1 U53 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U54 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U55 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U56 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U57 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U58 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U59 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U60 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U61 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U62 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U63 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U64 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
  FADDX1 U65 ( .A(in1[33]), .B(in2[33]), .CI(in3[33]), .CO(cout[33]), .S(
        sumout[33]) );
  FADDX1 U66 ( .A(in1[34]), .B(in2[34]), .CI(in3[34]), .CO(cout[34]), .S(
        sumout[34]) );
  FADDX1 U67 ( .A(in1[35]), .B(in2[35]), .CI(in3[35]), .CO(cout[35]), .S(
        sumout[35]) );
  FADDX1 U68 ( .A(in1[36]), .B(in2[36]), .CI(in3[36]), .CO(cout[36]), .S(
        sumout[36]) );
  FADDX1 U69 ( .A(in1[37]), .B(in2[37]), .CI(in3[37]), .CO(cout[37]), .S(
        sumout[37]) );
  FADDX1 U70 ( .A(in1[38]), .B(in2[38]), .CI(in3[38]), .CO(cout[38]), .S(
        sumout[38]) );
  FADDX1 U71 ( .A(in1[39]), .B(in2[39]), .CI(in3[39]), .CO(cout[39]), .S(
        sumout[39]) );
endmodule


module csa51squ_28 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17;

  NBUFFX2 U1 ( .INP(in1[6]), .Z(sumout[6]) );
  NBUFFX2 U2 ( .INP(in1[7]), .Z(sumout[7]) );
  NBUFFX2 U3 ( .INP(in1[8]), .Z(sumout[8]) );
  NBUFFX2 U4 ( .INP(in1[9]), .Z(sumout[9]) );
  NBUFFX2 U5 ( .INP(in1[10]), .Z(sumout[10]) );
  NBUFFX2 U6 ( .INP(in1[11]), .Z(sumout[11]) );
  AND2X1 U7 ( .IN1(in3[13]), .IN2(in1[13]), .Q(cout[13]) );
  NOR2X0 U8 ( .IN1(in3[13]), .IN2(in1[13]), .QN(n7) );
  NOR2X0 U9 ( .IN1(n7), .IN2(cout[13]), .QN(sumout[13]) );
  AND2X1 U10 ( .IN1(in3[15]), .IN2(in1[15]), .Q(cout[15]) );
  NOR2X0 U11 ( .IN1(in3[15]), .IN2(in1[15]), .QN(n8) );
  NOR2X0 U12 ( .IN1(n8), .IN2(cout[15]), .QN(sumout[15]) );
  AND2X1 U13 ( .IN1(in3[17]), .IN2(in1[17]), .Q(cout[17]) );
  NOR2X0 U14 ( .IN1(in3[17]), .IN2(in1[17]), .QN(n9) );
  NOR2X0 U15 ( .IN1(n9), .IN2(cout[17]), .QN(sumout[17]) );
  AND2X1 U16 ( .IN1(in3[43]), .IN2(in2[43]), .Q(cout[43]) );
  NOR2X0 U17 ( .IN1(in3[43]), .IN2(in2[43]), .QN(n10) );
  NOR2X0 U18 ( .IN1(n10), .IN2(cout[43]), .QN(sumout[43]) );
  AND2X1 U19 ( .IN1(in3[44]), .IN2(in2[44]), .Q(cout[44]) );
  NOR2X0 U20 ( .IN1(in3[44]), .IN2(in2[44]), .QN(n11) );
  NOR2X0 U21 ( .IN1(n11), .IN2(cout[44]), .QN(sumout[44]) );
  AND2X1 U22 ( .IN1(in3[45]), .IN2(in2[45]), .Q(cout[45]) );
  NOR2X0 U23 ( .IN1(in3[45]), .IN2(in2[45]), .QN(n12) );
  NOR2X0 U24 ( .IN1(n12), .IN2(cout[45]), .QN(sumout[45]) );
  AND2X1 U25 ( .IN1(in3[46]), .IN2(in2[46]), .Q(cout[46]) );
  NOR2X0 U26 ( .IN1(in3[46]), .IN2(in2[46]), .QN(n13) );
  NOR2X0 U27 ( .IN1(n13), .IN2(cout[46]), .QN(sumout[46]) );
  XOR2X1 U28 ( .IN1(in3[47]), .IN2(in2[47]), .Q(sumout[47]) );
  AND2X1 U29 ( .IN1(in3[12]), .IN2(in1[12]), .Q(cout[12]) );
  NOR2X0 U30 ( .IN1(in3[12]), .IN2(in1[12]), .QN(n14) );
  NOR2X0 U31 ( .IN1(n14), .IN2(cout[12]), .QN(sumout[12]) );
  AND2X1 U32 ( .IN1(in3[14]), .IN2(in1[14]), .Q(cout[14]) );
  NOR2X0 U33 ( .IN1(in3[14]), .IN2(in1[14]), .QN(n15) );
  NOR2X0 U34 ( .IN1(n15), .IN2(cout[14]), .QN(sumout[14]) );
  AND2X1 U35 ( .IN1(in3[16]), .IN2(in1[16]), .Q(cout[16]) );
  NOR2X0 U36 ( .IN1(in3[16]), .IN2(in1[16]), .QN(n16) );
  NOR2X0 U37 ( .IN1(n16), .IN2(cout[16]), .QN(sumout[16]) );
  AND2X1 U38 ( .IN1(in3[18]), .IN2(in1[18]), .Q(cout[18]) );
  NOR2X0 U39 ( .IN1(in3[18]), .IN2(in1[18]), .QN(n17) );
  NOR2X0 U40 ( .IN1(n17), .IN2(cout[18]), .QN(sumout[18]) );
  FADDX1 U41 ( .A(in1[19]), .B(in2[19]), .CI(in3[19]), .CO(cout[19]), .S(
        sumout[19]) );
  FADDX1 U42 ( .A(in1[20]), .B(in2[20]), .CI(in3[20]), .CO(cout[20]), .S(
        sumout[20]) );
  FADDX1 U43 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U44 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U45 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U46 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U47 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U48 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U49 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U50 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U51 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U52 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U53 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U54 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
  FADDX1 U55 ( .A(in1[33]), .B(in2[33]), .CI(in3[33]), .CO(cout[33]), .S(
        sumout[33]) );
  FADDX1 U56 ( .A(in1[34]), .B(in2[34]), .CI(in3[34]), .CO(cout[34]), .S(
        sumout[34]) );
  FADDX1 U57 ( .A(in1[35]), .B(in2[35]), .CI(in3[35]), .CO(cout[35]), .S(
        sumout[35]) );
  FADDX1 U58 ( .A(in1[36]), .B(in2[36]), .CI(in3[36]), .CO(cout[36]), .S(
        sumout[36]) );
  FADDX1 U59 ( .A(in1[37]), .B(in2[37]), .CI(in3[37]), .CO(cout[37]), .S(
        sumout[37]) );
  FADDX1 U60 ( .A(in1[38]), .B(in2[38]), .CI(in3[38]), .CO(cout[38]), .S(
        sumout[38]) );
  FADDX1 U61 ( .A(in1[39]), .B(in2[39]), .CI(in3[39]), .CO(cout[39]), .S(
        sumout[39]) );
  FADDX1 U62 ( .A(in1[40]), .B(in2[40]), .CI(in3[40]), .CO(cout[40]), .S(
        sumout[40]) );
  FADDX1 U63 ( .A(in1[41]), .B(in2[41]), .CI(in3[41]), .CO(cout[41]), .S(
        sumout[41]) );
  FADDX1 U64 ( .A(in1[42]), .B(in2[42]), .CI(in3[42]), .CO(cout[42]), .S(
        sumout[42]) );
endmodule


module csa51squ_29 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19;

  NBUFFX2 U1 ( .INP(in2[46]), .Z(sumout[46]) );
  NBUFFX2 U2 ( .INP(in2[45]), .Z(sumout[45]) );
  NBUFFX2 U3 ( .INP(in2[44]), .Z(sumout[44]) );
  NBUFFX2 U4 ( .INP(in2[43]), .Z(sumout[43]) );
  NBUFFX2 U5 ( .INP(in2[42]), .Z(sumout[42]) );
  NBUFFX2 U6 ( .INP(in2[41]), .Z(sumout[41]) );
  NBUFFX2 U7 ( .INP(in2[40]), .Z(sumout[40]) );
  NBUFFX2 U8 ( .INP(in2[39]), .Z(sumout[39]) );
  AND2X1 U9 ( .IN1(in2[7]), .IN2(in1[7]), .Q(cout[7]) );
  NOR2X0 U10 ( .IN1(in2[7]), .IN2(in1[7]), .QN(n9) );
  NOR2X0 U11 ( .IN1(n9), .IN2(cout[7]), .QN(sumout[7]) );
  AND2X1 U12 ( .IN1(in2[8]), .IN2(in1[8]), .Q(cout[8]) );
  NOR2X0 U13 ( .IN1(in2[8]), .IN2(in1[8]), .QN(n10) );
  NOR2X0 U14 ( .IN1(n10), .IN2(cout[8]), .QN(sumout[8]) );
  AND2X1 U15 ( .IN1(in2[9]), .IN2(in1[9]), .Q(cout[9]) );
  NOR2X0 U16 ( .IN1(in2[9]), .IN2(in1[9]), .QN(n11) );
  NOR2X0 U17 ( .IN1(n11), .IN2(cout[9]), .QN(sumout[9]) );
  AND2X1 U18 ( .IN1(in3[33]), .IN2(in2[33]), .Q(cout[33]) );
  NOR2X0 U19 ( .IN1(in3[33]), .IN2(in2[33]), .QN(n12) );
  NOR2X0 U20 ( .IN1(n12), .IN2(cout[33]), .QN(sumout[33]) );
  AND2X1 U21 ( .IN1(in3[34]), .IN2(in2[34]), .Q(cout[34]) );
  NOR2X0 U22 ( .IN1(in3[34]), .IN2(in2[34]), .QN(n13) );
  NOR2X0 U23 ( .IN1(n13), .IN2(cout[34]), .QN(sumout[34]) );
  AND2X1 U24 ( .IN1(in3[35]), .IN2(in2[35]), .Q(cout[35]) );
  NOR2X0 U25 ( .IN1(in3[35]), .IN2(in2[35]), .QN(n14) );
  NOR2X0 U26 ( .IN1(n14), .IN2(cout[35]), .QN(sumout[35]) );
  AND2X1 U27 ( .IN1(in3[36]), .IN2(in2[36]), .Q(cout[36]) );
  NOR2X0 U28 ( .IN1(in3[36]), .IN2(in2[36]), .QN(n15) );
  NOR2X0 U29 ( .IN1(n15), .IN2(cout[36]), .QN(sumout[36]) );
  AND2X1 U30 ( .IN1(in3[37]), .IN2(in2[37]), .Q(cout[37]) );
  NOR2X0 U31 ( .IN1(in3[37]), .IN2(in2[37]), .QN(n16) );
  NOR2X0 U32 ( .IN1(n16), .IN2(cout[37]), .QN(sumout[37]) );
  AND2X1 U33 ( .IN1(in3[38]), .IN2(in2[38]), .Q(cout[38]) );
  NOR2X0 U34 ( .IN1(in3[38]), .IN2(in2[38]), .QN(n17) );
  NOR2X0 U35 ( .IN1(n17), .IN2(cout[38]), .QN(sumout[38]) );
  AND2X1 U36 ( .IN1(in2[4]), .IN2(in1[4]), .Q(cout[4]) );
  AND2X1 U37 ( .IN1(in2[5]), .IN2(in1[5]), .Q(cout[5]) );
  NOR2X0 U38 ( .IN1(in2[5]), .IN2(in1[5]), .QN(n18) );
  NOR2X0 U39 ( .IN1(n18), .IN2(cout[5]), .QN(sumout[5]) );
  AND2X1 U40 ( .IN1(in2[6]), .IN2(in1[6]), .Q(cout[6]) );
  NOR2X0 U41 ( .IN1(in2[6]), .IN2(in1[6]), .QN(n19) );
  NOR2X0 U42 ( .IN1(n19), .IN2(cout[6]), .QN(sumout[6]) );
  FADDX1 U43 ( .A(in1[10]), .B(in2[10]), .CI(in3[10]), .CO(cout[10]), .S(
        sumout[10]) );
  FADDX1 U44 ( .A(in1[11]), .B(in2[11]), .CI(in3[11]), .CO(cout[11]), .S(
        sumout[11]) );
  FADDX1 U45 ( .A(in1[12]), .B(in2[12]), .CI(in3[12]), .CO(cout[12]), .S(
        sumout[12]) );
  FADDX1 U46 ( .A(in1[13]), .B(in2[13]), .CI(in3[13]), .CO(cout[13]), .S(
        sumout[13]) );
  FADDX1 U47 ( .A(in1[14]), .B(in2[14]), .CI(in3[14]), .CO(cout[14]), .S(
        sumout[14]) );
  FADDX1 U48 ( .A(in1[15]), .B(in2[15]), .CI(in3[15]), .CO(cout[15]), .S(
        sumout[15]) );
  FADDX1 U49 ( .A(in1[16]), .B(in2[16]), .CI(in3[16]), .CO(cout[16]), .S(
        sumout[16]) );
  FADDX1 U50 ( .A(in1[17]), .B(in2[17]), .CI(in3[17]), .CO(cout[17]), .S(
        sumout[17]) );
  FADDX1 U51 ( .A(in1[18]), .B(in2[18]), .CI(in3[18]), .CO(cout[18]), .S(
        sumout[18]) );
  FADDX1 U52 ( .A(in1[19]), .B(in2[19]), .CI(in3[19]), .CO(cout[19]), .S(
        sumout[19]) );
  FADDX1 U53 ( .A(in1[20]), .B(in2[20]), .CI(in3[20]), .CO(cout[20]), .S(
        sumout[20]) );
  FADDX1 U54 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U55 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U56 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U57 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U58 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U59 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U60 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U61 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U62 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U63 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U64 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U65 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
endmodule


module csa51squ_30 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n7, n8, n9, n10, n11, n12, n13;

  NBUFFX2 U1 ( .INP(in1[12]), .Z(sumout[12]) );
  NBUFFX2 U2 ( .INP(in1[13]), .Z(sumout[13]) );
  NBUFFX2 U3 ( .INP(in1[14]), .Z(sumout[14]) );
  NBUFFX2 U4 ( .INP(in1[15]), .Z(sumout[15]) );
  NBUFFX2 U5 ( .INP(in1[16]), .Z(sumout[16]) );
  NBUFFX2 U6 ( .INP(in1[17]), .Z(sumout[17]) );
  AND2X1 U7 ( .IN1(in3[19]), .IN2(in1[19]), .Q(cout[19]) );
  NOR2X0 U8 ( .IN1(in3[19]), .IN2(in1[19]), .QN(n7) );
  NOR2X0 U9 ( .IN1(n7), .IN2(cout[19]), .QN(sumout[19]) );
  AND2X1 U10 ( .IN1(in3[44]), .IN2(in2[44]), .Q(cout[44]) );
  NOR2X0 U11 ( .IN1(in3[44]), .IN2(in2[44]), .QN(n8) );
  NOR2X0 U12 ( .IN1(n8), .IN2(cout[44]), .QN(sumout[44]) );
  AND2X1 U13 ( .IN1(in3[45]), .IN2(in2[45]), .Q(cout[45]) );
  NOR2X0 U14 ( .IN1(in3[45]), .IN2(in2[45]), .QN(n9) );
  NOR2X0 U15 ( .IN1(n9), .IN2(cout[45]), .QN(sumout[45]) );
  AND2X1 U16 ( .IN1(in3[46]), .IN2(in2[46]), .Q(cout[46]) );
  NOR2X0 U17 ( .IN1(in3[46]), .IN2(in2[46]), .QN(n10) );
  NOR2X0 U18 ( .IN1(n10), .IN2(cout[46]), .QN(sumout[46]) );
  XOR2X1 U19 ( .IN1(in3[47]), .IN2(in2[47]), .Q(sumout[47]) );
  AND2X1 U20 ( .IN1(in3[18]), .IN2(in1[18]), .Q(cout[18]) );
  NOR2X0 U21 ( .IN1(in3[18]), .IN2(in1[18]), .QN(n11) );
  NOR2X0 U22 ( .IN1(n11), .IN2(cout[18]), .QN(sumout[18]) );
  AND2X1 U23 ( .IN1(in3[20]), .IN2(in1[20]), .Q(cout[20]) );
  NOR2X0 U24 ( .IN1(in3[20]), .IN2(in1[20]), .QN(n12) );
  NOR2X0 U25 ( .IN1(n12), .IN2(cout[20]), .QN(sumout[20]) );
  INVX0 U26 ( .INP(in1[42]), .ZN(n13) );
  FADDX1 U27 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U28 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U29 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U30 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U31 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U32 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U33 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U34 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U35 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U36 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U37 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U38 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
  FADDX1 U39 ( .A(in1[33]), .B(in2[33]), .CI(in3[33]), .CO(cout[33]), .S(
        sumout[33]) );
  FADDX1 U40 ( .A(in1[34]), .B(in2[34]), .CI(in3[34]), .CO(cout[34]), .S(
        sumout[34]) );
  FADDX1 U41 ( .A(in1[35]), .B(in2[35]), .CI(in3[35]), .CO(cout[35]), .S(
        sumout[35]) );
  FADDX1 U42 ( .A(in1[36]), .B(in2[36]), .CI(in3[36]), .CO(cout[36]), .S(
        sumout[36]) );
  FADDX1 U43 ( .A(in1[37]), .B(in2[37]), .CI(in3[37]), .CO(cout[37]), .S(
        sumout[37]) );
  FADDX1 U44 ( .A(in1[38]), .B(in2[38]), .CI(in3[38]), .CO(cout[38]), .S(
        sumout[38]) );
  FADDX1 U45 ( .A(in1[39]), .B(in2[39]), .CI(in3[39]), .CO(cout[39]), .S(
        sumout[39]) );
  FADDX1 U46 ( .A(in1[40]), .B(in2[40]), .CI(in3[40]), .CO(cout[40]), .S(
        sumout[40]) );
  FADDX1 U47 ( .A(in1[41]), .B(in2[41]), .CI(in3[41]), .CO(cout[41]), .S(
        sumout[41]) );
  FADDX1 U48 ( .A(in1[42]), .B(in2[42]), .CI(in3[42]), .CO(cout[42]), .S(
        sumout[42]) );
  FADDX1 U49 ( .A(in2[43]), .B(in3[43]), .CI(n13), .CO(cout[43]), .S(
        sumout[43]) );
endmodule


module csa51squ_31 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n9, n10, n11, n12, n13, n14, n15;

  NBUFFX2 U1 ( .INP(in2[6]), .Z(sumout[6]) );
  NBUFFX2 U2 ( .INP(in2[7]), .Z(sumout[7]) );
  NBUFFX2 U3 ( .INP(in2[8]), .Z(sumout[8]) );
  NBUFFX2 U4 ( .INP(in3[42]), .Z(sumout[42]) );
  NBUFFX2 U5 ( .INP(in3[41]), .Z(sumout[41]) );
  NBUFFX2 U6 ( .INP(in3[39]), .Z(sumout[39]) );
  NBUFFX2 U7 ( .INP(in3[38]), .Z(sumout[38]) );
  NBUFFX2 U8 ( .INP(in3[40]), .Z(sumout[40]) );
  AND2X1 U9 ( .IN1(in2[13]), .IN2(in1[13]), .Q(cout[13]) );
  NOR2X0 U10 ( .IN1(in2[13]), .IN2(in1[13]), .QN(n9) );
  NOR2X0 U11 ( .IN1(n9), .IN2(cout[13]), .QN(sumout[13]) );
  AND2X1 U12 ( .IN1(in2[37]), .IN2(in3[37]), .Q(cout[37]) );
  INVX0 U13 ( .INP(in2[37]), .ZN(n15) );
  MUX21X1 U14 ( .IN1(in2[37]), .IN2(n15), .S(in3[37]), .Q(sumout[37]) );
  AND2X1 U15 ( .IN1(in2[9]), .IN2(in1[9]), .Q(cout[9]) );
  NOR2X0 U16 ( .IN1(in2[9]), .IN2(in1[9]), .QN(n10) );
  NOR2X0 U17 ( .IN1(n10), .IN2(cout[9]), .QN(sumout[9]) );
  AND2X1 U18 ( .IN1(in2[10]), .IN2(in1[10]), .Q(cout[10]) );
  NOR2X0 U19 ( .IN1(in2[10]), .IN2(in1[10]), .QN(n11) );
  NOR2X0 U20 ( .IN1(n11), .IN2(cout[10]), .QN(sumout[10]) );
  AND2X1 U21 ( .IN1(in2[11]), .IN2(in1[11]), .Q(cout[11]) );
  NOR2X0 U22 ( .IN1(in2[11]), .IN2(in1[11]), .QN(n12) );
  NOR2X0 U23 ( .IN1(n12), .IN2(cout[11]), .QN(sumout[11]) );
  AND2X1 U24 ( .IN1(in2[12]), .IN2(in1[12]), .Q(cout[12]) );
  NOR2X0 U25 ( .IN1(in2[12]), .IN2(in1[12]), .QN(n13) );
  NOR2X0 U26 ( .IN1(n13), .IN2(cout[12]), .QN(sumout[12]) );
  AND2X1 U27 ( .IN1(in2[14]), .IN2(in1[14]), .Q(cout[14]) );
  NOR2X0 U28 ( .IN1(in2[14]), .IN2(in1[14]), .QN(n14) );
  NOR2X0 U29 ( .IN1(n14), .IN2(cout[14]), .QN(sumout[14]) );
  FADDX1 U30 ( .A(in1[15]), .B(in2[15]), .CI(in3[15]), .CO(cout[15]), .S(
        sumout[15]) );
  FADDX1 U31 ( .A(in1[16]), .B(in2[16]), .CI(in3[16]), .CO(cout[16]), .S(
        sumout[16]) );
  FADDX1 U32 ( .A(in1[17]), .B(in2[17]), .CI(in3[17]), .CO(cout[17]), .S(
        sumout[17]) );
  FADDX1 U33 ( .A(in1[18]), .B(in2[18]), .CI(in3[18]), .CO(cout[18]), .S(
        sumout[18]) );
  FADDX1 U34 ( .A(in1[19]), .B(in2[19]), .CI(in3[19]), .CO(cout[19]), .S(
        sumout[19]) );
  FADDX1 U35 ( .A(in1[20]), .B(in2[20]), .CI(in3[20]), .CO(cout[20]), .S(
        sumout[20]) );
  FADDX1 U36 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U37 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U38 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U39 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U40 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U41 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U42 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U43 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U44 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U45 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U46 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U47 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
  FADDX1 U48 ( .A(in1[33]), .B(in2[33]), .CI(in3[33]), .CO(cout[33]), .S(
        sumout[33]) );
  FADDX1 U49 ( .A(in1[34]), .B(in2[34]), .CI(in3[34]), .CO(cout[34]), .S(
        sumout[34]) );
  FADDX1 U50 ( .A(in1[35]), .B(in2[35]), .CI(in3[35]), .CO(cout[35]), .S(
        sumout[35]) );
  FADDX1 U51 ( .A(in1[36]), .B(in3[36]), .CI(n15), .CO(cout[36]), .S(
        sumout[36]) );
endmodule


module csa51squ_32 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36;

  NBUFFX2 U1 ( .INP(in3[46]), .Z(sumout[46]) );
  NBUFFX2 U2 ( .INP(in3[45]), .Z(sumout[45]) );
  NBUFFX2 U3 ( .INP(in3[44]), .Z(sumout[44]) );
  NBUFFX2 U4 ( .INP(in3[43]), .Z(sumout[43]) );
  NBUFFX2 U5 ( .INP(in3[42]), .Z(sumout[42]) );
  NBUFFX2 U6 ( .INP(in3[33]), .Z(sumout[33]) );
  NBUFFX2 U7 ( .INP(in3[32]), .Z(sumout[32]) );
  NBUFFX2 U8 ( .INP(in3[37]), .Z(sumout[37]) );
  NBUFFX2 U9 ( .INP(in3[36]), .Z(sumout[36]) );
  NBUFFX2 U10 ( .INP(in3[35]), .Z(sumout[35]) );
  NBUFFX2 U11 ( .INP(in3[34]), .Z(sumout[34]) );
  NBUFFX2 U12 ( .INP(in3[41]), .Z(sumout[41]) );
  NBUFFX2 U13 ( .INP(in3[40]), .Z(sumout[40]) );
  NBUFFX2 U14 ( .INP(in3[39]), .Z(sumout[39]) );
  NBUFFX2 U15 ( .INP(in3[38]), .Z(sumout[38]) );
  AND2X1 U16 ( .IN1(in2[31]), .IN2(in3[31]), .Q(cout[31]) );
  INVX0 U17 ( .INP(in2[31]), .ZN(n36) );
  MUX21X1 U18 ( .IN1(in2[31]), .IN2(n36), .S(in3[31]), .Q(sumout[31]) );
  AND2X1 U19 ( .IN1(in2[3]), .IN2(in1[3]), .Q(cout[3]) );
  AND2X1 U20 ( .IN1(in2[4]), .IN2(in1[4]), .Q(cout[4]) );
  NOR2X0 U21 ( .IN1(in2[4]), .IN2(in1[4]), .QN(n16) );
  NOR2X0 U22 ( .IN1(n16), .IN2(cout[4]), .QN(sumout[4]) );
  AND2X1 U23 ( .IN1(in2[5]), .IN2(in1[5]), .Q(cout[5]) );
  NOR2X0 U24 ( .IN1(in2[5]), .IN2(in1[5]), .QN(n17) );
  NOR2X0 U25 ( .IN1(n17), .IN2(cout[5]), .QN(sumout[5]) );
  AND2X1 U26 ( .IN1(in2[6]), .IN2(in1[6]), .Q(cout[6]) );
  NOR2X0 U27 ( .IN1(in2[6]), .IN2(in1[6]), .QN(n18) );
  NOR2X0 U28 ( .IN1(n18), .IN2(cout[6]), .QN(sumout[6]) );
  AND2X1 U29 ( .IN1(in2[7]), .IN2(in1[7]), .Q(cout[7]) );
  NOR2X0 U30 ( .IN1(in2[7]), .IN2(in1[7]), .QN(n19) );
  NOR2X0 U31 ( .IN1(n19), .IN2(cout[7]), .QN(sumout[7]) );
  AND2X1 U32 ( .IN1(in2[8]), .IN2(in1[8]), .Q(cout[8]) );
  NOR2X0 U33 ( .IN1(in2[8]), .IN2(in1[8]), .QN(n20) );
  NOR2X0 U34 ( .IN1(n20), .IN2(cout[8]), .QN(sumout[8]) );
  AND2X1 U35 ( .IN1(in2[9]), .IN2(in1[9]), .Q(cout[9]) );
  NOR2X0 U36 ( .IN1(in2[9]), .IN2(in1[9]), .QN(n21) );
  NOR2X0 U37 ( .IN1(n21), .IN2(cout[9]), .QN(sumout[9]) );
  AND2X1 U38 ( .IN1(in2[10]), .IN2(in1[10]), .Q(cout[10]) );
  NOR2X0 U39 ( .IN1(in2[10]), .IN2(in1[10]), .QN(n22) );
  NOR2X0 U40 ( .IN1(n22), .IN2(cout[10]), .QN(sumout[10]) );
  AND2X1 U41 ( .IN1(in2[11]), .IN2(in1[11]), .Q(cout[11]) );
  NOR2X0 U42 ( .IN1(in2[11]), .IN2(in1[11]), .QN(n23) );
  NOR2X0 U43 ( .IN1(n23), .IN2(cout[11]), .QN(sumout[11]) );
  AND2X1 U44 ( .IN1(in2[12]), .IN2(in1[12]), .Q(cout[12]) );
  NOR2X0 U45 ( .IN1(in2[12]), .IN2(in1[12]), .QN(n24) );
  NOR2X0 U46 ( .IN1(n24), .IN2(cout[12]), .QN(sumout[12]) );
  AND2X1 U47 ( .IN1(in2[13]), .IN2(in1[13]), .Q(cout[13]) );
  NOR2X0 U48 ( .IN1(in2[13]), .IN2(in1[13]), .QN(n25) );
  NOR2X0 U49 ( .IN1(n25), .IN2(cout[13]), .QN(sumout[13]) );
  AND2X1 U50 ( .IN1(in2[14]), .IN2(in1[14]), .Q(cout[14]) );
  NOR2X0 U51 ( .IN1(in2[14]), .IN2(in1[14]), .QN(n26) );
  NOR2X0 U52 ( .IN1(n26), .IN2(cout[14]), .QN(sumout[14]) );
  AND2X1 U53 ( .IN1(in2[15]), .IN2(in1[15]), .Q(cout[15]) );
  NOR2X0 U54 ( .IN1(in2[15]), .IN2(in1[15]), .QN(n27) );
  NOR2X0 U55 ( .IN1(n27), .IN2(cout[15]), .QN(sumout[15]) );
  AND2X1 U56 ( .IN1(in2[16]), .IN2(in1[16]), .Q(cout[16]) );
  NOR2X0 U57 ( .IN1(in2[16]), .IN2(in1[16]), .QN(n28) );
  NOR2X0 U58 ( .IN1(n28), .IN2(cout[16]), .QN(sumout[16]) );
  AND2X1 U59 ( .IN1(in2[17]), .IN2(in1[17]), .Q(cout[17]) );
  NOR2X0 U60 ( .IN1(in2[17]), .IN2(in1[17]), .QN(n29) );
  NOR2X0 U61 ( .IN1(n29), .IN2(cout[17]), .QN(sumout[17]) );
  AND2X1 U62 ( .IN1(in2[18]), .IN2(in1[18]), .Q(cout[18]) );
  NOR2X0 U63 ( .IN1(in2[18]), .IN2(in1[18]), .QN(n30) );
  NOR2X0 U64 ( .IN1(n30), .IN2(cout[18]), .QN(sumout[18]) );
  AND2X1 U65 ( .IN1(in2[19]), .IN2(in1[19]), .Q(cout[19]) );
  NOR2X0 U66 ( .IN1(in2[19]), .IN2(in1[19]), .QN(n31) );
  NOR2X0 U67 ( .IN1(n31), .IN2(cout[19]), .QN(sumout[19]) );
  AND2X1 U68 ( .IN1(in2[20]), .IN2(in1[20]), .Q(cout[20]) );
  NOR2X0 U69 ( .IN1(in2[20]), .IN2(in1[20]), .QN(n32) );
  NOR2X0 U70 ( .IN1(n32), .IN2(cout[20]), .QN(sumout[20]) );
  AND2X1 U71 ( .IN1(in2[21]), .IN2(in1[21]), .Q(cout[21]) );
  NOR2X0 U72 ( .IN1(in2[21]), .IN2(in1[21]), .QN(n33) );
  NOR2X0 U73 ( .IN1(n33), .IN2(cout[21]), .QN(sumout[21]) );
  AND2X1 U74 ( .IN1(in2[22]), .IN2(in1[22]), .Q(cout[22]) );
  NOR2X0 U75 ( .IN1(in2[22]), .IN2(in1[22]), .QN(n34) );
  NOR2X0 U76 ( .IN1(n34), .IN2(cout[22]), .QN(sumout[22]) );
  AND2X1 U77 ( .IN1(in2[23]), .IN2(in1[23]), .Q(cout[23]) );
  NOR2X0 U78 ( .IN1(in2[23]), .IN2(in1[23]), .QN(n35) );
  NOR2X0 U79 ( .IN1(n35), .IN2(cout[23]), .QN(sumout[23]) );
  FADDX1 U80 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U81 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U82 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U83 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U84 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U85 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U86 ( .A(in1[30]), .B(in3[30]), .CI(n36), .CO(cout[30]), .S(
        sumout[30]) );
endmodule


module csa51squ_33 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n3, n4, n5, n6, n7;

  NBUFFX2 U1 ( .INP(in1[18]), .Z(sumout[18]) );
  NBUFFX2 U2 ( .INP(in1[19]), .Z(sumout[19]) );
  AND2X1 U3 ( .IN1(in2[20]), .IN2(in1[20]), .Q(cout[20]) );
  NOR2X0 U4 ( .IN1(in2[20]), .IN2(in1[20]), .QN(n3) );
  NOR2X0 U5 ( .IN1(n3), .IN2(cout[20]), .QN(sumout[20]) );
  AND2X1 U6 ( .IN1(in2[21]), .IN2(in1[21]), .Q(cout[21]) );
  NOR2X0 U7 ( .IN1(in2[21]), .IN2(in1[21]), .QN(n4) );
  NOR2X0 U8 ( .IN1(n4), .IN2(cout[21]), .QN(sumout[21]) );
  AND2X1 U9 ( .IN1(in2[46]), .IN2(in3[46]), .Q(cout[46]) );
  NOR2X0 U10 ( .IN1(in2[46]), .IN2(in3[46]), .QN(n5) );
  NOR2X0 U11 ( .IN1(n5), .IN2(cout[46]), .QN(sumout[46]) );
  INVX0 U12 ( .INP(in2[46]), .ZN(n6) );
  MUX21X1 U13 ( .IN1(n6), .IN2(in2[46]), .S(in3[47]), .Q(sumout[47]) );
  INVX0 U14 ( .INP(in1[44]), .ZN(n7) );
  FADDX1 U15 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U16 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U17 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U18 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U19 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U20 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U21 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U22 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U23 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U24 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U25 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
  FADDX1 U26 ( .A(in1[33]), .B(in2[33]), .CI(in3[33]), .CO(cout[33]), .S(
        sumout[33]) );
  FADDX1 U27 ( .A(in1[34]), .B(in2[34]), .CI(in3[34]), .CO(cout[34]), .S(
        sumout[34]) );
  FADDX1 U28 ( .A(in1[35]), .B(in2[35]), .CI(in3[35]), .CO(cout[35]), .S(
        sumout[35]) );
  FADDX1 U29 ( .A(in1[36]), .B(in2[36]), .CI(in3[36]), .CO(cout[36]), .S(
        sumout[36]) );
  FADDX1 U30 ( .A(in1[37]), .B(in2[37]), .CI(in3[37]), .CO(cout[37]), .S(
        sumout[37]) );
  FADDX1 U31 ( .A(in1[38]), .B(in2[38]), .CI(in3[38]), .CO(cout[38]), .S(
        sumout[38]) );
  FADDX1 U32 ( .A(in1[39]), .B(in2[39]), .CI(in3[39]), .CO(cout[39]), .S(
        sumout[39]) );
  FADDX1 U33 ( .A(in1[40]), .B(in2[40]), .CI(in3[40]), .CO(cout[40]), .S(
        sumout[40]) );
  FADDX1 U34 ( .A(in1[41]), .B(in2[41]), .CI(in3[41]), .CO(cout[41]), .S(
        sumout[41]) );
  FADDX1 U35 ( .A(in1[42]), .B(in2[42]), .CI(in3[42]), .CO(cout[42]), .S(
        sumout[42]) );
  FADDX1 U36 ( .A(in1[43]), .B(in2[43]), .CI(in3[43]), .CO(cout[43]), .S(
        sumout[43]) );
  FADDX1 U37 ( .A(in1[44]), .B(in2[44]), .CI(in3[44]), .CO(cout[44]), .S(
        sumout[44]) );
  FADDX1 U38 ( .A(in2[45]), .B(in3[45]), .CI(n7), .CO(cout[45]), .S(sumout[45]) );
endmodule


module csa51squ_34 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n5, n6, n7, n8, n9, n10;

  AND2X1 U1 ( .IN1(in3[37]), .IN2(in2[37]), .Q(cout[37]) );
  NAND2X0 U2 ( .IN1(n5), .IN2(cout[39]), .QN(sumout[39]) );
  NAND2X0 U3 ( .IN1(in2[39]), .IN2(in3[39]), .QN(n5) );
  NBUFFX2 U4 ( .INP(in1[12]), .Z(sumout[12]) );
  NBUFFX2 U5 ( .INP(in1[13]), .Z(sumout[13]) );
  NBUFFX2 U6 ( .INP(in3[42]), .Z(sumout[42]) );
  XOR2X1 U7 ( .IN1(in2[37]), .IN2(in3[37]), .Q(sumout[37]) );
  OR2X1 U8 ( .IN1(in3[39]), .IN2(in2[39]), .Q(cout[39]) );
  AND2X1 U9 ( .IN1(in3[38]), .IN2(in2[38]), .Q(cout[38]) );
  NOR2X0 U10 ( .IN1(in3[38]), .IN2(in2[38]), .QN(n6) );
  NOR2X0 U11 ( .IN1(n6), .IN2(cout[38]), .QN(sumout[38]) );
  AND2X1 U12 ( .IN1(in2[14]), .IN2(in1[14]), .Q(cout[14]) );
  NOR2X0 U13 ( .IN1(in2[14]), .IN2(in1[14]), .QN(n7) );
  NOR2X0 U14 ( .IN1(n7), .IN2(cout[14]), .QN(sumout[14]) );
  AND2X1 U15 ( .IN1(in2[15]), .IN2(in1[15]), .Q(cout[15]) );
  NOR2X0 U16 ( .IN1(in2[15]), .IN2(in1[15]), .QN(n8) );
  NOR2X0 U17 ( .IN1(n8), .IN2(cout[15]), .QN(sumout[15]) );
  AND2X1 U18 ( .IN1(in2[40]), .IN2(in3[40]), .Q(cout[40]) );
  NOR2X0 U19 ( .IN1(in2[40]), .IN2(in3[40]), .QN(n9) );
  NOR2X0 U20 ( .IN1(n9), .IN2(cout[40]), .QN(sumout[40]) );
  INVX0 U21 ( .INP(in3[41]), .ZN(n10) );
  NOR2X0 U22 ( .IN1(in2[40]), .IN2(n10), .QN(cout[41]) );
  MUX21X1 U23 ( .IN1(n10), .IN2(in3[41]), .S(in2[40]), .Q(sumout[41]) );
  FADDX1 U24 ( .A(in1[16]), .B(in2[16]), .CI(in3[16]), .CO(cout[16]), .S(
        sumout[16]) );
  FADDX1 U25 ( .A(in1[17]), .B(in2[17]), .CI(in3[17]), .CO(cout[17]), .S(
        sumout[17]) );
  FADDX1 U26 ( .A(in1[18]), .B(in2[18]), .CI(in3[18]), .CO(cout[18]), .S(
        sumout[18]) );
  FADDX1 U27 ( .A(in1[19]), .B(in2[19]), .CI(in3[19]), .CO(cout[19]), .S(
        sumout[19]) );
  FADDX1 U28 ( .A(in1[20]), .B(in2[20]), .CI(in3[20]), .CO(cout[20]), .S(
        sumout[20]) );
  FADDX1 U29 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U30 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U31 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U32 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U33 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U34 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U35 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U36 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U37 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U38 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U39 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U40 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
  FADDX1 U41 ( .A(in1[33]), .B(in2[33]), .CI(in3[33]), .CO(cout[33]), .S(
        sumout[33]) );
  FADDX1 U42 ( .A(in1[34]), .B(in2[34]), .CI(in3[34]), .CO(cout[34]), .S(
        sumout[34]) );
  FADDX1 U43 ( .A(in1[35]), .B(in2[35]), .CI(in3[35]), .CO(cout[35]), .S(
        sumout[35]) );
  FADDX1 U44 ( .A(in1[36]), .B(in2[36]), .CI(in3[36]), .CO(cout[36]), .S(
        sumout[36]) );
endmodule


module csa51squ_35 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n4, n5, n6, n7, n8;

  NBUFFX2 U1 ( .INP(in1[6]), .Z(sumout[6]) );
  NBUFFX2 U2 ( .INP(in1[7]), .Z(sumout[7]) );
  NBUFFX2 U3 ( .INP(in3[37]), .Z(sumout[37]) );
  AND2X1 U4 ( .IN1(in2[8]), .IN2(in1[8]), .Q(cout[8]) );
  NOR2X0 U5 ( .IN1(in2[8]), .IN2(in1[8]), .QN(n4) );
  NOR2X0 U6 ( .IN1(n4), .IN2(cout[8]), .QN(sumout[8]) );
  AND2X1 U7 ( .IN1(in2[9]), .IN2(in1[9]), .Q(cout[9]) );
  NOR2X0 U8 ( .IN1(in2[9]), .IN2(in1[9]), .QN(n5) );
  NOR2X0 U9 ( .IN1(n5), .IN2(cout[9]), .QN(sumout[9]) );
  AND2X1 U10 ( .IN1(in2[34]), .IN2(in3[34]), .Q(cout[34]) );
  NOR2X0 U11 ( .IN1(in2[34]), .IN2(in3[34]), .QN(n6) );
  NOR2X0 U12 ( .IN1(n6), .IN2(cout[34]), .QN(sumout[34]) );
  INVX0 U13 ( .INP(in3[35]), .ZN(n7) );
  NOR2X0 U14 ( .IN1(in2[34]), .IN2(n7), .QN(cout[35]) );
  MUX21X1 U15 ( .IN1(n7), .IN2(in3[35]), .S(in2[34]), .Q(sumout[35]) );
  INVX0 U16 ( .INP(in1[32]), .ZN(n8) );
  FADDX1 U17 ( .A(in1[10]), .B(in2[10]), .CI(in3[10]), .CO(cout[10]), .S(
        sumout[10]) );
  FADDX1 U18 ( .A(in1[11]), .B(in2[11]), .CI(in3[11]), .CO(cout[11]), .S(
        sumout[11]) );
  FADDX1 U19 ( .A(in1[12]), .B(in2[12]), .CI(in3[12]), .CO(cout[12]), .S(
        sumout[12]) );
  FADDX1 U20 ( .A(in1[13]), .B(in2[13]), .CI(in3[13]), .CO(cout[13]), .S(
        sumout[13]) );
  FADDX1 U21 ( .A(in1[14]), .B(in2[14]), .CI(in3[14]), .CO(cout[14]), .S(
        sumout[14]) );
  FADDX1 U22 ( .A(in1[15]), .B(in2[15]), .CI(in3[15]), .CO(cout[15]), .S(
        sumout[15]) );
  FADDX1 U23 ( .A(in1[16]), .B(in2[16]), .CI(in3[16]), .CO(cout[16]), .S(
        sumout[16]) );
  FADDX1 U24 ( .A(in1[17]), .B(in2[17]), .CI(in3[17]), .CO(cout[17]), .S(
        sumout[17]) );
  FADDX1 U25 ( .A(in1[18]), .B(in2[18]), .CI(in3[18]), .CO(cout[18]), .S(
        sumout[18]) );
  FADDX1 U26 ( .A(in1[19]), .B(in2[19]), .CI(in3[19]), .CO(cout[19]), .S(
        sumout[19]) );
  FADDX1 U27 ( .A(in1[20]), .B(in2[20]), .CI(in3[20]), .CO(cout[20]), .S(
        sumout[20]) );
  FADDX1 U28 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U29 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U30 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U31 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U32 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U33 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U34 ( .A(in1[27]), .B(in2[27]), .CI(in3[27]), .CO(cout[27]), .S(
        sumout[27]) );
  FADDX1 U35 ( .A(in1[28]), .B(in2[28]), .CI(in3[28]), .CO(cout[28]), .S(
        sumout[28]) );
  FADDX1 U36 ( .A(in1[29]), .B(in2[29]), .CI(in3[29]), .CO(cout[29]), .S(
        sumout[29]) );
  FADDX1 U37 ( .A(in1[30]), .B(in2[30]), .CI(in3[30]), .CO(cout[30]), .S(
        sumout[30]) );
  FADDX1 U38 ( .A(in1[31]), .B(in2[31]), .CI(in3[31]), .CO(cout[31]), .S(
        sumout[31]) );
  FADDX1 U39 ( .A(in1[32]), .B(in2[32]), .CI(in3[32]), .CO(cout[32]), .S(
        sumout[32]) );
  FADDX1 U40 ( .A(in2[33]), .B(in3[33]), .CI(n8), .CO(cout[33]), .S(sumout[33]) );
endmodule


module csa51squ_36 ( cout, sumout, in1, in2, in3 );
  output [50:0] cout;
  output [50:0] sumout;
  input [50:0] in1;
  input [50:0] in2;
  input [50:0] in3;
  wire   n2, n3, n4, n5;

  NBUFFX2 U1 ( .INP(in3[31]), .Z(sumout[31]) );
  AND2X1 U2 ( .IN1(in2[2]), .IN2(in1[2]), .Q(cout[2]) );
  AND2X1 U3 ( .IN1(in2[3]), .IN2(in1[3]), .Q(cout[3]) );
  NOR2X0 U4 ( .IN1(in2[3]), .IN2(in1[3]), .QN(n2) );
  NOR2X0 U5 ( .IN1(n2), .IN2(cout[3]), .QN(sumout[3]) );
  AND2X1 U6 ( .IN1(in2[28]), .IN2(in3[28]), .Q(cout[28]) );
  NOR2X0 U7 ( .IN1(in2[28]), .IN2(in3[28]), .QN(n3) );
  NOR2X0 U8 ( .IN1(n3), .IN2(cout[28]), .QN(sumout[28]) );
  INVX0 U9 ( .INP(in3[29]), .ZN(n4) );
  NOR2X0 U10 ( .IN1(in2[28]), .IN2(n4), .QN(cout[29]) );
  MUX21X1 U11 ( .IN1(n4), .IN2(in3[29]), .S(in2[28]), .Q(sumout[29]) );
  INVX0 U12 ( .INP(in1[26]), .ZN(n5) );
  FADDX1 U13 ( .A(in1[10]), .B(in2[10]), .CI(in3[10]), .CO(cout[10]), .S(
        sumout[10]) );
  FADDX1 U14 ( .A(in1[11]), .B(in2[11]), .CI(in3[11]), .CO(cout[11]), .S(
        sumout[11]) );
  FADDX1 U15 ( .A(in1[12]), .B(in2[12]), .CI(in3[12]), .CO(cout[12]), .S(
        sumout[12]) );
  FADDX1 U16 ( .A(in1[13]), .B(in2[13]), .CI(in3[13]), .CO(cout[13]), .S(
        sumout[13]) );
  FADDX1 U17 ( .A(in1[14]), .B(in2[14]), .CI(in3[14]), .CO(cout[14]), .S(
        sumout[14]) );
  FADDX1 U18 ( .A(in1[15]), .B(in2[15]), .CI(in3[15]), .CO(cout[15]), .S(
        sumout[15]) );
  FADDX1 U19 ( .A(in1[16]), .B(in2[16]), .CI(in3[16]), .CO(cout[16]), .S(
        sumout[16]) );
  FADDX1 U20 ( .A(in1[17]), .B(in2[17]), .CI(in3[17]), .CO(cout[17]), .S(
        sumout[17]) );
  FADDX1 U21 ( .A(in1[18]), .B(in2[18]), .CI(in3[18]), .CO(cout[18]), .S(
        sumout[18]) );
  FADDX1 U22 ( .A(in1[19]), .B(in2[19]), .CI(in3[19]), .CO(cout[19]), .S(
        sumout[19]) );
  FADDX1 U23 ( .A(in1[20]), .B(in2[20]), .CI(in3[20]), .CO(cout[20]), .S(
        sumout[20]) );
  FADDX1 U24 ( .A(in1[21]), .B(in2[21]), .CI(in3[21]), .CO(cout[21]), .S(
        sumout[21]) );
  FADDX1 U25 ( .A(in1[22]), .B(in2[22]), .CI(in3[22]), .CO(cout[22]), .S(
        sumout[22]) );
  FADDX1 U26 ( .A(in1[23]), .B(in2[23]), .CI(in3[23]), .CO(cout[23]), .S(
        sumout[23]) );
  FADDX1 U27 ( .A(in1[24]), .B(in2[24]), .CI(in3[24]), .CO(cout[24]), .S(
        sumout[24]) );
  FADDX1 U28 ( .A(in1[25]), .B(in2[25]), .CI(in3[25]), .CO(cout[25]), .S(
        sumout[25]) );
  FADDX1 U29 ( .A(in1[26]), .B(in2[26]), .CI(in3[26]), .CO(cout[26]), .S(
        sumout[26]) );
  FADDX1 U30 ( .A(in2[27]), .B(in3[27]), .CI(n5), .CO(cout[27]), .S(sumout[27]) );
  FADDX1 U31 ( .A(in1[4]), .B(in2[4]), .CI(in3[4]), .CO(cout[4]), .S(sumout[4]) );
  FADDX1 U32 ( .A(in1[5]), .B(in2[5]), .CI(in3[5]), .CO(cout[5]), .S(sumout[5]) );
  FADDX1 U33 ( .A(in1[6]), .B(in2[6]), .CI(in3[6]), .CO(cout[6]), .S(sumout[6]) );
  FADDX1 U34 ( .A(in1[7]), .B(in2[7]), .CI(in3[7]), .CO(cout[7]), .S(sumout[7]) );
  FADDX1 U35 ( .A(in1[8]), .B(in2[8]), .CI(in3[8]), .CO(cout[8]), .S(sumout[8]) );
  FADDX1 U36 ( .A(in1[9]), .B(in2[9]), .CI(in3[9]), .CO(cout[9]), .S(sumout[9]) );
endmodule


module booth27_27 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;


  NBUFFX2 U3 ( .INP(in2[22]), .Z(out1[22]) );
  NBUFFX2 U4 ( .INP(in2[21]), .Z(out1[21]) );
  NBUFFX2 U5 ( .INP(in2[20]), .Z(out1[20]) );
  NBUFFX2 U6 ( .INP(in2[0]), .Z(out1[0]) );
  NBUFFX2 U7 ( .INP(in2[19]), .Z(out1[19]) );
  NBUFFX2 U8 ( .INP(in2[18]), .Z(out1[18]) );
  NBUFFX2 U9 ( .INP(in2[6]), .Z(out1[6]) );
  NBUFFX2 U10 ( .INP(in2[5]), .Z(out1[5]) );
  NBUFFX2 U11 ( .INP(in2[4]), .Z(out1[4]) );
  NBUFFX2 U12 ( .INP(in2[3]), .Z(out1[3]) );
  NBUFFX2 U13 ( .INP(in2[2]), .Z(out1[2]) );
  NBUFFX2 U14 ( .INP(in2[1]), .Z(out1[1]) );
  NBUFFX2 U15 ( .INP(in2[9]), .Z(out1[9]) );
  NBUFFX2 U16 ( .INP(in2[8]), .Z(out1[8]) );
  NBUFFX2 U17 ( .INP(in2[7]), .Z(out1[7]) );
  NBUFFX2 U18 ( .INP(in2[13]), .Z(out1[13]) );
  NBUFFX2 U19 ( .INP(in2[12]), .Z(out1[12]) );
  NBUFFX2 U20 ( .INP(in2[11]), .Z(out1[11]) );
  NBUFFX2 U21 ( .INP(in2[10]), .Z(out1[10]) );
  NBUFFX2 U22 ( .INP(in2[17]), .Z(out1[17]) );
  NBUFFX2 U23 ( .INP(in2[16]), .Z(out1[16]) );
  NBUFFX2 U24 ( .INP(in2[15]), .Z(out1[15]) );
  NBUFFX2 U25 ( .INP(in2[14]), .Z(out1[14]) );
endmodule


module booth27_28 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76;

  NAND2X0 U3 ( .IN1(n1), .IN2(n2), .QN(n8) );
  NAND2X0 U4 ( .IN1(n71), .IN2(in2[0]), .QN(n15) );
  NAND2X0 U5 ( .IN1(n16), .IN2(in2[4]), .QN(n17) );
  NAND2X0 U6 ( .IN1(n22), .IN2(in2[6]), .QN(n23) );
  NAND2X0 U7 ( .IN1(n28), .IN2(in2[8]), .QN(n29) );
  NAND2X0 U8 ( .IN1(n31), .IN2(in2[9]), .QN(n32) );
  NAND2X0 U9 ( .IN1(n34), .IN2(in2[10]), .QN(n35) );
  NAND2X0 U10 ( .IN1(n37), .IN2(in2[11]), .QN(n38) );
  NAND2X0 U11 ( .IN1(n40), .IN2(in2[12]), .QN(n41) );
  NAND2X0 U12 ( .IN1(n49), .IN2(in2[15]), .QN(n50) );
  NAND2X0 U13 ( .IN1(n7), .IN2(n15), .QN(out1[1]) );
  NAND2X0 U14 ( .IN1(n10), .IN2(n9), .QN(out1[2]) );
  NAND2X0 U15 ( .IN1(n58), .IN2(in2[18]), .QN(n59) );
  NAND2X0 U16 ( .IN1(in1[1]), .IN2(in1[0]), .QN(out1[25]) );
  NOR2X0 U17 ( .IN1(in1[1]), .IN2(in1[0]), .QN(n71) );
  INVX0 U18 ( .INP(in2[0]), .ZN(n1) );
  INVX0 U19 ( .INP(in2[1]), .ZN(n2) );
  INVX0 U20 ( .INP(in2[3]), .ZN(n3) );
  INVX0 U21 ( .INP(in2[21]), .ZN(n4) );
  INVX0 U22 ( .INP(in2[22]), .ZN(n5) );
  INVX0 U23 ( .INP(in1[1]), .ZN(n6) );
  MUX21X1 U24 ( .IN1(in1[1]), .IN2(n6), .S(in1[0]), .Q(n74) );
  INVX0 U25 ( .INP(n74), .ZN(n76) );
  AO221X1 U26 ( .IN1(in2[0]), .IN2(in2[1]), .IN3(n1), .IN4(n2), .IN5(n76), .Q(
        n7) );
  MUX21X1 U27 ( .IN1(n2), .IN2(n8), .S(in2[2]), .Q(n12) );
  AO221X1 U28 ( .IN1(n12), .IN2(in2[2]), .IN3(n12), .IN4(n1), .IN5(n76), .Q(
        n10) );
  INVX0 U29 ( .INP(n71), .ZN(n13) );
  AO221X1 U30 ( .IN1(in2[0]), .IN2(in2[1]), .IN3(n1), .IN4(n2), .IN5(n13), .Q(
        n9) );
  NOR3X0 U31 ( .IN1(in2[0]), .IN2(in2[2]), .IN3(in2[1]), .QN(n11) );
  OR4X1 U32 ( .IN1(in2[3]), .IN2(in2[0]), .IN3(in2[2]), .IN4(in2[1]), .Q(n16)
         );
  OA21X1 U33 ( .IN1(n11), .IN2(n3), .IN3(n16), .Q(n18) );
  INVX0 U34 ( .INP(n18), .ZN(n14) );
  OAI222X1 U35 ( .IN1(n15), .IN2(in2[2]), .IN3(n14), .IN4(n76), .IN5(n13), 
        .IN6(n12), .QN(out1[3]) );
  OR2X1 U36 ( .IN1(in2[4]), .IN2(n16), .Q(n19) );
  AND2X1 U37 ( .IN1(n19), .IN2(n17), .Q(n21) );
  AO22X1 U38 ( .IN1(n71), .IN2(n18), .IN3(n21), .IN4(n74), .Q(out1[4]) );
  OR2X1 U39 ( .IN1(in2[5]), .IN2(n19), .Q(n22) );
  NAND2X0 U40 ( .IN1(n19), .IN2(in2[5]), .QN(n20) );
  AND2X1 U41 ( .IN1(n22), .IN2(n20), .Q(n24) );
  AO22X1 U42 ( .IN1(n71), .IN2(n21), .IN3(n24), .IN4(n74), .Q(out1[5]) );
  OR2X1 U43 ( .IN1(in2[6]), .IN2(n22), .Q(n25) );
  AND2X1 U44 ( .IN1(n25), .IN2(n23), .Q(n27) );
  AO22X1 U45 ( .IN1(n71), .IN2(n24), .IN3(n27), .IN4(n74), .Q(out1[6]) );
  OR2X1 U46 ( .IN1(in2[7]), .IN2(n25), .Q(n28) );
  NAND2X0 U47 ( .IN1(n25), .IN2(in2[7]), .QN(n26) );
  AND2X1 U48 ( .IN1(n28), .IN2(n26), .Q(n30) );
  AO22X1 U49 ( .IN1(n71), .IN2(n27), .IN3(n30), .IN4(n74), .Q(out1[7]) );
  OR2X1 U50 ( .IN1(in2[8]), .IN2(n28), .Q(n31) );
  AND2X1 U51 ( .IN1(n31), .IN2(n29), .Q(n33) );
  AO22X1 U52 ( .IN1(n71), .IN2(n30), .IN3(n33), .IN4(n74), .Q(out1[8]) );
  OR2X1 U53 ( .IN1(in2[9]), .IN2(n31), .Q(n34) );
  AND2X1 U54 ( .IN1(n34), .IN2(n32), .Q(n36) );
  AO22X1 U55 ( .IN1(n71), .IN2(n33), .IN3(n36), .IN4(n74), .Q(out1[9]) );
  OR2X1 U56 ( .IN1(in2[10]), .IN2(n34), .Q(n37) );
  AND2X1 U57 ( .IN1(n37), .IN2(n35), .Q(n39) );
  AO22X1 U58 ( .IN1(n71), .IN2(n36), .IN3(n39), .IN4(n74), .Q(out1[10]) );
  OR2X1 U59 ( .IN1(in2[11]), .IN2(n37), .Q(n40) );
  AND2X1 U60 ( .IN1(n40), .IN2(n38), .Q(n42) );
  AO22X1 U61 ( .IN1(n71), .IN2(n39), .IN3(n42), .IN4(n74), .Q(out1[11]) );
  OR2X1 U62 ( .IN1(in2[12]), .IN2(n40), .Q(n43) );
  AND2X1 U63 ( .IN1(n43), .IN2(n41), .Q(n45) );
  AO22X1 U64 ( .IN1(n71), .IN2(n42), .IN3(n45), .IN4(n74), .Q(out1[12]) );
  OR2X1 U65 ( .IN1(in2[13]), .IN2(n43), .Q(n46) );
  NAND2X0 U66 ( .IN1(n43), .IN2(in2[13]), .QN(n44) );
  AND2X1 U67 ( .IN1(n46), .IN2(n44), .Q(n48) );
  AO22X1 U68 ( .IN1(n71), .IN2(n45), .IN3(n48), .IN4(n74), .Q(out1[13]) );
  OR2X1 U69 ( .IN1(in2[14]), .IN2(n46), .Q(n49) );
  NAND2X0 U70 ( .IN1(n46), .IN2(in2[14]), .QN(n47) );
  AND2X1 U71 ( .IN1(n49), .IN2(n47), .Q(n51) );
  AO22X1 U72 ( .IN1(n71), .IN2(n48), .IN3(n51), .IN4(n74), .Q(out1[14]) );
  OR2X1 U73 ( .IN1(in2[15]), .IN2(n49), .Q(n52) );
  AND2X1 U74 ( .IN1(n52), .IN2(n50), .Q(n54) );
  AO22X1 U75 ( .IN1(n71), .IN2(n51), .IN3(n54), .IN4(n74), .Q(out1[15]) );
  OR2X1 U76 ( .IN1(in2[16]), .IN2(n52), .Q(n55) );
  NAND2X0 U77 ( .IN1(n52), .IN2(in2[16]), .QN(n53) );
  AND2X1 U78 ( .IN1(n55), .IN2(n53), .Q(n57) );
  AO22X1 U79 ( .IN1(n71), .IN2(n54), .IN3(n57), .IN4(n74), .Q(out1[16]) );
  OR2X1 U80 ( .IN1(in2[17]), .IN2(n55), .Q(n58) );
  NAND2X0 U81 ( .IN1(n55), .IN2(in2[17]), .QN(n56) );
  AND2X1 U82 ( .IN1(n58), .IN2(n56), .Q(n60) );
  AO22X1 U83 ( .IN1(n71), .IN2(n57), .IN3(n60), .IN4(n74), .Q(out1[17]) );
  OR2X1 U84 ( .IN1(in2[18]), .IN2(n58), .Q(n61) );
  AND2X1 U85 ( .IN1(n61), .IN2(n59), .Q(n63) );
  AO22X1 U86 ( .IN1(n71), .IN2(n60), .IN3(n63), .IN4(n74), .Q(out1[18]) );
  OR2X1 U87 ( .IN1(in2[19]), .IN2(n61), .Q(n64) );
  NAND2X0 U88 ( .IN1(n61), .IN2(in2[19]), .QN(n62) );
  AND2X1 U89 ( .IN1(n64), .IN2(n62), .Q(n65) );
  AO22X1 U90 ( .IN1(n71), .IN2(n63), .IN3(n65), .IN4(n74), .Q(out1[19]) );
  NOR2X0 U91 ( .IN1(in2[20]), .IN2(n64), .QN(n72) );
  AOI21X1 U92 ( .IN1(in2[20]), .IN2(n64), .IN3(n72), .QN(n66) );
  AO22X1 U93 ( .IN1(n71), .IN2(n65), .IN3(n66), .IN4(n74), .Q(out1[20]) );
  MUX21X1 U94 ( .IN1(n4), .IN2(in2[21]), .S(n72), .Q(n69) );
  AO22X1 U95 ( .IN1(n71), .IN2(n66), .IN3(n69), .IN4(n74), .Q(out1[21]) );
  INVX0 U96 ( .INP(n72), .ZN(n67) );
  NOR2X0 U97 ( .IN1(in2[21]), .IN2(n67), .QN(n70) );
  MUX21X1 U98 ( .IN1(n5), .IN2(in2[22]), .S(n70), .Q(n68) );
  AO22X1 U99 ( .IN1(n71), .IN2(n69), .IN3(n68), .IN4(n74), .Q(out1[22]) );
  MUX21X1 U100 ( .IN1(n71), .IN2(n74), .S(n70), .Q(n73) );
  AND3X1 U101 ( .IN1(n72), .IN2(n71), .IN3(n4), .Q(n75) );
  MUX21X1 U102 ( .IN1(n73), .IN2(n75), .S(in2[22]), .Q(out1[23]) );
  AO21X1 U103 ( .IN1(n75), .IN2(n5), .IN3(n74), .Q(out1[24]) );
  NOR2X0 U104 ( .IN1(n76), .IN2(n1), .QN(out1[0]) );
endmodule


module booth27_29 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n25), .IN2(n6), .QN(n30) );
  NAND2X0 U4 ( .IN1(n33), .IN2(n7), .QN(n37) );
  NAND2X0 U5 ( .IN1(n41), .IN2(n8), .QN(n45) );
  NAND2X0 U6 ( .IN1(n49), .IN2(n9), .QN(n53) );
  NAND2X0 U7 ( .IN1(n57), .IN2(n10), .QN(n61) );
  NAND2X0 U8 ( .IN1(n65), .IN2(n11), .QN(n77) );
  NAND2X0 U9 ( .IN1(n81), .IN2(n13), .QN(n89) );
  NAND2X0 U10 ( .IN1(n93), .IN2(n15), .QN(n101) );
  NAND2X0 U11 ( .IN1(n105), .IN2(n17), .QN(n114) );
  NAND2X0 U12 ( .IN1(n27), .IN2(n132), .QN(n4) );
  NAND2X0 U13 ( .IN1(in1[2]), .IN2(n77), .QN(n71) );
  NAND2X0 U14 ( .IN1(n70), .IN2(n132), .QN(n74) );
  NAND2X0 U15 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U16 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U17 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U18 ( .IN1(n118), .IN2(n19), .QN(n125) );
  NAND2X0 U19 ( .IN1(n141), .IN2(n130), .QN(n24) );
  NAND2X0 U20 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NAND2X0 U21 ( .IN1(n32), .IN2(n31), .QN(out1[3]) );
  NAND2X0 U22 ( .IN1(n36), .IN2(n35), .QN(out1[4]) );
  NAND2X0 U23 ( .IN1(n40), .IN2(n39), .QN(out1[5]) );
  NAND2X0 U24 ( .IN1(n44), .IN2(n43), .QN(out1[6]) );
  NAND2X0 U25 ( .IN1(n48), .IN2(n47), .QN(out1[7]) );
  NAND2X0 U26 ( .IN1(n52), .IN2(n51), .QN(out1[8]) );
  NAND2X0 U27 ( .IN1(n56), .IN2(n55), .QN(out1[9]) );
  NAND2X0 U28 ( .IN1(n60), .IN2(n59), .QN(out1[10]) );
  NAND2X0 U29 ( .IN1(n64), .IN2(n63), .QN(out1[11]) );
  NAND2X0 U30 ( .IN1(n69), .IN2(n68), .QN(out1[12]) );
  NAND2X0 U31 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U32 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U33 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U34 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U35 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U36 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U37 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U38 ( .IN1(n23), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U39 ( .IN1(in1[2]), .IN2(n22), .QN(n23) );
  NOR2X0 U40 ( .IN1(n28), .IN2(n26), .QN(n3) );
  NOR2X0 U41 ( .IN1(n142), .IN2(n21), .QN(n1) );
  NOR2X0 U42 ( .IN1(n142), .IN2(n111), .QN(n138) );
  INVX0 U43 ( .INP(n130), .ZN(n137) );
  INVX0 U44 ( .INP(n132), .ZN(n141) );
  NOR3X0 U45 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  NAND3X0 U46 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  MUX21X1 U47 ( .IN1(n22), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  INVX0 U48 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U49 ( .INP(in2[2]), .ZN(n6) );
  INVX0 U50 ( .INP(in2[4]), .ZN(n7) );
  INVX0 U51 ( .INP(in2[6]), .ZN(n8) );
  INVX0 U52 ( .INP(in2[8]), .ZN(n9) );
  INVX0 U53 ( .INP(in2[10]), .ZN(n10) );
  INVX0 U54 ( .INP(in2[12]), .ZN(n11) );
  INVX0 U55 ( .INP(in2[13]), .ZN(n12) );
  INVX0 U56 ( .INP(in2[14]), .ZN(n13) );
  INVX0 U57 ( .INP(in2[15]), .ZN(n14) );
  INVX0 U58 ( .INP(in2[16]), .ZN(n15) );
  INVX0 U59 ( .INP(in2[17]), .ZN(n16) );
  INVX0 U60 ( .INP(in2[18]), .ZN(n17) );
  INVX0 U61 ( .INP(in2[19]), .ZN(n18) );
  INVX0 U62 ( .INP(in2[20]), .ZN(n19) );
  INVX0 U63 ( .INP(in2[21]), .ZN(n20) );
  INVX0 U64 ( .INP(in2[22]), .ZN(n21) );
  INVX0 U65 ( .INP(in1[1]), .ZN(n22) );
  INVX0 U66 ( .INP(in1[2]), .ZN(n111) );
  INVX0 U67 ( .INP(n138), .ZN(n140) );
  NOR2X0 U68 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n25) );
  AOI21X1 U69 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n25), .QN(n27) );
  NOR2X0 U70 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U71 ( .IN1(n24), .IN2(in2[0]), .IN3(n138), .IN4(n27), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U72 ( .INP(n133), .ZN(n67) );
  NOR2X0 U73 ( .IN1(n67), .IN2(n6), .QN(n28) );
  OA21X1 U74 ( .IN1(n25), .IN2(n6), .IN3(n30), .Q(n29) );
  AO22X1 U75 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n29), .Q(n26) );
  AOI22X1 U76 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n29), .QN(n32) );
  NOR2X0 U77 ( .IN1(in2[3]), .IN2(n30), .QN(n33) );
  AO21X1 U78 ( .IN1(in2[3]), .IN2(n30), .IN3(n33), .Q(n34) );
  OA22X1 U79 ( .IN1(n6), .IN2(n130), .IN3(n140), .IN4(n34), .Q(n31) );
  OA21X1 U80 ( .IN1(n33), .IN2(n7), .IN3(n37), .Q(n38) );
  AOI22X1 U81 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n38), .QN(n36) );
  OA22X1 U82 ( .IN1(n67), .IN2(n7), .IN3(n141), .IN4(n34), .Q(n35) );
  NOR2X0 U83 ( .IN1(in2[5]), .IN2(n37), .QN(n41) );
  AO21X1 U84 ( .IN1(in2[5]), .IN2(n37), .IN3(n41), .Q(n42) );
  OA22X1 U85 ( .IN1(n7), .IN2(n130), .IN3(n140), .IN4(n42), .Q(n40) );
  AOI22X1 U86 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n38), .QN(n39) );
  OA21X1 U87 ( .IN1(n41), .IN2(n8), .IN3(n45), .Q(n46) );
  AOI22X1 U88 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n46), .QN(n44) );
  OA22X1 U89 ( .IN1(n67), .IN2(n8), .IN3(n141), .IN4(n42), .Q(n43) );
  NOR2X0 U90 ( .IN1(in2[7]), .IN2(n45), .QN(n49) );
  AO21X1 U91 ( .IN1(in2[7]), .IN2(n45), .IN3(n49), .Q(n50) );
  OA22X1 U92 ( .IN1(n8), .IN2(n130), .IN3(n140), .IN4(n50), .Q(n48) );
  AOI22X1 U93 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n46), .QN(n47) );
  OA21X1 U94 ( .IN1(n49), .IN2(n9), .IN3(n53), .Q(n54) );
  AOI22X1 U95 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n54), .QN(n52) );
  OA22X1 U96 ( .IN1(n67), .IN2(n9), .IN3(n141), .IN4(n50), .Q(n51) );
  NOR2X0 U97 ( .IN1(in2[9]), .IN2(n53), .QN(n57) );
  AO21X1 U98 ( .IN1(in2[9]), .IN2(n53), .IN3(n57), .Q(n58) );
  OA22X1 U99 ( .IN1(n9), .IN2(n130), .IN3(n140), .IN4(n58), .Q(n56) );
  AOI22X1 U100 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n54), .QN(n55) );
  OA21X1 U101 ( .IN1(n57), .IN2(n10), .IN3(n61), .Q(n62) );
  AOI22X1 U102 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n62), .QN(n60) );
  OA22X1 U103 ( .IN1(n67), .IN2(n10), .IN3(n141), .IN4(n58), .Q(n59) );
  NOR2X0 U104 ( .IN1(in2[11]), .IN2(n61), .QN(n65) );
  AO21X1 U105 ( .IN1(in2[11]), .IN2(n61), .IN3(n65), .Q(n66) );
  OA22X1 U106 ( .IN1(n10), .IN2(n130), .IN3(n140), .IN4(n66), .Q(n64) );
  AOI22X1 U107 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n62), .QN(n63) );
  OA21X1 U108 ( .IN1(n65), .IN2(n11), .IN3(n77), .Q(n70) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n70), .QN(n69) );
  OA22X1 U110 ( .IN1(n67), .IN2(n11), .IN3(n141), .IN4(n66), .Q(n68) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n12), .S(n71), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n11), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n13), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n12), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n12), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n14), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n13), .IN4(n85), .IN5(n84), 
        .Q(out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n15), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n14), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n14), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n16), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n15), .IN4(n97), .IN5(n96), 
        .Q(out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n17), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n16), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n16), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n18), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n17), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n19), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n18), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n18), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n20), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n19), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n21), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n20), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n20), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n21), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_30 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n33), .IN2(n7), .QN(n37) );
  NAND2X0 U4 ( .IN1(n41), .IN2(n8), .QN(n45) );
  NAND2X0 U5 ( .IN1(n49), .IN2(n9), .QN(n53) );
  NAND2X0 U6 ( .IN1(n57), .IN2(n10), .QN(n61) );
  NAND2X0 U7 ( .IN1(n25), .IN2(n6), .QN(n30) );
  NAND2X0 U8 ( .IN1(n65), .IN2(n11), .QN(n77) );
  NAND2X0 U9 ( .IN1(n81), .IN2(n13), .QN(n89) );
  NAND2X0 U10 ( .IN1(n93), .IN2(n15), .QN(n101) );
  NAND2X0 U11 ( .IN1(n105), .IN2(n17), .QN(n114) );
  NAND2X0 U12 ( .IN1(n118), .IN2(n19), .QN(n125) );
  NAND2X0 U13 ( .IN1(in1[2]), .IN2(n77), .QN(n71) );
  NAND2X0 U14 ( .IN1(n70), .IN2(n132), .QN(n74) );
  NAND2X0 U15 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U16 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U17 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U18 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U19 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U20 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U21 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U22 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NAND2X0 U23 ( .IN1(n27), .IN2(n132), .QN(n4) );
  NAND2X0 U24 ( .IN1(n32), .IN2(n31), .QN(out1[3]) );
  NAND2X0 U25 ( .IN1(n36), .IN2(n35), .QN(out1[4]) );
  NAND2X0 U26 ( .IN1(n40), .IN2(n39), .QN(out1[5]) );
  NAND2X0 U27 ( .IN1(n44), .IN2(n43), .QN(out1[6]) );
  NAND2X0 U28 ( .IN1(n48), .IN2(n47), .QN(out1[7]) );
  NAND2X0 U29 ( .IN1(n52), .IN2(n51), .QN(out1[8]) );
  NAND2X0 U30 ( .IN1(n56), .IN2(n55), .QN(out1[9]) );
  NAND2X0 U31 ( .IN1(n60), .IN2(n59), .QN(out1[10]) );
  NAND2X0 U32 ( .IN1(n64), .IN2(n63), .QN(out1[11]) );
  NAND2X0 U33 ( .IN1(n69), .IN2(n68), .QN(out1[12]) );
  NAND2X0 U34 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U35 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U36 ( .IN1(n141), .IN2(n130), .QN(n24) );
  NAND2X0 U37 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U38 ( .IN1(n23), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U39 ( .IN1(in1[2]), .IN2(n22), .QN(n23) );
  NOR2X0 U40 ( .IN1(n28), .IN2(n26), .QN(n3) );
  NOR2X0 U41 ( .IN1(n142), .IN2(n111), .QN(n138) );
  NOR2X0 U42 ( .IN1(n142), .IN2(n21), .QN(n1) );
  INVX0 U43 ( .INP(n130), .ZN(n137) );
  INVX0 U44 ( .INP(n132), .ZN(n141) );
  NOR3X0 U45 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  NAND3X0 U46 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  MUX21X1 U47 ( .IN1(n22), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  INVX0 U48 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U49 ( .INP(in2[2]), .ZN(n6) );
  INVX0 U50 ( .INP(in2[4]), .ZN(n7) );
  INVX0 U51 ( .INP(in2[6]), .ZN(n8) );
  INVX0 U52 ( .INP(in2[8]), .ZN(n9) );
  INVX0 U53 ( .INP(in2[10]), .ZN(n10) );
  INVX0 U54 ( .INP(in2[12]), .ZN(n11) );
  INVX0 U55 ( .INP(in2[13]), .ZN(n12) );
  INVX0 U56 ( .INP(in2[14]), .ZN(n13) );
  INVX0 U57 ( .INP(in2[15]), .ZN(n14) );
  INVX0 U58 ( .INP(in2[16]), .ZN(n15) );
  INVX0 U59 ( .INP(in2[17]), .ZN(n16) );
  INVX0 U60 ( .INP(in2[18]), .ZN(n17) );
  INVX0 U61 ( .INP(in2[19]), .ZN(n18) );
  INVX0 U62 ( .INP(in2[20]), .ZN(n19) );
  INVX0 U63 ( .INP(in2[21]), .ZN(n20) );
  INVX0 U64 ( .INP(in2[22]), .ZN(n21) );
  INVX0 U65 ( .INP(in1[1]), .ZN(n22) );
  INVX0 U66 ( .INP(in1[2]), .ZN(n111) );
  INVX0 U67 ( .INP(n138), .ZN(n140) );
  NOR2X0 U68 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n25) );
  AOI21X1 U69 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n25), .QN(n27) );
  NOR2X0 U70 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U71 ( .IN1(n24), .IN2(in2[0]), .IN3(n138), .IN4(n27), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U72 ( .INP(n133), .ZN(n67) );
  NOR2X0 U73 ( .IN1(n67), .IN2(n6), .QN(n28) );
  OA21X1 U74 ( .IN1(n25), .IN2(n6), .IN3(n30), .Q(n29) );
  AO22X1 U75 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n29), .Q(n26) );
  AOI22X1 U76 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n29), .QN(n32) );
  NOR2X0 U77 ( .IN1(in2[3]), .IN2(n30), .QN(n33) );
  AO21X1 U78 ( .IN1(in2[3]), .IN2(n30), .IN3(n33), .Q(n34) );
  OA22X1 U79 ( .IN1(n6), .IN2(n130), .IN3(n140), .IN4(n34), .Q(n31) );
  OA21X1 U80 ( .IN1(n33), .IN2(n7), .IN3(n37), .Q(n38) );
  AOI22X1 U81 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n38), .QN(n36) );
  OA22X1 U82 ( .IN1(n67), .IN2(n7), .IN3(n141), .IN4(n34), .Q(n35) );
  NOR2X0 U83 ( .IN1(in2[5]), .IN2(n37), .QN(n41) );
  AO21X1 U84 ( .IN1(in2[5]), .IN2(n37), .IN3(n41), .Q(n42) );
  OA22X1 U85 ( .IN1(n7), .IN2(n130), .IN3(n140), .IN4(n42), .Q(n40) );
  AOI22X1 U86 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n38), .QN(n39) );
  OA21X1 U87 ( .IN1(n41), .IN2(n8), .IN3(n45), .Q(n46) );
  AOI22X1 U88 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n46), .QN(n44) );
  OA22X1 U89 ( .IN1(n67), .IN2(n8), .IN3(n141), .IN4(n42), .Q(n43) );
  NOR2X0 U90 ( .IN1(in2[7]), .IN2(n45), .QN(n49) );
  AO21X1 U91 ( .IN1(in2[7]), .IN2(n45), .IN3(n49), .Q(n50) );
  OA22X1 U92 ( .IN1(n8), .IN2(n130), .IN3(n140), .IN4(n50), .Q(n48) );
  AOI22X1 U93 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n46), .QN(n47) );
  OA21X1 U94 ( .IN1(n49), .IN2(n9), .IN3(n53), .Q(n54) );
  AOI22X1 U95 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n54), .QN(n52) );
  OA22X1 U96 ( .IN1(n67), .IN2(n9), .IN3(n141), .IN4(n50), .Q(n51) );
  NOR2X0 U97 ( .IN1(in2[9]), .IN2(n53), .QN(n57) );
  AO21X1 U98 ( .IN1(in2[9]), .IN2(n53), .IN3(n57), .Q(n58) );
  OA22X1 U99 ( .IN1(n9), .IN2(n130), .IN3(n140), .IN4(n58), .Q(n56) );
  AOI22X1 U100 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n54), .QN(n55) );
  OA21X1 U101 ( .IN1(n57), .IN2(n10), .IN3(n61), .Q(n62) );
  AOI22X1 U102 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n62), .QN(n60) );
  OA22X1 U103 ( .IN1(n67), .IN2(n10), .IN3(n141), .IN4(n58), .Q(n59) );
  NOR2X0 U104 ( .IN1(in2[11]), .IN2(n61), .QN(n65) );
  AO21X1 U105 ( .IN1(in2[11]), .IN2(n61), .IN3(n65), .Q(n66) );
  OA22X1 U106 ( .IN1(n10), .IN2(n130), .IN3(n140), .IN4(n66), .Q(n64) );
  AOI22X1 U107 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n62), .QN(n63) );
  OA21X1 U108 ( .IN1(n65), .IN2(n11), .IN3(n77), .Q(n70) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n70), .QN(n69) );
  OA22X1 U110 ( .IN1(n67), .IN2(n11), .IN3(n141), .IN4(n66), .Q(n68) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n12), .S(n71), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n11), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n13), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n12), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n12), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n14), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n13), .IN4(n85), .IN5(n84), 
        .Q(out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n15), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n14), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n14), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n16), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n15), .IN4(n97), .IN5(n96), 
        .Q(out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n17), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n16), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n16), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n18), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n17), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n19), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n18), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n18), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n20), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n19), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n21), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n20), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n20), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n21), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_31 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n41), .IN2(n8), .QN(n45) );
  NAND2X0 U4 ( .IN1(n49), .IN2(n9), .QN(n53) );
  NAND2X0 U5 ( .IN1(n57), .IN2(n10), .QN(n61) );
  NAND2X0 U6 ( .IN1(n33), .IN2(n7), .QN(n37) );
  NAND2X0 U7 ( .IN1(n25), .IN2(n6), .QN(n30) );
  NAND2X0 U8 ( .IN1(n65), .IN2(n11), .QN(n77) );
  NAND2X0 U9 ( .IN1(n81), .IN2(n13), .QN(n89) );
  NAND2X0 U10 ( .IN1(n93), .IN2(n15), .QN(n101) );
  NAND2X0 U11 ( .IN1(in1[2]), .IN2(n77), .QN(n71) );
  NAND2X0 U12 ( .IN1(n70), .IN2(n132), .QN(n74) );
  NAND2X0 U13 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U14 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U15 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U16 ( .IN1(n118), .IN2(n19), .QN(n125) );
  NAND2X0 U17 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U18 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U19 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U20 ( .IN1(n27), .IN2(n132), .QN(n4) );
  NAND2X0 U21 ( .IN1(n141), .IN2(n130), .QN(n24) );
  NAND2X0 U22 ( .IN1(n40), .IN2(n39), .QN(out1[5]) );
  NAND2X0 U23 ( .IN1(n44), .IN2(n43), .QN(out1[6]) );
  NAND2X0 U24 ( .IN1(n48), .IN2(n47), .QN(out1[7]) );
  NAND2X0 U25 ( .IN1(n52), .IN2(n51), .QN(out1[8]) );
  NAND2X0 U26 ( .IN1(n56), .IN2(n55), .QN(out1[9]) );
  NAND2X0 U27 ( .IN1(n60), .IN2(n59), .QN(out1[10]) );
  NAND2X0 U28 ( .IN1(n64), .IN2(n63), .QN(out1[11]) );
  NAND2X0 U29 ( .IN1(n69), .IN2(n68), .QN(out1[12]) );
  NAND2X0 U30 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U31 ( .IN1(n105), .IN2(n17), .QN(n114) );
  NAND2X0 U32 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U33 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U34 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U35 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NAND2X0 U36 ( .IN1(n32), .IN2(n31), .QN(out1[3]) );
  NAND2X0 U37 ( .IN1(n36), .IN2(n35), .QN(out1[4]) );
  NAND2X0 U38 ( .IN1(n23), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U39 ( .IN1(in1[2]), .IN2(n22), .QN(n23) );
  INVX0 U40 ( .INP(in1[2]), .ZN(n111) );
  NOR2X0 U41 ( .IN1(n28), .IN2(n26), .QN(n3) );
  NOR2X0 U42 ( .IN1(n142), .IN2(n21), .QN(n1) );
  INVX0 U43 ( .INP(n132), .ZN(n141) );
  INVX0 U44 ( .INP(n130), .ZN(n137) );
  NOR2X0 U45 ( .IN1(n142), .IN2(n111), .QN(n138) );
  MUX21X1 U46 ( .IN1(n22), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  NAND3X0 U47 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  NOR3X0 U48 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  INVX0 U49 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U50 ( .INP(in2[2]), .ZN(n6) );
  INVX0 U51 ( .INP(in2[4]), .ZN(n7) );
  INVX0 U52 ( .INP(in2[6]), .ZN(n8) );
  INVX0 U53 ( .INP(in2[8]), .ZN(n9) );
  INVX0 U54 ( .INP(in2[10]), .ZN(n10) );
  INVX0 U55 ( .INP(in2[12]), .ZN(n11) );
  INVX0 U56 ( .INP(in2[13]), .ZN(n12) );
  INVX0 U57 ( .INP(in2[14]), .ZN(n13) );
  INVX0 U58 ( .INP(in2[15]), .ZN(n14) );
  INVX0 U59 ( .INP(in2[16]), .ZN(n15) );
  INVX0 U60 ( .INP(in2[17]), .ZN(n16) );
  INVX0 U61 ( .INP(in2[18]), .ZN(n17) );
  INVX0 U62 ( .INP(in2[19]), .ZN(n18) );
  INVX0 U63 ( .INP(in2[20]), .ZN(n19) );
  INVX0 U64 ( .INP(in2[21]), .ZN(n20) );
  INVX0 U65 ( .INP(in2[22]), .ZN(n21) );
  INVX0 U66 ( .INP(in1[1]), .ZN(n22) );
  INVX0 U67 ( .INP(n138), .ZN(n140) );
  NOR2X0 U68 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n25) );
  AOI21X1 U69 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n25), .QN(n27) );
  NOR2X0 U70 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U71 ( .IN1(n24), .IN2(in2[0]), .IN3(n138), .IN4(n27), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U72 ( .INP(n133), .ZN(n67) );
  NOR2X0 U73 ( .IN1(n67), .IN2(n6), .QN(n28) );
  OA21X1 U74 ( .IN1(n25), .IN2(n6), .IN3(n30), .Q(n29) );
  AO22X1 U75 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n29), .Q(n26) );
  AOI22X1 U76 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n29), .QN(n32) );
  NOR2X0 U77 ( .IN1(in2[3]), .IN2(n30), .QN(n33) );
  AO21X1 U78 ( .IN1(in2[3]), .IN2(n30), .IN3(n33), .Q(n34) );
  OA22X1 U79 ( .IN1(n6), .IN2(n130), .IN3(n140), .IN4(n34), .Q(n31) );
  OA21X1 U80 ( .IN1(n33), .IN2(n7), .IN3(n37), .Q(n38) );
  AOI22X1 U81 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n38), .QN(n36) );
  OA22X1 U82 ( .IN1(n67), .IN2(n7), .IN3(n141), .IN4(n34), .Q(n35) );
  NOR2X0 U83 ( .IN1(in2[5]), .IN2(n37), .QN(n41) );
  AO21X1 U84 ( .IN1(in2[5]), .IN2(n37), .IN3(n41), .Q(n42) );
  OA22X1 U85 ( .IN1(n7), .IN2(n130), .IN3(n140), .IN4(n42), .Q(n40) );
  AOI22X1 U86 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n38), .QN(n39) );
  OA21X1 U87 ( .IN1(n41), .IN2(n8), .IN3(n45), .Q(n46) );
  AOI22X1 U88 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n46), .QN(n44) );
  OA22X1 U89 ( .IN1(n67), .IN2(n8), .IN3(n141), .IN4(n42), .Q(n43) );
  NOR2X0 U90 ( .IN1(in2[7]), .IN2(n45), .QN(n49) );
  AO21X1 U91 ( .IN1(in2[7]), .IN2(n45), .IN3(n49), .Q(n50) );
  OA22X1 U92 ( .IN1(n8), .IN2(n130), .IN3(n140), .IN4(n50), .Q(n48) );
  AOI22X1 U93 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n46), .QN(n47) );
  OA21X1 U94 ( .IN1(n49), .IN2(n9), .IN3(n53), .Q(n54) );
  AOI22X1 U95 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n54), .QN(n52) );
  OA22X1 U96 ( .IN1(n67), .IN2(n9), .IN3(n141), .IN4(n50), .Q(n51) );
  NOR2X0 U97 ( .IN1(in2[9]), .IN2(n53), .QN(n57) );
  AO21X1 U98 ( .IN1(in2[9]), .IN2(n53), .IN3(n57), .Q(n58) );
  OA22X1 U99 ( .IN1(n9), .IN2(n130), .IN3(n140), .IN4(n58), .Q(n56) );
  AOI22X1 U100 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n54), .QN(n55) );
  OA21X1 U101 ( .IN1(n57), .IN2(n10), .IN3(n61), .Q(n62) );
  AOI22X1 U102 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n62), .QN(n60) );
  OA22X1 U103 ( .IN1(n67), .IN2(n10), .IN3(n141), .IN4(n58), .Q(n59) );
  NOR2X0 U104 ( .IN1(in2[11]), .IN2(n61), .QN(n65) );
  AO21X1 U105 ( .IN1(in2[11]), .IN2(n61), .IN3(n65), .Q(n66) );
  OA22X1 U106 ( .IN1(n10), .IN2(n130), .IN3(n140), .IN4(n66), .Q(n64) );
  AOI22X1 U107 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n62), .QN(n63) );
  OA21X1 U108 ( .IN1(n65), .IN2(n11), .IN3(n77), .Q(n70) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n70), .QN(n69) );
  OA22X1 U110 ( .IN1(n67), .IN2(n11), .IN3(n141), .IN4(n66), .Q(n68) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n12), .S(n71), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n11), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n13), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n12), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n12), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n14), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n13), .IN4(n85), .IN5(n84), 
        .Q(out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n15), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n14), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n14), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n16), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n15), .IN4(n97), .IN5(n96), 
        .Q(out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n17), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n16), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n16), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n18), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n17), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n19), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n18), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n18), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n20), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n19), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n21), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n20), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n20), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n21), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_32 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90;

  NAND2X0 U3 ( .IN1(n31), .IN2(n6), .QN(n33) );
  NAND2X0 U4 ( .IN1(n35), .IN2(n7), .QN(n37) );
  NAND2X0 U5 ( .IN1(n39), .IN2(n8), .QN(n44) );
  NAND2X0 U6 ( .IN1(n23), .IN2(n4), .QN(n25) );
  NAND2X0 U7 ( .IN1(n27), .IN2(n5), .QN(n29) );
  NAND2X0 U8 ( .IN1(in1[2]), .IN2(n44), .QN(n41) );
  NAND2X0 U9 ( .IN1(n49), .IN2(n10), .QN(n52) );
  NAND2X0 U10 ( .IN1(in1[2]), .IN2(n52), .QN(n48) );
  NAND2X0 U11 ( .IN1(n57), .IN2(n12), .QN(n60) );
  NAND2X0 U12 ( .IN1(in1[2]), .IN2(n60), .QN(n56) );
  NAND2X0 U13 ( .IN1(n65), .IN2(n14), .QN(n68) );
  NAND2X0 U14 ( .IN1(in1[2]), .IN2(n68), .QN(n64) );
  NAND2X0 U15 ( .IN1(n75), .IN2(n16), .QN(n79) );
  NAND2X0 U16 ( .IN1(n72), .IN2(in1[2]), .QN(n83) );
  NAND2X0 U17 ( .IN1(in1[2]), .IN2(n79), .QN(n74) );
  INVX0 U18 ( .INP(n83), .ZN(n86) );
  NOR2X0 U19 ( .IN1(n72), .IN2(n69), .QN(n89) );
  NOR2X0 U20 ( .IN1(in1[2]), .IN2(n72), .QN(n87) );
  NBUFFX2 U21 ( .INP(in1[2]), .Z(out1[26]) );
  NBUFFX2 U22 ( .INP(in1[2]), .Z(out1[25]) );
  INVX0 U23 ( .INP(in2[2]), .ZN(n3) );
  INVX0 U24 ( .INP(in2[4]), .ZN(n4) );
  INVX0 U25 ( .INP(in2[6]), .ZN(n5) );
  INVX0 U26 ( .INP(in2[8]), .ZN(n6) );
  INVX0 U27 ( .INP(in2[10]), .ZN(n7) );
  INVX0 U28 ( .INP(in2[12]), .ZN(n8) );
  INVX0 U29 ( .INP(in2[13]), .ZN(n9) );
  INVX0 U30 ( .INP(in2[14]), .ZN(n10) );
  INVX0 U31 ( .INP(in2[15]), .ZN(n11) );
  INVX0 U32 ( .INP(in2[16]), .ZN(n12) );
  INVX0 U33 ( .INP(in2[17]), .ZN(n13) );
  INVX0 U34 ( .INP(in2[18]), .ZN(n14) );
  INVX0 U35 ( .INP(in2[19]), .ZN(n15) );
  INVX0 U36 ( .INP(in2[20]), .ZN(n16) );
  INVX0 U37 ( .INP(in2[21]), .ZN(n17) );
  INVX0 U38 ( .INP(in2[22]), .ZN(n18) );
  INVX0 U39 ( .INP(in1[1]), .ZN(n72) );
  INVX0 U40 ( .INP(in1[2]), .ZN(n69) );
  NOR2X0 U41 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n19) );
  AOI21X1 U42 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n19), .QN(n20) );
  AO222X1 U43 ( .IN1(in2[0]), .IN2(n86), .IN3(in2[1]), .IN4(n87), .IN5(n89), 
        .IN6(n20), .Q(out1[1]) );
  OR3X1 U44 ( .IN1(in2[2]), .IN2(in2[0]), .IN3(in2[1]), .Q(n21) );
  OA21X1 U45 ( .IN1(n19), .IN2(n3), .IN3(n21), .Q(n22) );
  AO222X1 U46 ( .IN1(in2[2]), .IN2(n87), .IN3(n86), .IN4(n20), .IN5(n22), 
        .IN6(n89), .Q(out1[2]) );
  NOR2X0 U47 ( .IN1(in2[3]), .IN2(n21), .QN(n23) );
  AOI21X1 U48 ( .IN1(in2[3]), .IN2(n21), .IN3(n23), .QN(n24) );
  AO222X1 U49 ( .IN1(in2[3]), .IN2(n87), .IN3(n86), .IN4(n22), .IN5(n24), 
        .IN6(n89), .Q(out1[3]) );
  OA21X1 U50 ( .IN1(n23), .IN2(n4), .IN3(n25), .Q(n26) );
  AO222X1 U51 ( .IN1(in2[4]), .IN2(n87), .IN3(n86), .IN4(n24), .IN5(n26), 
        .IN6(n89), .Q(out1[4]) );
  NOR2X0 U52 ( .IN1(in2[5]), .IN2(n25), .QN(n27) );
  AOI21X1 U53 ( .IN1(in2[5]), .IN2(n25), .IN3(n27), .QN(n28) );
  AO222X1 U54 ( .IN1(in2[5]), .IN2(n87), .IN3(n86), .IN4(n26), .IN5(n28), 
        .IN6(n89), .Q(out1[5]) );
  OA21X1 U55 ( .IN1(n27), .IN2(n5), .IN3(n29), .Q(n30) );
  AO222X1 U56 ( .IN1(in2[6]), .IN2(n87), .IN3(n86), .IN4(n28), .IN5(n30), 
        .IN6(n89), .Q(out1[6]) );
  NOR2X0 U57 ( .IN1(in2[7]), .IN2(n29), .QN(n31) );
  AOI21X1 U58 ( .IN1(in2[7]), .IN2(n29), .IN3(n31), .QN(n32) );
  AO222X1 U59 ( .IN1(in2[7]), .IN2(n87), .IN3(n86), .IN4(n30), .IN5(n32), 
        .IN6(n89), .Q(out1[7]) );
  OA21X1 U60 ( .IN1(n31), .IN2(n6), .IN3(n33), .Q(n34) );
  AO222X1 U61 ( .IN1(in2[8]), .IN2(n87), .IN3(n86), .IN4(n32), .IN5(n34), 
        .IN6(n89), .Q(out1[8]) );
  NOR2X0 U62 ( .IN1(in2[9]), .IN2(n33), .QN(n35) );
  AOI21X1 U63 ( .IN1(in2[9]), .IN2(n33), .IN3(n35), .QN(n36) );
  AO222X1 U64 ( .IN1(in2[9]), .IN2(n87), .IN3(n86), .IN4(n34), .IN5(n36), 
        .IN6(n89), .Q(out1[9]) );
  OA21X1 U65 ( .IN1(n35), .IN2(n7), .IN3(n37), .Q(n38) );
  AO222X1 U66 ( .IN1(in2[10]), .IN2(n87), .IN3(n86), .IN4(n36), .IN5(n38), 
        .IN6(n89), .Q(out1[10]) );
  NOR2X0 U67 ( .IN1(in2[11]), .IN2(n37), .QN(n39) );
  AOI21X1 U68 ( .IN1(in2[11]), .IN2(n37), .IN3(n39), .QN(n40) );
  AO222X1 U69 ( .IN1(in2[11]), .IN2(n87), .IN3(n86), .IN4(n38), .IN5(n40), 
        .IN6(n89), .Q(out1[11]) );
  OA21X1 U70 ( .IN1(n39), .IN2(n8), .IN3(n44), .Q(n42) );
  AO222X1 U71 ( .IN1(in2[12]), .IN2(n87), .IN3(n86), .IN4(n40), .IN5(n42), 
        .IN6(n89), .Q(out1[12]) );
  MUX21X1 U72 ( .IN1(n9), .IN2(in2[13]), .S(n41), .Q(n43) );
  AO22X1 U73 ( .IN1(in1[1]), .IN2(n43), .IN3(n86), .IN4(n42), .Q(out1[13]) );
  NOR2X0 U74 ( .IN1(in2[13]), .IN2(n44), .QN(n49) );
  AO21X1 U75 ( .IN1(in2[13]), .IN2(n44), .IN3(n83), .Q(n47) );
  NOR2X0 U76 ( .IN1(n49), .IN2(n69), .QN(n45) );
  MUX21X1 U77 ( .IN1(n10), .IN2(in2[14]), .S(n45), .Q(n46) );
  OAI22X1 U78 ( .IN1(n49), .IN2(n47), .IN3(n72), .IN4(n46), .QN(out1[14]) );
  MUX21X1 U79 ( .IN1(n11), .IN2(in2[15]), .S(n48), .Q(n51) );
  OA21X1 U80 ( .IN1(n49), .IN2(n10), .IN3(n86), .Q(n50) );
  AO22X1 U81 ( .IN1(in1[1]), .IN2(n51), .IN3(n50), .IN4(n52), .Q(out1[15]) );
  NOR2X0 U82 ( .IN1(in2[15]), .IN2(n52), .QN(n57) );
  AO21X1 U83 ( .IN1(in2[15]), .IN2(n52), .IN3(n83), .Q(n55) );
  NOR2X0 U84 ( .IN1(n57), .IN2(n69), .QN(n53) );
  MUX21X1 U85 ( .IN1(n12), .IN2(in2[16]), .S(n53), .Q(n54) );
  OAI22X1 U86 ( .IN1(n57), .IN2(n55), .IN3(n72), .IN4(n54), .QN(out1[16]) );
  MUX21X1 U87 ( .IN1(n13), .IN2(in2[17]), .S(n56), .Q(n59) );
  OA21X1 U88 ( .IN1(n57), .IN2(n12), .IN3(n86), .Q(n58) );
  AO22X1 U89 ( .IN1(in1[1]), .IN2(n59), .IN3(n58), .IN4(n60), .Q(out1[17]) );
  NOR2X0 U90 ( .IN1(in2[17]), .IN2(n60), .QN(n65) );
  AO21X1 U91 ( .IN1(in2[17]), .IN2(n60), .IN3(n83), .Q(n63) );
  NOR2X0 U92 ( .IN1(n65), .IN2(n69), .QN(n61) );
  MUX21X1 U93 ( .IN1(n14), .IN2(in2[18]), .S(n61), .Q(n62) );
  OAI22X1 U94 ( .IN1(n65), .IN2(n63), .IN3(n72), .IN4(n62), .QN(out1[18]) );
  MUX21X1 U95 ( .IN1(n15), .IN2(in2[19]), .S(n64), .Q(n67) );
  OA21X1 U96 ( .IN1(n65), .IN2(n14), .IN3(n86), .Q(n66) );
  AO22X1 U97 ( .IN1(in1[1]), .IN2(n67), .IN3(n66), .IN4(n68), .Q(out1[19]) );
  NOR2X0 U98 ( .IN1(in2[19]), .IN2(n68), .QN(n75) );
  AO21X1 U99 ( .IN1(in2[19]), .IN2(n68), .IN3(n83), .Q(n73) );
  NOR2X0 U100 ( .IN1(n75), .IN2(n69), .QN(n70) );
  MUX21X1 U101 ( .IN1(n16), .IN2(in2[20]), .S(n70), .Q(n71) );
  OAI22X1 U102 ( .IN1(n75), .IN2(n73), .IN3(n72), .IN4(n71), .QN(out1[20]) );
  MUX21X1 U103 ( .IN1(n17), .IN2(in2[21]), .S(n74), .Q(n77) );
  MUX21X1 U104 ( .IN1(n16), .IN2(in2[20]), .S(n75), .Q(n76) );
  AO22X1 U105 ( .IN1(in1[1]), .IN2(n77), .IN3(n86), .IN4(n76), .Q(out1[21]) );
  INVX0 U106 ( .INP(n89), .ZN(n78) );
  OR2X1 U107 ( .IN1(n79), .IN2(in2[21]), .Q(n85) );
  NOR2X0 U108 ( .IN1(n78), .IN2(n85), .QN(n84) );
  NOR2X0 U109 ( .IN1(in2[22]), .IN2(n78), .QN(n81) );
  NAND2X0 U110 ( .IN1(in2[21]), .IN2(n79), .QN(n80) );
  OA221X1 U111 ( .IN1(n81), .IN2(n86), .IN3(n81), .IN4(n80), .IN5(n85), .Q(n82) );
  AO221X1 U112 ( .IN1(in2[22]), .IN2(n87), .IN3(in2[22]), .IN4(n84), .IN5(n82), 
        .Q(out1[22]) );
  NOR2X0 U113 ( .IN1(n83), .IN2(n85), .QN(n90) );
  AO21X1 U114 ( .IN1(n86), .IN2(n85), .IN3(n84), .Q(n88) );
  AO221X1 U115 ( .IN1(in2[22]), .IN2(n90), .IN3(n18), .IN4(n88), .IN5(n87), 
        .Q(out1[23]) );
  AO21X1 U116 ( .IN1(n90), .IN2(n18), .IN3(n89), .Q(out1[24]) );
  AND2X1 U117 ( .IN1(in1[1]), .IN2(in2[0]), .Q(out1[0]) );
endmodule


module booth27_33 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2;

  AND2X1 U3 ( .IN1(in1[1]), .IN2(in1[0]), .Q(out1[24]) );
  INVX0 U4 ( .INP(in1[1]), .ZN(n1) );
  MUX21X1 U5 ( .IN1(in1[1]), .IN2(n1), .S(in1[0]), .Q(n2) );
  AO22X1 U6 ( .IN1(in2[0]), .IN2(out1[24]), .IN3(in2[1]), .IN4(n2), .Q(out1[1]) );
  AO22X1 U7 ( .IN1(out1[24]), .IN2(in2[1]), .IN3(in2[2]), .IN4(n2), .Q(out1[2]) );
  AO22X1 U8 ( .IN1(out1[24]), .IN2(in2[2]), .IN3(in2[3]), .IN4(n2), .Q(out1[3]) );
  AO22X1 U9 ( .IN1(out1[24]), .IN2(in2[3]), .IN3(in2[4]), .IN4(n2), .Q(out1[4]) );
  AO22X1 U10 ( .IN1(out1[24]), .IN2(in2[4]), .IN3(in2[5]), .IN4(n2), .Q(
        out1[5]) );
  AO22X1 U11 ( .IN1(out1[24]), .IN2(in2[5]), .IN3(in2[6]), .IN4(n2), .Q(
        out1[6]) );
  AO22X1 U12 ( .IN1(out1[24]), .IN2(in2[6]), .IN3(in2[7]), .IN4(n2), .Q(
        out1[7]) );
  AO22X1 U13 ( .IN1(out1[24]), .IN2(in2[7]), .IN3(in2[8]), .IN4(n2), .Q(
        out1[8]) );
  AO22X1 U14 ( .IN1(out1[24]), .IN2(in2[8]), .IN3(in2[9]), .IN4(n2), .Q(
        out1[9]) );
  AO22X1 U15 ( .IN1(out1[24]), .IN2(in2[9]), .IN3(in2[10]), .IN4(n2), .Q(
        out1[10]) );
  AO22X1 U16 ( .IN1(out1[24]), .IN2(in2[10]), .IN3(in2[11]), .IN4(n2), .Q(
        out1[11]) );
  AO22X1 U17 ( .IN1(out1[24]), .IN2(in2[11]), .IN3(in2[12]), .IN4(n2), .Q(
        out1[12]) );
  AO22X1 U18 ( .IN1(out1[24]), .IN2(in2[12]), .IN3(in2[13]), .IN4(n2), .Q(
        out1[13]) );
  AO22X1 U19 ( .IN1(out1[24]), .IN2(in2[13]), .IN3(in2[14]), .IN4(n2), .Q(
        out1[14]) );
  AO22X1 U20 ( .IN1(out1[24]), .IN2(in2[14]), .IN3(in2[15]), .IN4(n2), .Q(
        out1[15]) );
  AO22X1 U21 ( .IN1(out1[24]), .IN2(in2[15]), .IN3(in2[16]), .IN4(n2), .Q(
        out1[16]) );
  AO22X1 U22 ( .IN1(out1[24]), .IN2(in2[16]), .IN3(in2[17]), .IN4(n2), .Q(
        out1[17]) );
  AO22X1 U23 ( .IN1(out1[24]), .IN2(in2[17]), .IN3(in2[18]), .IN4(n2), .Q(
        out1[18]) );
  AO22X1 U24 ( .IN1(out1[24]), .IN2(in2[18]), .IN3(in2[19]), .IN4(n2), .Q(
        out1[19]) );
  AO22X1 U25 ( .IN1(out1[24]), .IN2(in2[19]), .IN3(in2[20]), .IN4(n2), .Q(
        out1[20]) );
  AO22X1 U26 ( .IN1(out1[24]), .IN2(in2[20]), .IN3(in2[21]), .IN4(n2), .Q(
        out1[21]) );
  AO22X1 U27 ( .IN1(out1[24]), .IN2(in2[21]), .IN3(in2[22]), .IN4(n2), .Q(
        out1[22]) );
  AO21X1 U28 ( .IN1(out1[24]), .IN2(in2[22]), .IN3(n2), .Q(out1[23]) );
  AND2X1 U29 ( .IN1(in2[0]), .IN2(n2), .Q(out1[0]) );
endmodule


module booth27_34 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n57), .IN2(n10), .QN(n61) );
  NAND2X0 U4 ( .IN1(n25), .IN2(n6), .QN(n30) );
  NAND2X0 U5 ( .IN1(n33), .IN2(n7), .QN(n37) );
  NAND2X0 U6 ( .IN1(n49), .IN2(n9), .QN(n53) );
  NAND2X0 U7 ( .IN1(n41), .IN2(n8), .QN(n45) );
  NAND2X0 U8 ( .IN1(n65), .IN2(n11), .QN(n77) );
  NAND2X0 U9 ( .IN1(n81), .IN2(n13), .QN(n89) );
  NAND2X0 U10 ( .IN1(n93), .IN2(n15), .QN(n101) );
  NAND2X0 U11 ( .IN1(n105), .IN2(n17), .QN(n114) );
  NAND2X0 U12 ( .IN1(n118), .IN2(n19), .QN(n125) );
  NAND2X0 U13 ( .IN1(in1[2]), .IN2(n77), .QN(n71) );
  NAND2X0 U14 ( .IN1(n70), .IN2(n132), .QN(n74) );
  NAND2X0 U15 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U16 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U17 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U18 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U19 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U20 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U21 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U22 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U23 ( .IN1(n141), .IN2(n130), .QN(n24) );
  NAND2X0 U24 ( .IN1(n27), .IN2(n132), .QN(n4) );
  NAND2X0 U25 ( .IN1(n56), .IN2(n55), .QN(out1[9]) );
  NAND2X0 U26 ( .IN1(n60), .IN2(n59), .QN(out1[10]) );
  NAND2X0 U27 ( .IN1(n64), .IN2(n63), .QN(out1[11]) );
  NAND2X0 U28 ( .IN1(n69), .IN2(n68), .QN(out1[12]) );
  NAND2X0 U29 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U30 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U31 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NAND2X0 U32 ( .IN1(n32), .IN2(n31), .QN(out1[3]) );
  NAND2X0 U33 ( .IN1(n36), .IN2(n35), .QN(out1[4]) );
  NAND2X0 U34 ( .IN1(n40), .IN2(n39), .QN(out1[5]) );
  NAND2X0 U35 ( .IN1(n44), .IN2(n43), .QN(out1[6]) );
  NAND2X0 U36 ( .IN1(n48), .IN2(n47), .QN(out1[7]) );
  NAND2X0 U37 ( .IN1(n52), .IN2(n51), .QN(out1[8]) );
  NAND2X0 U38 ( .IN1(n23), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U39 ( .IN1(in1[2]), .IN2(n22), .QN(n23) );
  NOR2X0 U40 ( .IN1(n28), .IN2(n26), .QN(n3) );
  INVX0 U41 ( .INP(n130), .ZN(n137) );
  NAND3X0 U42 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  NOR2X0 U43 ( .IN1(n142), .IN2(n21), .QN(n1) );
  INVX0 U44 ( .INP(n132), .ZN(n141) );
  NOR3X0 U45 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  NOR2X0 U46 ( .IN1(n142), .IN2(n111), .QN(n138) );
  MUX21X1 U47 ( .IN1(n22), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  INVX0 U48 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U49 ( .INP(in2[2]), .ZN(n6) );
  INVX0 U50 ( .INP(in2[4]), .ZN(n7) );
  INVX0 U51 ( .INP(in2[6]), .ZN(n8) );
  INVX0 U52 ( .INP(in2[8]), .ZN(n9) );
  INVX0 U53 ( .INP(in2[10]), .ZN(n10) );
  INVX0 U54 ( .INP(in2[12]), .ZN(n11) );
  INVX0 U55 ( .INP(in2[13]), .ZN(n12) );
  INVX0 U56 ( .INP(in2[14]), .ZN(n13) );
  INVX0 U57 ( .INP(in2[15]), .ZN(n14) );
  INVX0 U58 ( .INP(in2[16]), .ZN(n15) );
  INVX0 U59 ( .INP(in2[17]), .ZN(n16) );
  INVX0 U60 ( .INP(in2[18]), .ZN(n17) );
  INVX0 U61 ( .INP(in2[19]), .ZN(n18) );
  INVX0 U62 ( .INP(in2[20]), .ZN(n19) );
  INVX0 U63 ( .INP(in2[21]), .ZN(n20) );
  INVX0 U64 ( .INP(in2[22]), .ZN(n21) );
  INVX0 U65 ( .INP(in1[1]), .ZN(n22) );
  INVX0 U66 ( .INP(in1[2]), .ZN(n111) );
  INVX0 U67 ( .INP(n138), .ZN(n140) );
  NOR2X0 U68 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n25) );
  AOI21X1 U69 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n25), .QN(n27) );
  NOR2X0 U70 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U71 ( .IN1(n24), .IN2(in2[0]), .IN3(n138), .IN4(n27), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U72 ( .INP(n133), .ZN(n67) );
  NOR2X0 U73 ( .IN1(n67), .IN2(n6), .QN(n28) );
  OA21X1 U74 ( .IN1(n25), .IN2(n6), .IN3(n30), .Q(n29) );
  AO22X1 U75 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n29), .Q(n26) );
  AOI22X1 U76 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n29), .QN(n32) );
  NOR2X0 U77 ( .IN1(in2[3]), .IN2(n30), .QN(n33) );
  AO21X1 U78 ( .IN1(in2[3]), .IN2(n30), .IN3(n33), .Q(n34) );
  OA22X1 U79 ( .IN1(n6), .IN2(n130), .IN3(n140), .IN4(n34), .Q(n31) );
  OA21X1 U80 ( .IN1(n33), .IN2(n7), .IN3(n37), .Q(n38) );
  AOI22X1 U81 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n38), .QN(n36) );
  OA22X1 U82 ( .IN1(n67), .IN2(n7), .IN3(n141), .IN4(n34), .Q(n35) );
  NOR2X0 U83 ( .IN1(in2[5]), .IN2(n37), .QN(n41) );
  AO21X1 U84 ( .IN1(in2[5]), .IN2(n37), .IN3(n41), .Q(n42) );
  OA22X1 U85 ( .IN1(n7), .IN2(n130), .IN3(n140), .IN4(n42), .Q(n40) );
  AOI22X1 U86 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n38), .QN(n39) );
  OA21X1 U87 ( .IN1(n41), .IN2(n8), .IN3(n45), .Q(n46) );
  AOI22X1 U88 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n46), .QN(n44) );
  OA22X1 U89 ( .IN1(n67), .IN2(n8), .IN3(n141), .IN4(n42), .Q(n43) );
  NOR2X0 U90 ( .IN1(in2[7]), .IN2(n45), .QN(n49) );
  AO21X1 U91 ( .IN1(in2[7]), .IN2(n45), .IN3(n49), .Q(n50) );
  OA22X1 U92 ( .IN1(n8), .IN2(n130), .IN3(n140), .IN4(n50), .Q(n48) );
  AOI22X1 U93 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n46), .QN(n47) );
  OA21X1 U94 ( .IN1(n49), .IN2(n9), .IN3(n53), .Q(n54) );
  AOI22X1 U95 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n54), .QN(n52) );
  OA22X1 U96 ( .IN1(n67), .IN2(n9), .IN3(n141), .IN4(n50), .Q(n51) );
  NOR2X0 U97 ( .IN1(in2[9]), .IN2(n53), .QN(n57) );
  AO21X1 U98 ( .IN1(in2[9]), .IN2(n53), .IN3(n57), .Q(n58) );
  OA22X1 U99 ( .IN1(n9), .IN2(n130), .IN3(n140), .IN4(n58), .Q(n56) );
  AOI22X1 U100 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n54), .QN(n55) );
  OA21X1 U101 ( .IN1(n57), .IN2(n10), .IN3(n61), .Q(n62) );
  AOI22X1 U102 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n62), .QN(n60) );
  OA22X1 U103 ( .IN1(n67), .IN2(n10), .IN3(n141), .IN4(n58), .Q(n59) );
  NOR2X0 U104 ( .IN1(in2[11]), .IN2(n61), .QN(n65) );
  AO21X1 U105 ( .IN1(in2[11]), .IN2(n61), .IN3(n65), .Q(n66) );
  OA22X1 U106 ( .IN1(n10), .IN2(n130), .IN3(n140), .IN4(n66), .Q(n64) );
  AOI22X1 U107 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n62), .QN(n63) );
  OA21X1 U108 ( .IN1(n65), .IN2(n11), .IN3(n77), .Q(n70) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n70), .QN(n69) );
  OA22X1 U110 ( .IN1(n67), .IN2(n11), .IN3(n141), .IN4(n66), .Q(n68) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n12), .S(n71), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n11), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n13), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n12), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n12), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n14), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n13), .IN4(n85), .IN5(n84), 
        .Q(out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n15), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n14), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n14), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n16), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n15), .IN4(n97), .IN5(n96), 
        .Q(out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n17), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n16), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n16), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n18), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n17), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n19), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n18), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n18), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n20), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n19), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n21), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n20), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n20), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n21), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_35 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n25), .IN2(n6), .QN(n30) );
  NAND2X0 U4 ( .IN1(n33), .IN2(n7), .QN(n37) );
  NAND2X0 U5 ( .IN1(n41), .IN2(n8), .QN(n45) );
  NAND2X0 U6 ( .IN1(n57), .IN2(n10), .QN(n61) );
  NAND2X0 U7 ( .IN1(n49), .IN2(n9), .QN(n53) );
  NAND2X0 U8 ( .IN1(n65), .IN2(n11), .QN(n77) );
  NAND2X0 U9 ( .IN1(n81), .IN2(n13), .QN(n89) );
  NAND2X0 U10 ( .IN1(n93), .IN2(n15), .QN(n101) );
  NAND2X0 U11 ( .IN1(n105), .IN2(n17), .QN(n114) );
  NAND2X0 U12 ( .IN1(n118), .IN2(n19), .QN(n125) );
  NAND2X0 U13 ( .IN1(in1[2]), .IN2(n77), .QN(n71) );
  NAND2X0 U14 ( .IN1(n70), .IN2(n132), .QN(n74) );
  NAND2X0 U15 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U16 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U17 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U18 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U19 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U20 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U21 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U22 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U23 ( .IN1(n141), .IN2(n130), .QN(n24) );
  NAND2X0 U24 ( .IN1(n27), .IN2(n132), .QN(n4) );
  NAND2X0 U25 ( .IN1(n64), .IN2(n63), .QN(out1[11]) );
  NAND2X0 U26 ( .IN1(n69), .IN2(n68), .QN(out1[12]) );
  NAND2X0 U27 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U28 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U29 ( .IN1(n23), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U30 ( .IN1(in1[2]), .IN2(n22), .QN(n23) );
  NAND2X0 U31 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NAND2X0 U32 ( .IN1(n32), .IN2(n31), .QN(out1[3]) );
  NAND2X0 U33 ( .IN1(n36), .IN2(n35), .QN(out1[4]) );
  NAND2X0 U34 ( .IN1(n40), .IN2(n39), .QN(out1[5]) );
  NAND2X0 U35 ( .IN1(n44), .IN2(n43), .QN(out1[6]) );
  NAND2X0 U36 ( .IN1(n48), .IN2(n47), .QN(out1[7]) );
  NAND2X0 U37 ( .IN1(n52), .IN2(n51), .QN(out1[8]) );
  NAND2X0 U38 ( .IN1(n56), .IN2(n55), .QN(out1[9]) );
  NAND2X0 U39 ( .IN1(n60), .IN2(n59), .QN(out1[10]) );
  NOR2X0 U40 ( .IN1(n28), .IN2(n26), .QN(n3) );
  NOR2X0 U41 ( .IN1(n142), .IN2(n21), .QN(n1) );
  INVX0 U42 ( .INP(n132), .ZN(n141) );
  INVX0 U43 ( .INP(n130), .ZN(n137) );
  NAND3X0 U44 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  NOR3X0 U45 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  NOR2X0 U46 ( .IN1(n142), .IN2(n111), .QN(n138) );
  MUX21X1 U47 ( .IN1(n22), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  INVX0 U48 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U49 ( .INP(in2[2]), .ZN(n6) );
  INVX0 U50 ( .INP(in2[4]), .ZN(n7) );
  INVX0 U51 ( .INP(in2[6]), .ZN(n8) );
  INVX0 U52 ( .INP(in2[8]), .ZN(n9) );
  INVX0 U53 ( .INP(in2[10]), .ZN(n10) );
  INVX0 U54 ( .INP(in2[12]), .ZN(n11) );
  INVX0 U55 ( .INP(in2[13]), .ZN(n12) );
  INVX0 U56 ( .INP(in2[14]), .ZN(n13) );
  INVX0 U57 ( .INP(in2[15]), .ZN(n14) );
  INVX0 U58 ( .INP(in2[16]), .ZN(n15) );
  INVX0 U59 ( .INP(in2[17]), .ZN(n16) );
  INVX0 U60 ( .INP(in2[18]), .ZN(n17) );
  INVX0 U61 ( .INP(in2[19]), .ZN(n18) );
  INVX0 U62 ( .INP(in2[20]), .ZN(n19) );
  INVX0 U63 ( .INP(in2[21]), .ZN(n20) );
  INVX0 U64 ( .INP(in2[22]), .ZN(n21) );
  INVX0 U65 ( .INP(in1[1]), .ZN(n22) );
  INVX0 U66 ( .INP(in1[2]), .ZN(n111) );
  INVX0 U67 ( .INP(n138), .ZN(n140) );
  NOR2X0 U68 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n25) );
  AOI21X1 U69 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n25), .QN(n27) );
  NOR2X0 U70 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U71 ( .IN1(n24), .IN2(in2[0]), .IN3(n138), .IN4(n27), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U72 ( .INP(n133), .ZN(n67) );
  NOR2X0 U73 ( .IN1(n67), .IN2(n6), .QN(n28) );
  OA21X1 U74 ( .IN1(n25), .IN2(n6), .IN3(n30), .Q(n29) );
  AO22X1 U75 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n29), .Q(n26) );
  AOI22X1 U76 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n29), .QN(n32) );
  NOR2X0 U77 ( .IN1(in2[3]), .IN2(n30), .QN(n33) );
  AO21X1 U78 ( .IN1(in2[3]), .IN2(n30), .IN3(n33), .Q(n34) );
  OA22X1 U79 ( .IN1(n6), .IN2(n130), .IN3(n140), .IN4(n34), .Q(n31) );
  OA21X1 U80 ( .IN1(n33), .IN2(n7), .IN3(n37), .Q(n38) );
  AOI22X1 U81 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n38), .QN(n36) );
  OA22X1 U82 ( .IN1(n67), .IN2(n7), .IN3(n141), .IN4(n34), .Q(n35) );
  NOR2X0 U83 ( .IN1(in2[5]), .IN2(n37), .QN(n41) );
  AO21X1 U84 ( .IN1(in2[5]), .IN2(n37), .IN3(n41), .Q(n42) );
  OA22X1 U85 ( .IN1(n7), .IN2(n130), .IN3(n140), .IN4(n42), .Q(n40) );
  AOI22X1 U86 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n38), .QN(n39) );
  OA21X1 U87 ( .IN1(n41), .IN2(n8), .IN3(n45), .Q(n46) );
  AOI22X1 U88 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n46), .QN(n44) );
  OA22X1 U89 ( .IN1(n67), .IN2(n8), .IN3(n141), .IN4(n42), .Q(n43) );
  NOR2X0 U90 ( .IN1(in2[7]), .IN2(n45), .QN(n49) );
  AO21X1 U91 ( .IN1(in2[7]), .IN2(n45), .IN3(n49), .Q(n50) );
  OA22X1 U92 ( .IN1(n8), .IN2(n130), .IN3(n140), .IN4(n50), .Q(n48) );
  AOI22X1 U93 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n46), .QN(n47) );
  OA21X1 U94 ( .IN1(n49), .IN2(n9), .IN3(n53), .Q(n54) );
  AOI22X1 U95 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n54), .QN(n52) );
  OA22X1 U96 ( .IN1(n67), .IN2(n9), .IN3(n141), .IN4(n50), .Q(n51) );
  NOR2X0 U97 ( .IN1(in2[9]), .IN2(n53), .QN(n57) );
  AO21X1 U98 ( .IN1(in2[9]), .IN2(n53), .IN3(n57), .Q(n58) );
  OA22X1 U99 ( .IN1(n9), .IN2(n130), .IN3(n140), .IN4(n58), .Q(n56) );
  AOI22X1 U100 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n54), .QN(n55) );
  OA21X1 U101 ( .IN1(n57), .IN2(n10), .IN3(n61), .Q(n62) );
  AOI22X1 U102 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n62), .QN(n60) );
  OA22X1 U103 ( .IN1(n67), .IN2(n10), .IN3(n141), .IN4(n58), .Q(n59) );
  NOR2X0 U104 ( .IN1(in2[11]), .IN2(n61), .QN(n65) );
  AO21X1 U105 ( .IN1(in2[11]), .IN2(n61), .IN3(n65), .Q(n66) );
  OA22X1 U106 ( .IN1(n10), .IN2(n130), .IN3(n140), .IN4(n66), .Q(n64) );
  AOI22X1 U107 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n62), .QN(n63) );
  OA21X1 U108 ( .IN1(n65), .IN2(n11), .IN3(n77), .Q(n70) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n70), .QN(n69) );
  OA22X1 U110 ( .IN1(n67), .IN2(n11), .IN3(n141), .IN4(n66), .Q(n68) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n12), .S(n71), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n11), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n13), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n12), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n12), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n14), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n13), .IN4(n85), .IN5(n84), 
        .Q(out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n15), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n14), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n14), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n16), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n15), .IN4(n97), .IN5(n96), 
        .Q(out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n17), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n16), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n16), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n18), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n17), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n19), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n18), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n18), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n20), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n19), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n21), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n20), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n20), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n21), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_36 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90;

  NAND2X0 U3 ( .IN1(n75), .IN2(n16), .QN(n79) );
  NAND2X0 U4 ( .IN1(n23), .IN2(n4), .QN(n25) );
  NAND2X0 U5 ( .IN1(n27), .IN2(n5), .QN(n29) );
  NAND2X0 U6 ( .IN1(n31), .IN2(n6), .QN(n33) );
  NAND2X0 U7 ( .IN1(n35), .IN2(n7), .QN(n37) );
  NAND2X0 U8 ( .IN1(n39), .IN2(n8), .QN(n44) );
  NAND2X0 U9 ( .IN1(in1[2]), .IN2(n44), .QN(n41) );
  NAND2X0 U10 ( .IN1(n49), .IN2(n10), .QN(n52) );
  NAND2X0 U11 ( .IN1(in1[2]), .IN2(n52), .QN(n48) );
  NAND2X0 U12 ( .IN1(n57), .IN2(n12), .QN(n60) );
  NAND2X0 U13 ( .IN1(in1[2]), .IN2(n60), .QN(n56) );
  NAND2X0 U14 ( .IN1(n65), .IN2(n14), .QN(n68) );
  NAND2X0 U15 ( .IN1(in1[2]), .IN2(n68), .QN(n64) );
  NAND2X0 U16 ( .IN1(in1[2]), .IN2(n79), .QN(n74) );
  NAND2X0 U17 ( .IN1(n72), .IN2(in1[2]), .QN(n83) );
  INVX0 U18 ( .INP(n83), .ZN(n86) );
  INVX0 U19 ( .INP(in1[0]), .ZN(n72) );
  NOR2X0 U20 ( .IN1(in1[2]), .IN2(n72), .QN(n87) );
  NOR2X0 U21 ( .IN1(n72), .IN2(n69), .QN(n89) );
  NBUFFX2 U22 ( .INP(in1[2]), .Z(out1[25]) );
  NBUFFX2 U23 ( .INP(in1[2]), .Z(out1[26]) );
  INVX0 U24 ( .INP(in2[2]), .ZN(n3) );
  INVX0 U25 ( .INP(in2[4]), .ZN(n4) );
  INVX0 U26 ( .INP(in2[6]), .ZN(n5) );
  INVX0 U27 ( .INP(in2[8]), .ZN(n6) );
  INVX0 U28 ( .INP(in2[10]), .ZN(n7) );
  INVX0 U29 ( .INP(in2[12]), .ZN(n8) );
  INVX0 U30 ( .INP(in2[13]), .ZN(n9) );
  INVX0 U31 ( .INP(in2[14]), .ZN(n10) );
  INVX0 U32 ( .INP(in2[15]), .ZN(n11) );
  INVX0 U33 ( .INP(in2[16]), .ZN(n12) );
  INVX0 U34 ( .INP(in2[17]), .ZN(n13) );
  INVX0 U35 ( .INP(in2[18]), .ZN(n14) );
  INVX0 U36 ( .INP(in2[19]), .ZN(n15) );
  INVX0 U37 ( .INP(in2[20]), .ZN(n16) );
  INVX0 U38 ( .INP(in2[21]), .ZN(n17) );
  INVX0 U39 ( .INP(in2[22]), .ZN(n18) );
  INVX0 U40 ( .INP(in1[2]), .ZN(n69) );
  NOR2X0 U41 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n19) );
  AOI21X1 U42 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n19), .QN(n20) );
  AO222X1 U43 ( .IN1(in2[0]), .IN2(n86), .IN3(in2[1]), .IN4(n87), .IN5(n89), 
        .IN6(n20), .Q(out1[1]) );
  OR3X1 U44 ( .IN1(in2[2]), .IN2(in2[0]), .IN3(in2[1]), .Q(n21) );
  OA21X1 U45 ( .IN1(n19), .IN2(n3), .IN3(n21), .Q(n22) );
  AO222X1 U46 ( .IN1(in2[2]), .IN2(n87), .IN3(n86), .IN4(n20), .IN5(n22), 
        .IN6(n89), .Q(out1[2]) );
  NOR2X0 U47 ( .IN1(in2[3]), .IN2(n21), .QN(n23) );
  AOI21X1 U48 ( .IN1(in2[3]), .IN2(n21), .IN3(n23), .QN(n24) );
  AO222X1 U49 ( .IN1(in2[3]), .IN2(n87), .IN3(n86), .IN4(n22), .IN5(n24), 
        .IN6(n89), .Q(out1[3]) );
  OA21X1 U50 ( .IN1(n23), .IN2(n4), .IN3(n25), .Q(n26) );
  AO222X1 U51 ( .IN1(in2[4]), .IN2(n87), .IN3(n86), .IN4(n24), .IN5(n26), 
        .IN6(n89), .Q(out1[4]) );
  NOR2X0 U52 ( .IN1(in2[5]), .IN2(n25), .QN(n27) );
  AOI21X1 U53 ( .IN1(in2[5]), .IN2(n25), .IN3(n27), .QN(n28) );
  AO222X1 U54 ( .IN1(in2[5]), .IN2(n87), .IN3(n86), .IN4(n26), .IN5(n28), 
        .IN6(n89), .Q(out1[5]) );
  OA21X1 U55 ( .IN1(n27), .IN2(n5), .IN3(n29), .Q(n30) );
  AO222X1 U56 ( .IN1(in2[6]), .IN2(n87), .IN3(n86), .IN4(n28), .IN5(n30), 
        .IN6(n89), .Q(out1[6]) );
  NOR2X0 U57 ( .IN1(in2[7]), .IN2(n29), .QN(n31) );
  AOI21X1 U58 ( .IN1(in2[7]), .IN2(n29), .IN3(n31), .QN(n32) );
  AO222X1 U59 ( .IN1(in2[7]), .IN2(n87), .IN3(n86), .IN4(n30), .IN5(n32), 
        .IN6(n89), .Q(out1[7]) );
  OA21X1 U60 ( .IN1(n31), .IN2(n6), .IN3(n33), .Q(n34) );
  AO222X1 U61 ( .IN1(in2[8]), .IN2(n87), .IN3(n86), .IN4(n32), .IN5(n34), 
        .IN6(n89), .Q(out1[8]) );
  NOR2X0 U62 ( .IN1(in2[9]), .IN2(n33), .QN(n35) );
  AOI21X1 U63 ( .IN1(in2[9]), .IN2(n33), .IN3(n35), .QN(n36) );
  AO222X1 U64 ( .IN1(in2[9]), .IN2(n87), .IN3(n86), .IN4(n34), .IN5(n36), 
        .IN6(n89), .Q(out1[9]) );
  OA21X1 U65 ( .IN1(n35), .IN2(n7), .IN3(n37), .Q(n38) );
  AO222X1 U66 ( .IN1(in2[10]), .IN2(n87), .IN3(n86), .IN4(n36), .IN5(n38), 
        .IN6(n89), .Q(out1[10]) );
  NOR2X0 U67 ( .IN1(in2[11]), .IN2(n37), .QN(n39) );
  AOI21X1 U68 ( .IN1(in2[11]), .IN2(n37), .IN3(n39), .QN(n40) );
  AO222X1 U69 ( .IN1(in2[11]), .IN2(n87), .IN3(n86), .IN4(n38), .IN5(n40), 
        .IN6(n89), .Q(out1[11]) );
  OA21X1 U70 ( .IN1(n39), .IN2(n8), .IN3(n44), .Q(n42) );
  AO222X1 U71 ( .IN1(in2[12]), .IN2(n87), .IN3(n86), .IN4(n40), .IN5(n42), 
        .IN6(n89), .Q(out1[12]) );
  MUX21X1 U72 ( .IN1(n9), .IN2(in2[13]), .S(n41), .Q(n43) );
  AO22X1 U73 ( .IN1(in1[0]), .IN2(n43), .IN3(n86), .IN4(n42), .Q(out1[13]) );
  NOR2X0 U74 ( .IN1(in2[13]), .IN2(n44), .QN(n49) );
  AO21X1 U75 ( .IN1(in2[13]), .IN2(n44), .IN3(n83), .Q(n47) );
  NOR2X0 U76 ( .IN1(n49), .IN2(n69), .QN(n45) );
  MUX21X1 U77 ( .IN1(n10), .IN2(in2[14]), .S(n45), .Q(n46) );
  OAI22X1 U78 ( .IN1(n49), .IN2(n47), .IN3(n72), .IN4(n46), .QN(out1[14]) );
  MUX21X1 U79 ( .IN1(n11), .IN2(in2[15]), .S(n48), .Q(n51) );
  OA21X1 U80 ( .IN1(n49), .IN2(n10), .IN3(n86), .Q(n50) );
  AO22X1 U81 ( .IN1(in1[0]), .IN2(n51), .IN3(n50), .IN4(n52), .Q(out1[15]) );
  NOR2X0 U82 ( .IN1(in2[15]), .IN2(n52), .QN(n57) );
  AO21X1 U83 ( .IN1(in2[15]), .IN2(n52), .IN3(n83), .Q(n55) );
  NOR2X0 U84 ( .IN1(n57), .IN2(n69), .QN(n53) );
  MUX21X1 U85 ( .IN1(n12), .IN2(in2[16]), .S(n53), .Q(n54) );
  OAI22X1 U86 ( .IN1(n57), .IN2(n55), .IN3(n72), .IN4(n54), .QN(out1[16]) );
  MUX21X1 U87 ( .IN1(n13), .IN2(in2[17]), .S(n56), .Q(n59) );
  OA21X1 U88 ( .IN1(n57), .IN2(n12), .IN3(n86), .Q(n58) );
  AO22X1 U89 ( .IN1(in1[0]), .IN2(n59), .IN3(n58), .IN4(n60), .Q(out1[17]) );
  NOR2X0 U90 ( .IN1(in2[17]), .IN2(n60), .QN(n65) );
  AO21X1 U91 ( .IN1(in2[17]), .IN2(n60), .IN3(n83), .Q(n63) );
  NOR2X0 U92 ( .IN1(n65), .IN2(n69), .QN(n61) );
  MUX21X1 U93 ( .IN1(n14), .IN2(in2[18]), .S(n61), .Q(n62) );
  OAI22X1 U94 ( .IN1(n65), .IN2(n63), .IN3(n72), .IN4(n62), .QN(out1[18]) );
  MUX21X1 U95 ( .IN1(n15), .IN2(in2[19]), .S(n64), .Q(n67) );
  OA21X1 U96 ( .IN1(n65), .IN2(n14), .IN3(n86), .Q(n66) );
  AO22X1 U97 ( .IN1(in1[0]), .IN2(n67), .IN3(n66), .IN4(n68), .Q(out1[19]) );
  NOR2X0 U98 ( .IN1(in2[19]), .IN2(n68), .QN(n75) );
  AO21X1 U99 ( .IN1(in2[19]), .IN2(n68), .IN3(n83), .Q(n73) );
  NOR2X0 U100 ( .IN1(n75), .IN2(n69), .QN(n70) );
  MUX21X1 U101 ( .IN1(n16), .IN2(in2[20]), .S(n70), .Q(n71) );
  OAI22X1 U102 ( .IN1(n75), .IN2(n73), .IN3(n72), .IN4(n71), .QN(out1[20]) );
  MUX21X1 U103 ( .IN1(n17), .IN2(in2[21]), .S(n74), .Q(n77) );
  MUX21X1 U104 ( .IN1(n16), .IN2(in2[20]), .S(n75), .Q(n76) );
  AO22X1 U105 ( .IN1(in1[0]), .IN2(n77), .IN3(n86), .IN4(n76), .Q(out1[21]) );
  INVX0 U106 ( .INP(n89), .ZN(n78) );
  OR2X1 U107 ( .IN1(n79), .IN2(in2[21]), .Q(n85) );
  NOR2X0 U108 ( .IN1(n78), .IN2(n85), .QN(n84) );
  NOR2X0 U109 ( .IN1(in2[22]), .IN2(n78), .QN(n81) );
  NAND2X0 U110 ( .IN1(in2[21]), .IN2(n79), .QN(n80) );
  OA221X1 U111 ( .IN1(n81), .IN2(n86), .IN3(n81), .IN4(n80), .IN5(n85), .Q(n82) );
  AO221X1 U112 ( .IN1(in2[22]), .IN2(n87), .IN3(in2[22]), .IN4(n84), .IN5(n82), 
        .Q(out1[22]) );
  NOR2X0 U113 ( .IN1(n83), .IN2(n85), .QN(n90) );
  AO21X1 U114 ( .IN1(n86), .IN2(n85), .IN3(n84), .Q(n88) );
  AO221X1 U115 ( .IN1(in2[22]), .IN2(n90), .IN3(n18), .IN4(n88), .IN5(n87), 
        .Q(out1[23]) );
  AO21X1 U116 ( .IN1(n90), .IN2(n18), .IN3(n89), .Q(out1[24]) );
  AND2X1 U117 ( .IN1(in1[0]), .IN2(in2[0]), .Q(out1[0]) );
endmodule


module booth27_37 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n25), .IN2(n6), .QN(n30) );
  NAND2X0 U4 ( .IN1(n33), .IN2(n7), .QN(n37) );
  NAND2X0 U5 ( .IN1(n41), .IN2(n8), .QN(n45) );
  NAND2X0 U6 ( .IN1(n49), .IN2(n9), .QN(n53) );
  NAND2X0 U7 ( .IN1(n57), .IN2(n10), .QN(n61) );
  NAND2X0 U8 ( .IN1(n118), .IN2(n19), .QN(n125) );
  NAND2X0 U9 ( .IN1(n65), .IN2(n11), .QN(n77) );
  NAND2X0 U10 ( .IN1(n81), .IN2(n13), .QN(n89) );
  NAND2X0 U11 ( .IN1(n105), .IN2(n17), .QN(n114) );
  NAND2X0 U12 ( .IN1(n93), .IN2(n15), .QN(n101) );
  NAND2X0 U13 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U14 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U15 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U16 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U17 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U18 ( .IN1(n27), .IN2(n132), .QN(n4) );
  NAND2X0 U19 ( .IN1(n141), .IN2(n130), .QN(n24) );
  NAND2X0 U20 ( .IN1(n32), .IN2(n31), .QN(out1[3]) );
  NAND2X0 U21 ( .IN1(n36), .IN2(n35), .QN(out1[4]) );
  NAND2X0 U22 ( .IN1(in1[2]), .IN2(n77), .QN(n71) );
  NAND2X0 U23 ( .IN1(n70), .IN2(n132), .QN(n74) );
  NAND2X0 U24 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U25 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U26 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U27 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U28 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NAND2X0 U29 ( .IN1(n40), .IN2(n39), .QN(out1[5]) );
  NAND2X0 U30 ( .IN1(n44), .IN2(n43), .QN(out1[6]) );
  NAND2X0 U31 ( .IN1(n48), .IN2(n47), .QN(out1[7]) );
  NAND2X0 U32 ( .IN1(n52), .IN2(n51), .QN(out1[8]) );
  NAND2X0 U33 ( .IN1(n56), .IN2(n55), .QN(out1[9]) );
  NAND2X0 U34 ( .IN1(n60), .IN2(n59), .QN(out1[10]) );
  NAND2X0 U35 ( .IN1(n64), .IN2(n63), .QN(out1[11]) );
  NAND2X0 U36 ( .IN1(n69), .IN2(n68), .QN(out1[12]) );
  NAND2X0 U37 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U38 ( .IN1(n23), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U39 ( .IN1(in1[2]), .IN2(n22), .QN(n23) );
  NOR2X0 U40 ( .IN1(n28), .IN2(n26), .QN(n3) );
  NOR2X0 U41 ( .IN1(n142), .IN2(n21), .QN(n1) );
  INVX0 U42 ( .INP(n130), .ZN(n137) );
  INVX0 U43 ( .INP(n132), .ZN(n141) );
  NOR3X0 U44 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  NAND3X0 U45 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  NOR2X0 U46 ( .IN1(n142), .IN2(n111), .QN(n138) );
  MUX21X1 U47 ( .IN1(n22), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  INVX0 U48 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U49 ( .INP(in2[2]), .ZN(n6) );
  INVX0 U50 ( .INP(in2[4]), .ZN(n7) );
  INVX0 U51 ( .INP(in2[6]), .ZN(n8) );
  INVX0 U52 ( .INP(in2[8]), .ZN(n9) );
  INVX0 U53 ( .INP(in2[10]), .ZN(n10) );
  INVX0 U54 ( .INP(in2[12]), .ZN(n11) );
  INVX0 U55 ( .INP(in2[13]), .ZN(n12) );
  INVX0 U56 ( .INP(in2[14]), .ZN(n13) );
  INVX0 U57 ( .INP(in2[15]), .ZN(n14) );
  INVX0 U58 ( .INP(in2[16]), .ZN(n15) );
  INVX0 U59 ( .INP(in2[17]), .ZN(n16) );
  INVX0 U60 ( .INP(in2[18]), .ZN(n17) );
  INVX0 U61 ( .INP(in2[19]), .ZN(n18) );
  INVX0 U62 ( .INP(in2[20]), .ZN(n19) );
  INVX0 U63 ( .INP(in2[21]), .ZN(n20) );
  INVX0 U64 ( .INP(in2[22]), .ZN(n21) );
  INVX0 U65 ( .INP(in1[1]), .ZN(n22) );
  INVX0 U66 ( .INP(in1[2]), .ZN(n111) );
  INVX0 U67 ( .INP(n138), .ZN(n140) );
  NOR2X0 U68 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n25) );
  AOI21X1 U69 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n25), .QN(n27) );
  NOR2X0 U70 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U71 ( .IN1(n24), .IN2(in2[0]), .IN3(n138), .IN4(n27), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U72 ( .INP(n133), .ZN(n67) );
  NOR2X0 U73 ( .IN1(n67), .IN2(n6), .QN(n28) );
  OA21X1 U74 ( .IN1(n25), .IN2(n6), .IN3(n30), .Q(n29) );
  AO22X1 U75 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n29), .Q(n26) );
  AOI22X1 U76 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n29), .QN(n32) );
  NOR2X0 U77 ( .IN1(in2[3]), .IN2(n30), .QN(n33) );
  AO21X1 U78 ( .IN1(in2[3]), .IN2(n30), .IN3(n33), .Q(n34) );
  OA22X1 U79 ( .IN1(n6), .IN2(n130), .IN3(n140), .IN4(n34), .Q(n31) );
  OA21X1 U80 ( .IN1(n33), .IN2(n7), .IN3(n37), .Q(n38) );
  AOI22X1 U81 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n38), .QN(n36) );
  OA22X1 U82 ( .IN1(n67), .IN2(n7), .IN3(n141), .IN4(n34), .Q(n35) );
  NOR2X0 U83 ( .IN1(in2[5]), .IN2(n37), .QN(n41) );
  AO21X1 U84 ( .IN1(in2[5]), .IN2(n37), .IN3(n41), .Q(n42) );
  OA22X1 U85 ( .IN1(n7), .IN2(n130), .IN3(n140), .IN4(n42), .Q(n40) );
  AOI22X1 U86 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n38), .QN(n39) );
  OA21X1 U87 ( .IN1(n41), .IN2(n8), .IN3(n45), .Q(n46) );
  AOI22X1 U88 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n46), .QN(n44) );
  OA22X1 U89 ( .IN1(n67), .IN2(n8), .IN3(n141), .IN4(n42), .Q(n43) );
  NOR2X0 U90 ( .IN1(in2[7]), .IN2(n45), .QN(n49) );
  AO21X1 U91 ( .IN1(in2[7]), .IN2(n45), .IN3(n49), .Q(n50) );
  OA22X1 U92 ( .IN1(n8), .IN2(n130), .IN3(n140), .IN4(n50), .Q(n48) );
  AOI22X1 U93 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n46), .QN(n47) );
  OA21X1 U94 ( .IN1(n49), .IN2(n9), .IN3(n53), .Q(n54) );
  AOI22X1 U95 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n54), .QN(n52) );
  OA22X1 U96 ( .IN1(n67), .IN2(n9), .IN3(n141), .IN4(n50), .Q(n51) );
  NOR2X0 U97 ( .IN1(in2[9]), .IN2(n53), .QN(n57) );
  AO21X1 U98 ( .IN1(in2[9]), .IN2(n53), .IN3(n57), .Q(n58) );
  OA22X1 U99 ( .IN1(n9), .IN2(n130), .IN3(n140), .IN4(n58), .Q(n56) );
  AOI22X1 U100 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n54), .QN(n55) );
  OA21X1 U101 ( .IN1(n57), .IN2(n10), .IN3(n61), .Q(n62) );
  AOI22X1 U102 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n62), .QN(n60) );
  OA22X1 U103 ( .IN1(n67), .IN2(n10), .IN3(n141), .IN4(n58), .Q(n59) );
  NOR2X0 U104 ( .IN1(in2[11]), .IN2(n61), .QN(n65) );
  AO21X1 U105 ( .IN1(in2[11]), .IN2(n61), .IN3(n65), .Q(n66) );
  OA22X1 U106 ( .IN1(n10), .IN2(n130), .IN3(n140), .IN4(n66), .Q(n64) );
  AOI22X1 U107 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n62), .QN(n63) );
  OA21X1 U108 ( .IN1(n65), .IN2(n11), .IN3(n77), .Q(n70) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n70), .QN(n69) );
  OA22X1 U110 ( .IN1(n67), .IN2(n11), .IN3(n141), .IN4(n66), .Q(n68) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n12), .S(n71), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n11), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n13), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n12), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n12), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n14), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n13), .IN4(n85), .IN5(n84), 
        .Q(out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n15), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n14), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n14), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n16), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n15), .IN4(n97), .IN5(n96), 
        .Q(out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n17), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n16), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n16), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n18), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n17), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n19), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n18), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n18), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n20), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n19), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n21), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n20), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n20), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n21), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_38 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X0 U3 ( .IN1(n33), .IN2(n7), .QN(n37) );
  NAND2X0 U4 ( .IN1(n41), .IN2(n8), .QN(n45) );
  NAND2X0 U5 ( .IN1(n49), .IN2(n9), .QN(n53) );
  NAND2X0 U6 ( .IN1(n57), .IN2(n10), .QN(n61) );
  NAND2X0 U7 ( .IN1(n25), .IN2(n6), .QN(n30) );
  NAND2X0 U8 ( .IN1(n65), .IN2(n11), .QN(n77) );
  NAND2X0 U9 ( .IN1(n81), .IN2(n13), .QN(n89) );
  NAND2X0 U10 ( .IN1(n93), .IN2(n15), .QN(n101) );
  NAND2X0 U11 ( .IN1(n118), .IN2(n19), .QN(n125) );
  NAND2X0 U12 ( .IN1(n105), .IN2(n17), .QN(n114) );
  NAND2X0 U13 ( .IN1(n1), .IN2(n2), .QN(n129) );
  NAND2X0 U14 ( .IN1(in1[2]), .IN2(n124), .QN(n2) );
  NAND2X0 U15 ( .IN1(n136), .IN2(n130), .QN(n135) );
  NAND2X0 U16 ( .IN1(n132), .IN2(n131), .QN(n136) );
  NAND2X0 U17 ( .IN1(n40), .IN2(n39), .QN(out1[5]) );
  NAND2X0 U18 ( .IN1(n44), .IN2(n43), .QN(out1[6]) );
  NAND2X0 U19 ( .IN1(in1[2]), .IN2(n77), .QN(n71) );
  NAND2X0 U20 ( .IN1(n70), .IN2(n132), .QN(n74) );
  NAND2X0 U21 ( .IN1(in1[2]), .IN2(n89), .QN(n82) );
  NAND2X0 U22 ( .IN1(in1[2]), .IN2(n101), .QN(n94) );
  NAND2X0 U23 ( .IN1(in1[2]), .IN2(n114), .QN(n106) );
  NAND2X0 U24 ( .IN1(in1[2]), .IN2(n125), .QN(n119) );
  NAND2X0 U25 ( .IN1(n141), .IN2(n140), .QN(out1[25]) );
  NAND2X0 U26 ( .IN1(n23), .IN2(n140), .QN(out1[26]) );
  NAND2X0 U27 ( .IN1(in1[2]), .IN2(n22), .QN(n23) );
  NAND2X0 U28 ( .IN1(n36), .IN2(n35), .QN(out1[4]) );
  NAND2X0 U29 ( .IN1(n32), .IN2(n31), .QN(out1[3]) );
  NAND2X0 U30 ( .IN1(n27), .IN2(n132), .QN(n4) );
  NAND2X0 U31 ( .IN1(n48), .IN2(n47), .QN(out1[7]) );
  NAND2X0 U32 ( .IN1(n52), .IN2(n51), .QN(out1[8]) );
  NAND2X0 U33 ( .IN1(n56), .IN2(n55), .QN(out1[9]) );
  NAND2X0 U34 ( .IN1(n60), .IN2(n59), .QN(out1[10]) );
  NAND2X0 U35 ( .IN1(n64), .IN2(n63), .QN(out1[11]) );
  NAND2X0 U36 ( .IN1(n69), .IN2(n68), .QN(out1[12]) );
  NAND2X0 U37 ( .IN1(n74), .IN2(n73), .QN(out1[13]) );
  NAND2X0 U38 ( .IN1(n141), .IN2(n130), .QN(n24) );
  NAND2X0 U39 ( .IN1(n3), .IN2(n4), .QN(out1[2]) );
  NOR2X0 U40 ( .IN1(n28), .IN2(n26), .QN(n3) );
  INVX0 U41 ( .INP(n130), .ZN(n137) );
  INVX0 U42 ( .INP(n132), .ZN(n141) );
  NOR3X0 U43 ( .IN1(in1[0]), .IN2(in1[1]), .IN3(n111), .QN(n132) );
  NAND3X0 U44 ( .IN1(in1[1]), .IN2(in1[0]), .IN3(n111), .QN(n130) );
  NOR2X0 U45 ( .IN1(n142), .IN2(n111), .QN(n138) );
  NOR2X0 U46 ( .IN1(n142), .IN2(n21), .QN(n1) );
  MUX21X1 U47 ( .IN1(n22), .IN2(in1[1]), .S(in1[0]), .Q(n142) );
  INVX0 U48 ( .INP(in2[0]), .ZN(n5) );
  INVX0 U49 ( .INP(in2[2]), .ZN(n6) );
  INVX0 U50 ( .INP(in2[4]), .ZN(n7) );
  INVX0 U51 ( .INP(in2[6]), .ZN(n8) );
  INVX0 U52 ( .INP(in2[8]), .ZN(n9) );
  INVX0 U53 ( .INP(in2[10]), .ZN(n10) );
  INVX0 U54 ( .INP(in2[12]), .ZN(n11) );
  INVX0 U55 ( .INP(in2[13]), .ZN(n12) );
  INVX0 U56 ( .INP(in2[14]), .ZN(n13) );
  INVX0 U57 ( .INP(in2[15]), .ZN(n14) );
  INVX0 U58 ( .INP(in2[16]), .ZN(n15) );
  INVX0 U59 ( .INP(in2[17]), .ZN(n16) );
  INVX0 U60 ( .INP(in2[18]), .ZN(n17) );
  INVX0 U61 ( .INP(in2[19]), .ZN(n18) );
  INVX0 U62 ( .INP(in2[20]), .ZN(n19) );
  INVX0 U63 ( .INP(in2[21]), .ZN(n20) );
  INVX0 U64 ( .INP(in2[22]), .ZN(n21) );
  INVX0 U65 ( .INP(in1[1]), .ZN(n22) );
  INVX0 U66 ( .INP(in1[2]), .ZN(n111) );
  INVX0 U67 ( .INP(n138), .ZN(n140) );
  NOR2X0 U68 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n25) );
  AOI21X1 U69 ( .IN1(in2[1]), .IN2(in2[0]), .IN3(n25), .QN(n27) );
  NOR2X0 U70 ( .IN1(n142), .IN2(in1[2]), .QN(n133) );
  AO222X1 U71 ( .IN1(n24), .IN2(in2[0]), .IN3(n138), .IN4(n27), .IN5(n133), 
        .IN6(in2[1]), .Q(out1[1]) );
  INVX0 U72 ( .INP(n133), .ZN(n67) );
  NOR2X0 U73 ( .IN1(n67), .IN2(n6), .QN(n28) );
  OA21X1 U74 ( .IN1(n25), .IN2(n6), .IN3(n30), .Q(n29) );
  AO22X1 U75 ( .IN1(in2[1]), .IN2(n137), .IN3(n138), .IN4(n29), .Q(n26) );
  AOI22X1 U76 ( .IN1(n133), .IN2(in2[3]), .IN3(n132), .IN4(n29), .QN(n32) );
  NOR2X0 U77 ( .IN1(in2[3]), .IN2(n30), .QN(n33) );
  AO21X1 U78 ( .IN1(in2[3]), .IN2(n30), .IN3(n33), .Q(n34) );
  OA22X1 U79 ( .IN1(n6), .IN2(n130), .IN3(n140), .IN4(n34), .Q(n31) );
  OA21X1 U80 ( .IN1(n33), .IN2(n7), .IN3(n37), .Q(n38) );
  AOI22X1 U81 ( .IN1(in2[3]), .IN2(n137), .IN3(n138), .IN4(n38), .QN(n36) );
  OA22X1 U82 ( .IN1(n67), .IN2(n7), .IN3(n141), .IN4(n34), .Q(n35) );
  NOR2X0 U83 ( .IN1(in2[5]), .IN2(n37), .QN(n41) );
  AO21X1 U84 ( .IN1(in2[5]), .IN2(n37), .IN3(n41), .Q(n42) );
  OA22X1 U85 ( .IN1(n7), .IN2(n130), .IN3(n140), .IN4(n42), .Q(n40) );
  AOI22X1 U86 ( .IN1(n133), .IN2(in2[5]), .IN3(n132), .IN4(n38), .QN(n39) );
  OA21X1 U87 ( .IN1(n41), .IN2(n8), .IN3(n45), .Q(n46) );
  AOI22X1 U88 ( .IN1(in2[5]), .IN2(n137), .IN3(n138), .IN4(n46), .QN(n44) );
  OA22X1 U89 ( .IN1(n67), .IN2(n8), .IN3(n141), .IN4(n42), .Q(n43) );
  NOR2X0 U90 ( .IN1(in2[7]), .IN2(n45), .QN(n49) );
  AO21X1 U91 ( .IN1(in2[7]), .IN2(n45), .IN3(n49), .Q(n50) );
  OA22X1 U92 ( .IN1(n8), .IN2(n130), .IN3(n140), .IN4(n50), .Q(n48) );
  AOI22X1 U93 ( .IN1(n133), .IN2(in2[7]), .IN3(n132), .IN4(n46), .QN(n47) );
  OA21X1 U94 ( .IN1(n49), .IN2(n9), .IN3(n53), .Q(n54) );
  AOI22X1 U95 ( .IN1(in2[7]), .IN2(n137), .IN3(n138), .IN4(n54), .QN(n52) );
  OA22X1 U96 ( .IN1(n67), .IN2(n9), .IN3(n141), .IN4(n50), .Q(n51) );
  NOR2X0 U97 ( .IN1(in2[9]), .IN2(n53), .QN(n57) );
  AO21X1 U98 ( .IN1(in2[9]), .IN2(n53), .IN3(n57), .Q(n58) );
  OA22X1 U99 ( .IN1(n9), .IN2(n130), .IN3(n140), .IN4(n58), .Q(n56) );
  AOI22X1 U100 ( .IN1(n133), .IN2(in2[9]), .IN3(n132), .IN4(n54), .QN(n55) );
  OA21X1 U101 ( .IN1(n57), .IN2(n10), .IN3(n61), .Q(n62) );
  AOI22X1 U102 ( .IN1(in2[9]), .IN2(n137), .IN3(n138), .IN4(n62), .QN(n60) );
  OA22X1 U103 ( .IN1(n67), .IN2(n10), .IN3(n141), .IN4(n58), .Q(n59) );
  NOR2X0 U104 ( .IN1(in2[11]), .IN2(n61), .QN(n65) );
  AO21X1 U105 ( .IN1(in2[11]), .IN2(n61), .IN3(n65), .Q(n66) );
  OA22X1 U106 ( .IN1(n10), .IN2(n130), .IN3(n140), .IN4(n66), .Q(n64) );
  AOI22X1 U107 ( .IN1(n133), .IN2(in2[11]), .IN3(n132), .IN4(n62), .QN(n63) );
  OA21X1 U108 ( .IN1(n65), .IN2(n11), .IN3(n77), .Q(n70) );
  AOI22X1 U109 ( .IN1(in2[11]), .IN2(n137), .IN3(n138), .IN4(n70), .QN(n69) );
  OA22X1 U110 ( .IN1(n67), .IN2(n11), .IN3(n141), .IN4(n66), .Q(n68) );
  MUX21X1 U111 ( .IN1(in2[13]), .IN2(n12), .S(n71), .Q(n72) );
  OA22X1 U112 ( .IN1(n142), .IN2(n72), .IN3(n130), .IN4(n11), .Q(n73) );
  NOR2X0 U113 ( .IN1(in2[13]), .IN2(n77), .QN(n81) );
  NOR2X0 U114 ( .IN1(n81), .IN2(n111), .QN(n76) );
  INVX0 U115 ( .INP(n76), .ZN(n75) );
  AO221X1 U116 ( .IN1(in2[14]), .IN2(n76), .IN3(n13), .IN4(n75), .IN5(n142), 
        .Q(n80) );
  AO221X1 U117 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n77), .IN5(n12), .Q(
        n79) );
  NAND3X0 U118 ( .IN1(n132), .IN2(n12), .IN3(n77), .QN(n78) );
  NAND3X0 U119 ( .IN1(n80), .IN2(n79), .IN3(n78), .QN(out1[14]) );
  AO21X1 U120 ( .IN1(n81), .IN2(n132), .IN3(n137), .Q(n86) );
  NOR2X0 U121 ( .IN1(n81), .IN2(n141), .QN(n85) );
  MUX21X1 U122 ( .IN1(in2[15]), .IN2(n14), .S(n82), .Q(n83) );
  NOR2X0 U123 ( .IN1(n142), .IN2(n83), .QN(n84) );
  AO221X1 U124 ( .IN1(in2[14]), .IN2(n86), .IN3(n13), .IN4(n85), .IN5(n84), 
        .Q(out1[15]) );
  NOR2X0 U125 ( .IN1(in2[15]), .IN2(n89), .QN(n93) );
  NOR2X0 U126 ( .IN1(n93), .IN2(n111), .QN(n88) );
  INVX0 U127 ( .INP(n88), .ZN(n87) );
  AO221X1 U128 ( .IN1(in2[16]), .IN2(n88), .IN3(n15), .IN4(n87), .IN5(n142), 
        .Q(n92) );
  AO221X1 U129 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n89), .IN5(n14), .Q(
        n91) );
  NAND3X0 U130 ( .IN1(n132), .IN2(n14), .IN3(n89), .QN(n90) );
  NAND3X0 U131 ( .IN1(n92), .IN2(n91), .IN3(n90), .QN(out1[16]) );
  AO21X1 U132 ( .IN1(n93), .IN2(n132), .IN3(n137), .Q(n98) );
  NOR2X0 U133 ( .IN1(n93), .IN2(n141), .QN(n97) );
  MUX21X1 U134 ( .IN1(in2[17]), .IN2(n16), .S(n94), .Q(n95) );
  NOR2X0 U135 ( .IN1(n142), .IN2(n95), .QN(n96) );
  AO221X1 U136 ( .IN1(in2[16]), .IN2(n98), .IN3(n15), .IN4(n97), .IN5(n96), 
        .Q(out1[17]) );
  NOR2X0 U137 ( .IN1(in2[17]), .IN2(n101), .QN(n105) );
  NOR2X0 U138 ( .IN1(n105), .IN2(n111), .QN(n100) );
  INVX0 U139 ( .INP(n100), .ZN(n99) );
  AO221X1 U140 ( .IN1(in2[18]), .IN2(n100), .IN3(n17), .IN4(n99), .IN5(n142), 
        .Q(n104) );
  AO221X1 U141 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n101), .IN5(n16), 
        .Q(n103) );
  NAND3X0 U142 ( .IN1(n132), .IN2(n16), .IN3(n101), .QN(n102) );
  NAND3X0 U143 ( .IN1(n104), .IN2(n103), .IN3(n102), .QN(out1[18]) );
  AO21X1 U144 ( .IN1(n105), .IN2(n132), .IN3(n137), .Q(n110) );
  NOR2X0 U145 ( .IN1(n105), .IN2(n141), .QN(n109) );
  MUX21X1 U146 ( .IN1(in2[19]), .IN2(n18), .S(n106), .Q(n107) );
  NOR2X0 U147 ( .IN1(n142), .IN2(n107), .QN(n108) );
  AO221X1 U148 ( .IN1(in2[18]), .IN2(n110), .IN3(n17), .IN4(n109), .IN5(n108), 
        .Q(out1[19]) );
  NOR2X0 U149 ( .IN1(in2[19]), .IN2(n114), .QN(n118) );
  NOR2X0 U150 ( .IN1(n118), .IN2(n111), .QN(n113) );
  INVX0 U151 ( .INP(n113), .ZN(n112) );
  AO221X1 U152 ( .IN1(in2[20]), .IN2(n113), .IN3(n19), .IN4(n112), .IN5(n142), 
        .Q(n117) );
  AO221X1 U153 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n114), .IN5(n18), 
        .Q(n116) );
  NAND3X0 U154 ( .IN1(n132), .IN2(n18), .IN3(n114), .QN(n115) );
  NAND3X0 U155 ( .IN1(n117), .IN2(n116), .IN3(n115), .QN(out1[20]) );
  AO21X1 U156 ( .IN1(n118), .IN2(n132), .IN3(n137), .Q(n123) );
  NOR2X0 U157 ( .IN1(n118), .IN2(n141), .QN(n122) );
  MUX21X1 U158 ( .IN1(in2[21]), .IN2(n20), .S(n119), .Q(n120) );
  NOR2X0 U159 ( .IN1(n142), .IN2(n120), .QN(n121) );
  AO221X1 U160 ( .IN1(in2[20]), .IN2(n123), .IN3(n19), .IN4(n122), .IN5(n121), 
        .Q(out1[21]) );
  NOR2X0 U161 ( .IN1(in2[21]), .IN2(n125), .QN(n131) );
  INVX0 U162 ( .INP(n131), .ZN(n124) );
  NAND3X0 U163 ( .IN1(n138), .IN2(n21), .IN3(n124), .QN(n128) );
  AO221X1 U164 ( .IN1(n130), .IN2(n141), .IN3(n130), .IN4(n125), .IN5(n20), 
        .Q(n127) );
  NAND3X0 U165 ( .IN1(n132), .IN2(n20), .IN3(n125), .QN(n126) );
  NAND4X0 U166 ( .IN1(n129), .IN2(n128), .IN3(n127), .IN4(n126), .QN(out1[22])
         );
  MUX21X1 U167 ( .IN1(n132), .IN2(n138), .S(n131), .Q(n134) );
  AO221X1 U168 ( .IN1(in2[22]), .IN2(n135), .IN3(n21), .IN4(n134), .IN5(n133), 
        .Q(out1[23]) );
  NOR2X0 U169 ( .IN1(in2[22]), .IN2(n136), .QN(n139) );
  OR3X1 U170 ( .IN1(n139), .IN2(n138), .IN3(n137), .Q(out1[24]) );
  NOR2X0 U171 ( .IN1(n142), .IN2(n5), .QN(out1[0]) );
endmodule


module booth27_39 ( out1, in1, in2 );
  output [26:0] out1;
  input [2:0] in1;
  input [25:0] in2;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93;

  NAND2X0 U3 ( .IN1(n30), .IN2(n7), .QN(n32) );
  NAND2X0 U4 ( .IN1(n34), .IN2(n8), .QN(n36) );
  NAND2X0 U5 ( .IN1(n38), .IN2(n9), .QN(n40) );
  NAND2X0 U6 ( .IN1(n42), .IN2(n10), .QN(n47) );
  NAND2X0 U7 ( .IN1(n78), .IN2(n18), .QN(n82) );
  NAND2X0 U8 ( .IN1(n26), .IN2(n6), .QN(n28) );
  NAND2X0 U9 ( .IN1(in1[2]), .IN2(n47), .QN(n44) );
  NAND2X0 U10 ( .IN1(n52), .IN2(n12), .QN(n55) );
  NAND2X0 U11 ( .IN1(in1[2]), .IN2(n55), .QN(n51) );
  NAND2X0 U12 ( .IN1(n60), .IN2(n14), .QN(n63) );
  NAND2X0 U13 ( .IN1(in1[2]), .IN2(n63), .QN(n59) );
  NAND2X0 U14 ( .IN1(n68), .IN2(n16), .QN(n71) );
  NAND2X0 U15 ( .IN1(in1[2]), .IN2(n71), .QN(n67) );
  NAND2X0 U16 ( .IN1(in1[2]), .IN2(n82), .QN(n77) );
  NAND2X0 U17 ( .IN1(n75), .IN2(in1[2]), .QN(n86) );
  NAND2X0 U18 ( .IN1(n3), .IN2(n4), .QN(n22) );
  NAND2X0 U19 ( .IN1(in2[1]), .IN2(in2[0]), .QN(n4) );
  NAND2X0 U20 ( .IN1(n23), .IN2(n22), .QN(out1[2]) );
  INVX0 U21 ( .INP(n86), .ZN(n89) );
  NOR2X0 U22 ( .IN1(n21), .IN2(n86), .QN(n3) );
  NOR2X0 U23 ( .IN1(in1[2]), .IN2(n75), .QN(n90) );
  NOR2X0 U24 ( .IN1(n75), .IN2(n72), .QN(n92) );
  NBUFFX2 U25 ( .INP(in1[2]), .Z(out1[26]) );
  NBUFFX2 U26 ( .INP(in1[2]), .Z(out1[25]) );
  INVX0 U27 ( .INP(in2[2]), .ZN(n5) );
  INVX0 U28 ( .INP(in2[4]), .ZN(n6) );
  INVX0 U29 ( .INP(in2[6]), .ZN(n7) );
  INVX0 U30 ( .INP(in2[8]), .ZN(n8) );
  INVX0 U31 ( .INP(in2[10]), .ZN(n9) );
  INVX0 U32 ( .INP(in2[12]), .ZN(n10) );
  INVX0 U33 ( .INP(in2[13]), .ZN(n11) );
  INVX0 U34 ( .INP(in2[14]), .ZN(n12) );
  INVX0 U35 ( .INP(in2[15]), .ZN(n13) );
  INVX0 U36 ( .INP(in2[16]), .ZN(n14) );
  INVX0 U37 ( .INP(in2[17]), .ZN(n15) );
  INVX0 U38 ( .INP(in2[18]), .ZN(n16) );
  INVX0 U39 ( .INP(in2[19]), .ZN(n17) );
  INVX0 U40 ( .INP(in2[20]), .ZN(n18) );
  INVX0 U41 ( .INP(in2[21]), .ZN(n19) );
  INVX0 U42 ( .INP(in2[22]), .ZN(n20) );
  INVX0 U43 ( .INP(in1[1]), .ZN(n75) );
  INVX0 U44 ( .INP(in1[2]), .ZN(n72) );
  NOR2X0 U45 ( .IN1(in2[0]), .IN2(in2[1]), .QN(n21) );
  OR3X1 U46 ( .IN1(in2[2]), .IN2(in2[0]), .IN3(in2[1]), .Q(n24) );
  OA21X1 U47 ( .IN1(n21), .IN2(n5), .IN3(n24), .Q(n25) );
  AOI22X1 U48 ( .IN1(in2[2]), .IN2(n90), .IN3(n92), .IN4(n25), .QN(n23) );
  NOR2X0 U49 ( .IN1(in2[3]), .IN2(n24), .QN(n26) );
  AOI21X1 U50 ( .IN1(in2[3]), .IN2(n24), .IN3(n26), .QN(n27) );
  AO222X1 U51 ( .IN1(in2[3]), .IN2(n90), .IN3(n92), .IN4(n27), .IN5(n89), 
        .IN6(n25), .Q(out1[3]) );
  OA21X1 U52 ( .IN1(n26), .IN2(n6), .IN3(n28), .Q(n29) );
  AO222X1 U53 ( .IN1(in2[4]), .IN2(n90), .IN3(n92), .IN4(n29), .IN5(n89), 
        .IN6(n27), .Q(out1[4]) );
  NOR2X0 U54 ( .IN1(in2[5]), .IN2(n28), .QN(n30) );
  AOI21X1 U55 ( .IN1(in2[5]), .IN2(n28), .IN3(n30), .QN(n31) );
  AO222X1 U56 ( .IN1(in2[5]), .IN2(n90), .IN3(n92), .IN4(n31), .IN5(n89), 
        .IN6(n29), .Q(out1[5]) );
  OA21X1 U57 ( .IN1(n30), .IN2(n7), .IN3(n32), .Q(n33) );
  AO222X1 U58 ( .IN1(in2[6]), .IN2(n90), .IN3(n92), .IN4(n33), .IN5(n89), 
        .IN6(n31), .Q(out1[6]) );
  NOR2X0 U59 ( .IN1(in2[7]), .IN2(n32), .QN(n34) );
  AOI21X1 U60 ( .IN1(in2[7]), .IN2(n32), .IN3(n34), .QN(n35) );
  AO222X1 U61 ( .IN1(in2[7]), .IN2(n90), .IN3(n92), .IN4(n35), .IN5(n89), 
        .IN6(n33), .Q(out1[7]) );
  OA21X1 U62 ( .IN1(n34), .IN2(n8), .IN3(n36), .Q(n37) );
  AO222X1 U63 ( .IN1(in2[8]), .IN2(n90), .IN3(n92), .IN4(n37), .IN5(n89), 
        .IN6(n35), .Q(out1[8]) );
  NOR2X0 U64 ( .IN1(in2[9]), .IN2(n36), .QN(n38) );
  AOI21X1 U65 ( .IN1(in2[9]), .IN2(n36), .IN3(n38), .QN(n39) );
  AO222X1 U66 ( .IN1(in2[9]), .IN2(n90), .IN3(n92), .IN4(n39), .IN5(n89), 
        .IN6(n37), .Q(out1[9]) );
  OA21X1 U67 ( .IN1(n38), .IN2(n9), .IN3(n40), .Q(n41) );
  AO222X1 U68 ( .IN1(in2[10]), .IN2(n90), .IN3(n92), .IN4(n41), .IN5(n89), 
        .IN6(n39), .Q(out1[10]) );
  NOR2X0 U69 ( .IN1(in2[11]), .IN2(n40), .QN(n42) );
  AOI21X1 U70 ( .IN1(in2[11]), .IN2(n40), .IN3(n42), .QN(n43) );
  AO222X1 U71 ( .IN1(in2[11]), .IN2(n90), .IN3(n92), .IN4(n43), .IN5(n89), 
        .IN6(n41), .Q(out1[11]) );
  OA21X1 U72 ( .IN1(n42), .IN2(n10), .IN3(n47), .Q(n45) );
  AO222X1 U73 ( .IN1(in2[12]), .IN2(n90), .IN3(n92), .IN4(n45), .IN5(n89), 
        .IN6(n43), .Q(out1[12]) );
  MUX21X1 U74 ( .IN1(n11), .IN2(in2[13]), .S(n44), .Q(n46) );
  AO22X1 U75 ( .IN1(in1[1]), .IN2(n46), .IN3(n89), .IN4(n45), .Q(out1[13]) );
  NOR2X0 U76 ( .IN1(in2[13]), .IN2(n47), .QN(n52) );
  AO21X1 U77 ( .IN1(in2[13]), .IN2(n47), .IN3(n86), .Q(n50) );
  NOR2X0 U78 ( .IN1(n52), .IN2(n72), .QN(n48) );
  MUX21X1 U79 ( .IN1(n12), .IN2(in2[14]), .S(n48), .Q(n49) );
  OAI22X1 U80 ( .IN1(n52), .IN2(n50), .IN3(n75), .IN4(n49), .QN(out1[14]) );
  MUX21X1 U81 ( .IN1(n13), .IN2(in2[15]), .S(n51), .Q(n54) );
  OA21X1 U82 ( .IN1(n52), .IN2(n12), .IN3(n89), .Q(n53) );
  AO22X1 U83 ( .IN1(in1[1]), .IN2(n54), .IN3(n53), .IN4(n55), .Q(out1[15]) );
  NOR2X0 U84 ( .IN1(in2[15]), .IN2(n55), .QN(n60) );
  AO21X1 U85 ( .IN1(in2[15]), .IN2(n55), .IN3(n86), .Q(n58) );
  NOR2X0 U86 ( .IN1(n60), .IN2(n72), .QN(n56) );
  MUX21X1 U87 ( .IN1(n14), .IN2(in2[16]), .S(n56), .Q(n57) );
  OAI22X1 U88 ( .IN1(n60), .IN2(n58), .IN3(n75), .IN4(n57), .QN(out1[16]) );
  MUX21X1 U89 ( .IN1(n15), .IN2(in2[17]), .S(n59), .Q(n62) );
  OA21X1 U90 ( .IN1(n60), .IN2(n14), .IN3(n89), .Q(n61) );
  AO22X1 U91 ( .IN1(in1[1]), .IN2(n62), .IN3(n61), .IN4(n63), .Q(out1[17]) );
  NOR2X0 U92 ( .IN1(in2[17]), .IN2(n63), .QN(n68) );
  AO21X1 U93 ( .IN1(in2[17]), .IN2(n63), .IN3(n86), .Q(n66) );
  NOR2X0 U94 ( .IN1(n68), .IN2(n72), .QN(n64) );
  MUX21X1 U95 ( .IN1(n16), .IN2(in2[18]), .S(n64), .Q(n65) );
  OAI22X1 U96 ( .IN1(n68), .IN2(n66), .IN3(n75), .IN4(n65), .QN(out1[18]) );
  MUX21X1 U97 ( .IN1(n17), .IN2(in2[19]), .S(n67), .Q(n70) );
  OA21X1 U98 ( .IN1(n68), .IN2(n16), .IN3(n89), .Q(n69) );
  AO22X1 U99 ( .IN1(in1[1]), .IN2(n70), .IN3(n69), .IN4(n71), .Q(out1[19]) );
  NOR2X0 U100 ( .IN1(in2[19]), .IN2(n71), .QN(n78) );
  AO21X1 U101 ( .IN1(in2[19]), .IN2(n71), .IN3(n86), .Q(n76) );
  NOR2X0 U102 ( .IN1(n78), .IN2(n72), .QN(n73) );
  MUX21X1 U103 ( .IN1(n18), .IN2(in2[20]), .S(n73), .Q(n74) );
  OAI22X1 U104 ( .IN1(n78), .IN2(n76), .IN3(n75), .IN4(n74), .QN(out1[20]) );
  MUX21X1 U105 ( .IN1(n19), .IN2(in2[21]), .S(n77), .Q(n80) );
  MUX21X1 U106 ( .IN1(n18), .IN2(in2[20]), .S(n78), .Q(n79) );
  AO22X1 U107 ( .IN1(in1[1]), .IN2(n80), .IN3(n89), .IN4(n79), .Q(out1[21]) );
  INVX0 U108 ( .INP(n92), .ZN(n81) );
  OR2X1 U109 ( .IN1(n82), .IN2(in2[21]), .Q(n88) );
  NOR2X0 U110 ( .IN1(n81), .IN2(n88), .QN(n87) );
  NOR2X0 U111 ( .IN1(in2[22]), .IN2(n81), .QN(n84) );
  NAND2X0 U112 ( .IN1(in2[21]), .IN2(n82), .QN(n83) );
  OA221X1 U113 ( .IN1(n84), .IN2(n89), .IN3(n84), .IN4(n83), .IN5(n88), .Q(n85) );
  AO221X1 U114 ( .IN1(in2[22]), .IN2(n87), .IN3(in2[22]), .IN4(n90), .IN5(n85), 
        .Q(out1[22]) );
  NOR2X0 U115 ( .IN1(n86), .IN2(n88), .QN(n93) );
  AO21X1 U116 ( .IN1(n89), .IN2(n88), .IN3(n87), .Q(n91) );
  AO221X1 U117 ( .IN1(in2[22]), .IN2(n93), .IN3(n20), .IN4(n91), .IN5(n90), 
        .Q(out1[23]) );
  AO21X1 U118 ( .IN1(n93), .IN2(n20), .IN3(n92), .Q(out1[24]) );
endmodule


module mul26_3 ( clk, rst_n, in1, in2, en, mulout );
  input [25:0] in1;
  input [25:0] in2;
  output [50:0] mulout;
  input clk, rst_n, en;
  wire   N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24,
         N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38,
         N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N62, N63,
         N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77,
         N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91,
         N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, n18, n19, n20,
         n21, n22, n23, n24, n25, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n124, n125, SYNOPSYS_UNCONNECTED_1,
         SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3,
         SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5,
         SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7,
         SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9,
         SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11,
         SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13,
         SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15,
         SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17,
         SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19,
         SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21,
         SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_23,
         SYNOPSYS_UNCONNECTED_24, SYNOPSYS_UNCONNECTED_25,
         SYNOPSYS_UNCONNECTED_26, SYNOPSYS_UNCONNECTED_27,
         SYNOPSYS_UNCONNECTED_28, SYNOPSYS_UNCONNECTED_29,
         SYNOPSYS_UNCONNECTED_30, SYNOPSYS_UNCONNECTED_31,
         SYNOPSYS_UNCONNECTED_32, SYNOPSYS_UNCONNECTED_33,
         SYNOPSYS_UNCONNECTED_34, SYNOPSYS_UNCONNECTED_35,
         SYNOPSYS_UNCONNECTED_36, SYNOPSYS_UNCONNECTED_37,
         SYNOPSYS_UNCONNECTED_38, SYNOPSYS_UNCONNECTED_39,
         SYNOPSYS_UNCONNECTED_40, SYNOPSYS_UNCONNECTED_41,
         SYNOPSYS_UNCONNECTED_42, SYNOPSYS_UNCONNECTED_43,
         SYNOPSYS_UNCONNECTED_44, SYNOPSYS_UNCONNECTED_45,
         SYNOPSYS_UNCONNECTED_46, SYNOPSYS_UNCONNECTED_47,
         SYNOPSYS_UNCONNECTED_48, SYNOPSYS_UNCONNECTED_49,
         SYNOPSYS_UNCONNECTED_50, SYNOPSYS_UNCONNECTED_51,
         SYNOPSYS_UNCONNECTED_52, SYNOPSYS_UNCONNECTED_53,
         SYNOPSYS_UNCONNECTED_54, SYNOPSYS_UNCONNECTED_55,
         SYNOPSYS_UNCONNECTED_56, SYNOPSYS_UNCONNECTED_57,
         SYNOPSYS_UNCONNECTED_58, SYNOPSYS_UNCONNECTED_59,
         SYNOPSYS_UNCONNECTED_60, SYNOPSYS_UNCONNECTED_61,
         SYNOPSYS_UNCONNECTED_62, SYNOPSYS_UNCONNECTED_63,
         SYNOPSYS_UNCONNECTED_64, SYNOPSYS_UNCONNECTED_65,
         SYNOPSYS_UNCONNECTED_66, SYNOPSYS_UNCONNECTED_67,
         SYNOPSYS_UNCONNECTED_68, SYNOPSYS_UNCONNECTED_69,
         SYNOPSYS_UNCONNECTED_70, SYNOPSYS_UNCONNECTED_71,
         SYNOPSYS_UNCONNECTED_72, SYNOPSYS_UNCONNECTED_73,
         SYNOPSYS_UNCONNECTED_74, SYNOPSYS_UNCONNECTED_75,
         SYNOPSYS_UNCONNECTED_76, SYNOPSYS_UNCONNECTED_77,
         SYNOPSYS_UNCONNECTED_78, SYNOPSYS_UNCONNECTED_79,
         SYNOPSYS_UNCONNECTED_80, SYNOPSYS_UNCONNECTED_81,
         SYNOPSYS_UNCONNECTED_82, SYNOPSYS_UNCONNECTED_83,
         SYNOPSYS_UNCONNECTED_84, SYNOPSYS_UNCONNECTED_85,
         SYNOPSYS_UNCONNECTED_86, SYNOPSYS_UNCONNECTED_87,
         SYNOPSYS_UNCONNECTED_88, SYNOPSYS_UNCONNECTED_89,
         SYNOPSYS_UNCONNECTED_90, SYNOPSYS_UNCONNECTED_91,
         SYNOPSYS_UNCONNECTED_92, SYNOPSYS_UNCONNECTED_93,
         SYNOPSYS_UNCONNECTED_94, SYNOPSYS_UNCONNECTED_95,
         SYNOPSYS_UNCONNECTED_96, SYNOPSYS_UNCONNECTED_97,
         SYNOPSYS_UNCONNECTED_98, SYNOPSYS_UNCONNECTED_99,
         SYNOPSYS_UNCONNECTED_100, SYNOPSYS_UNCONNECTED_101,
         SYNOPSYS_UNCONNECTED_102, SYNOPSYS_UNCONNECTED_103,
         SYNOPSYS_UNCONNECTED_104, SYNOPSYS_UNCONNECTED_105,
         SYNOPSYS_UNCONNECTED_106, SYNOPSYS_UNCONNECTED_107,
         SYNOPSYS_UNCONNECTED_108, SYNOPSYS_UNCONNECTED_109,
         SYNOPSYS_UNCONNECTED_110, SYNOPSYS_UNCONNECTED_111,
         SYNOPSYS_UNCONNECTED_112, SYNOPSYS_UNCONNECTED_113,
         SYNOPSYS_UNCONNECTED_114, SYNOPSYS_UNCONNECTED_115,
         SYNOPSYS_UNCONNECTED_116, SYNOPSYS_UNCONNECTED_117,
         SYNOPSYS_UNCONNECTED_118, SYNOPSYS_UNCONNECTED_119,
         SYNOPSYS_UNCONNECTED_120, SYNOPSYS_UNCONNECTED_121,
         SYNOPSYS_UNCONNECTED_122, SYNOPSYS_UNCONNECTED_123,
         SYNOPSYS_UNCONNECTED_124, SYNOPSYS_UNCONNECTED_125,
         SYNOPSYS_UNCONNECTED_126, SYNOPSYS_UNCONNECTED_127,
         SYNOPSYS_UNCONNECTED_128, SYNOPSYS_UNCONNECTED_129,
         SYNOPSYS_UNCONNECTED_130, SYNOPSYS_UNCONNECTED_131,
         SYNOPSYS_UNCONNECTED_132, SYNOPSYS_UNCONNECTED_133,
         SYNOPSYS_UNCONNECTED_134, SYNOPSYS_UNCONNECTED_135,
         SYNOPSYS_UNCONNECTED_136, SYNOPSYS_UNCONNECTED_137,
         SYNOPSYS_UNCONNECTED_138, SYNOPSYS_UNCONNECTED_139,
         SYNOPSYS_UNCONNECTED_140, SYNOPSYS_UNCONNECTED_141,
         SYNOPSYS_UNCONNECTED_142, SYNOPSYS_UNCONNECTED_143,
         SYNOPSYS_UNCONNECTED_144, SYNOPSYS_UNCONNECTED_145,
         SYNOPSYS_UNCONNECTED_146, SYNOPSYS_UNCONNECTED_147,
         SYNOPSYS_UNCONNECTED_148, SYNOPSYS_UNCONNECTED_149,
         SYNOPSYS_UNCONNECTED_150, SYNOPSYS_UNCONNECTED_151,
         SYNOPSYS_UNCONNECTED_152, SYNOPSYS_UNCONNECTED_153,
         SYNOPSYS_UNCONNECTED_154, SYNOPSYS_UNCONNECTED_155,
         SYNOPSYS_UNCONNECTED_156, SYNOPSYS_UNCONNECTED_157,
         SYNOPSYS_UNCONNECTED_158, SYNOPSYS_UNCONNECTED_159,
         SYNOPSYS_UNCONNECTED_160, SYNOPSYS_UNCONNECTED_161,
         SYNOPSYS_UNCONNECTED_162, SYNOPSYS_UNCONNECTED_163,
         SYNOPSYS_UNCONNECTED_164, SYNOPSYS_UNCONNECTED_165,
         SYNOPSYS_UNCONNECTED_166, SYNOPSYS_UNCONNECTED_167,
         SYNOPSYS_UNCONNECTED_168, SYNOPSYS_UNCONNECTED_169,
         SYNOPSYS_UNCONNECTED_170, SYNOPSYS_UNCONNECTED_171,
         SYNOPSYS_UNCONNECTED_172, SYNOPSYS_UNCONNECTED_173,
         SYNOPSYS_UNCONNECTED_174, SYNOPSYS_UNCONNECTED_175,
         SYNOPSYS_UNCONNECTED_176, SYNOPSYS_UNCONNECTED_177,
         SYNOPSYS_UNCONNECTED_178, SYNOPSYS_UNCONNECTED_179,
         SYNOPSYS_UNCONNECTED_180, SYNOPSYS_UNCONNECTED_181,
         SYNOPSYS_UNCONNECTED_182, SYNOPSYS_UNCONNECTED_183,
         SYNOPSYS_UNCONNECTED_184, SYNOPSYS_UNCONNECTED_185,
         SYNOPSYS_UNCONNECTED_186, SYNOPSYS_UNCONNECTED_187,
         SYNOPSYS_UNCONNECTED_188, SYNOPSYS_UNCONNECTED_189,
         SYNOPSYS_UNCONNECTED_190, SYNOPSYS_UNCONNECTED_191,
         SYNOPSYS_UNCONNECTED_192, SYNOPSYS_UNCONNECTED_193,
         SYNOPSYS_UNCONNECTED_194, SYNOPSYS_UNCONNECTED_195,
         SYNOPSYS_UNCONNECTED_196, SYNOPSYS_UNCONNECTED_197,
         SYNOPSYS_UNCONNECTED_198, SYNOPSYS_UNCONNECTED_199,
         SYNOPSYS_UNCONNECTED_200, SYNOPSYS_UNCONNECTED_201,
         SYNOPSYS_UNCONNECTED_202, SYNOPSYS_UNCONNECTED_203,
         SYNOPSYS_UNCONNECTED_204, SYNOPSYS_UNCONNECTED_205,
         SYNOPSYS_UNCONNECTED_206, SYNOPSYS_UNCONNECTED_207,
         SYNOPSYS_UNCONNECTED_208, SYNOPSYS_UNCONNECTED_209,
         SYNOPSYS_UNCONNECTED_210, SYNOPSYS_UNCONNECTED_211,
         SYNOPSYS_UNCONNECTED_212, SYNOPSYS_UNCONNECTED_213,
         SYNOPSYS_UNCONNECTED_214, SYNOPSYS_UNCONNECTED_215,
         SYNOPSYS_UNCONNECTED_216, SYNOPSYS_UNCONNECTED_217,
         SYNOPSYS_UNCONNECTED_218, SYNOPSYS_UNCONNECTED_219,
         SYNOPSYS_UNCONNECTED_220, SYNOPSYS_UNCONNECTED_221,
         SYNOPSYS_UNCONNECTED_222, SYNOPSYS_UNCONNECTED_223,
         SYNOPSYS_UNCONNECTED_224, SYNOPSYS_UNCONNECTED_225,
         SYNOPSYS_UNCONNECTED_226, SYNOPSYS_UNCONNECTED_227,
         SYNOPSYS_UNCONNECTED_228, SYNOPSYS_UNCONNECTED_229,
         SYNOPSYS_UNCONNECTED_230, SYNOPSYS_UNCONNECTED_231,
         SYNOPSYS_UNCONNECTED_232, SYNOPSYS_UNCONNECTED_233,
         SYNOPSYS_UNCONNECTED_234, SYNOPSYS_UNCONNECTED_235,
         SYNOPSYS_UNCONNECTED_236, SYNOPSYS_UNCONNECTED_237,
         SYNOPSYS_UNCONNECTED_238, SYNOPSYS_UNCONNECTED_239,
         SYNOPSYS_UNCONNECTED_240, SYNOPSYS_UNCONNECTED_241,
         SYNOPSYS_UNCONNECTED_242, SYNOPSYS_UNCONNECTED_243,
         SYNOPSYS_UNCONNECTED_244, SYNOPSYS_UNCONNECTED_245,
         SYNOPSYS_UNCONNECTED_246, SYNOPSYS_UNCONNECTED_247,
         SYNOPSYS_UNCONNECTED_248, SYNOPSYS_UNCONNECTED_249,
         SYNOPSYS_UNCONNECTED_250, SYNOPSYS_UNCONNECTED_251,
         SYNOPSYS_UNCONNECTED_252, SYNOPSYS_UNCONNECTED_253,
         SYNOPSYS_UNCONNECTED_254, SYNOPSYS_UNCONNECTED_255,
         SYNOPSYS_UNCONNECTED_256, SYNOPSYS_UNCONNECTED_257,
         SYNOPSYS_UNCONNECTED_258, SYNOPSYS_UNCONNECTED_259,
         SYNOPSYS_UNCONNECTED_260, SYNOPSYS_UNCONNECTED_261,
         SYNOPSYS_UNCONNECTED_262, SYNOPSYS_UNCONNECTED_263,
         SYNOPSYS_UNCONNECTED_264, SYNOPSYS_UNCONNECTED_265,
         SYNOPSYS_UNCONNECTED_266, SYNOPSYS_UNCONNECTED_267,
         SYNOPSYS_UNCONNECTED_268, SYNOPSYS_UNCONNECTED_269,
         SYNOPSYS_UNCONNECTED_270, SYNOPSYS_UNCONNECTED_271,
         SYNOPSYS_UNCONNECTED_272, SYNOPSYS_UNCONNECTED_273,
         SYNOPSYS_UNCONNECTED_274, SYNOPSYS_UNCONNECTED_275,
         SYNOPSYS_UNCONNECTED_276, SYNOPSYS_UNCONNECTED_277,
         SYNOPSYS_UNCONNECTED_278, SYNOPSYS_UNCONNECTED_279,
         SYNOPSYS_UNCONNECTED_280, SYNOPSYS_UNCONNECTED_281,
         SYNOPSYS_UNCONNECTED_282, SYNOPSYS_UNCONNECTED_283,
         SYNOPSYS_UNCONNECTED_284, SYNOPSYS_UNCONNECTED_285,
         SYNOPSYS_UNCONNECTED_286, SYNOPSYS_UNCONNECTED_287,
         SYNOPSYS_UNCONNECTED_288, SYNOPSYS_UNCONNECTED_289,
         SYNOPSYS_UNCONNECTED_290, SYNOPSYS_UNCONNECTED_291,
         SYNOPSYS_UNCONNECTED_292, SYNOPSYS_UNCONNECTED_293,
         SYNOPSYS_UNCONNECTED_294, SYNOPSYS_UNCONNECTED_295,
         SYNOPSYS_UNCONNECTED_296, SYNOPSYS_UNCONNECTED_297,
         SYNOPSYS_UNCONNECTED_298, SYNOPSYS_UNCONNECTED_299,
         SYNOPSYS_UNCONNECTED_300, SYNOPSYS_UNCONNECTED_301,
         SYNOPSYS_UNCONNECTED_302, SYNOPSYS_UNCONNECTED_303,
         SYNOPSYS_UNCONNECTED_304, SYNOPSYS_UNCONNECTED_305,
         SYNOPSYS_UNCONNECTED_306, SYNOPSYS_UNCONNECTED_307,
         SYNOPSYS_UNCONNECTED_308, SYNOPSYS_UNCONNECTED_309,
         SYNOPSYS_UNCONNECTED_310, SYNOPSYS_UNCONNECTED_311,
         SYNOPSYS_UNCONNECTED_312, SYNOPSYS_UNCONNECTED_313,
         SYNOPSYS_UNCONNECTED_314, SYNOPSYS_UNCONNECTED_315,
         SYNOPSYS_UNCONNECTED_316, SYNOPSYS_UNCONNECTED_317,
         SYNOPSYS_UNCONNECTED_318, SYNOPSYS_UNCONNECTED_319,
         SYNOPSYS_UNCONNECTED_320, SYNOPSYS_UNCONNECTED_321,
         SYNOPSYS_UNCONNECTED_322, SYNOPSYS_UNCONNECTED_323,
         SYNOPSYS_UNCONNECTED_324, SYNOPSYS_UNCONNECTED_325,
         SYNOPSYS_UNCONNECTED_326, SYNOPSYS_UNCONNECTED_327,
         SYNOPSYS_UNCONNECTED_328, SYNOPSYS_UNCONNECTED_329,
         SYNOPSYS_UNCONNECTED_330, SYNOPSYS_UNCONNECTED_331,
         SYNOPSYS_UNCONNECTED_332, SYNOPSYS_UNCONNECTED_333,
         SYNOPSYS_UNCONNECTED_334, SYNOPSYS_UNCONNECTED_335,
         SYNOPSYS_UNCONNECTED_336, SYNOPSYS_UNCONNECTED_337,
         SYNOPSYS_UNCONNECTED_338, SYNOPSYS_UNCONNECTED_339,
         SYNOPSYS_UNCONNECTED_340, SYNOPSYS_UNCONNECTED_341,
         SYNOPSYS_UNCONNECTED_342, SYNOPSYS_UNCONNECTED_343,
         SYNOPSYS_UNCONNECTED_344, SYNOPSYS_UNCONNECTED_345,
         SYNOPSYS_UNCONNECTED_346, SYNOPSYS_UNCONNECTED_347,
         SYNOPSYS_UNCONNECTED_348, SYNOPSYS_UNCONNECTED_349,
         SYNOPSYS_UNCONNECTED_350, SYNOPSYS_UNCONNECTED_351,
         SYNOPSYS_UNCONNECTED_352, SYNOPSYS_UNCONNECTED_353,
         SYNOPSYS_UNCONNECTED_354, SYNOPSYS_UNCONNECTED_355,
         SYNOPSYS_UNCONNECTED_356, SYNOPSYS_UNCONNECTED_357,
         SYNOPSYS_UNCONNECTED_358, SYNOPSYS_UNCONNECTED_359,
         SYNOPSYS_UNCONNECTED_360, SYNOPSYS_UNCONNECTED_361,
         SYNOPSYS_UNCONNECTED_362, SYNOPSYS_UNCONNECTED_363,
         SYNOPSYS_UNCONNECTED_364, SYNOPSYS_UNCONNECTED_365,
         SYNOPSYS_UNCONNECTED_366, SYNOPSYS_UNCONNECTED_367,
         SYNOPSYS_UNCONNECTED_368, SYNOPSYS_UNCONNECTED_369,
         SYNOPSYS_UNCONNECTED_370, SYNOPSYS_UNCONNECTED_371,
         SYNOPSYS_UNCONNECTED_372, SYNOPSYS_UNCONNECTED_373,
         SYNOPSYS_UNCONNECTED_374, SYNOPSYS_UNCONNECTED_375,
         SYNOPSYS_UNCONNECTED_376, SYNOPSYS_UNCONNECTED_377,
         SYNOPSYS_UNCONNECTED_378, SYNOPSYS_UNCONNECTED_379,
         SYNOPSYS_UNCONNECTED_380, SYNOPSYS_UNCONNECTED_381,
         SYNOPSYS_UNCONNECTED_382, SYNOPSYS_UNCONNECTED_383,
         SYNOPSYS_UNCONNECTED_384, SYNOPSYS_UNCONNECTED_385,
         SYNOPSYS_UNCONNECTED_386, SYNOPSYS_UNCONNECTED_387,
         SYNOPSYS_UNCONNECTED_388, SYNOPSYS_UNCONNECTED_389,
         SYNOPSYS_UNCONNECTED_390, SYNOPSYS_UNCONNECTED_391,
         SYNOPSYS_UNCONNECTED_392, SYNOPSYS_UNCONNECTED_393,
         SYNOPSYS_UNCONNECTED_394, SYNOPSYS_UNCONNECTED_395,
         SYNOPSYS_UNCONNECTED_396, SYNOPSYS_UNCONNECTED_397,
         SYNOPSYS_UNCONNECTED_398, SYNOPSYS_UNCONNECTED_399,
         SYNOPSYS_UNCONNECTED_400, SYNOPSYS_UNCONNECTED_401,
         SYNOPSYS_UNCONNECTED_402, SYNOPSYS_UNCONNECTED_403,
         SYNOPSYS_UNCONNECTED_404, SYNOPSYS_UNCONNECTED_405,
         SYNOPSYS_UNCONNECTED_406, SYNOPSYS_UNCONNECTED_407,
         SYNOPSYS_UNCONNECTED_408, SYNOPSYS_UNCONNECTED_409,
         SYNOPSYS_UNCONNECTED_410, SYNOPSYS_UNCONNECTED_411,
         SYNOPSYS_UNCONNECTED_412, SYNOPSYS_UNCONNECTED_413,
         SYNOPSYS_UNCONNECTED_414;
  wire   [26:2] boothout1;
  wire   [26:0] boothout2;
  wire   [26:0] boothout3;
  wire   [26:0] boothout4;
  wire   [26:0] boothout5;
  wire   [26:0] boothout6;
  wire   [24:0] boothout7;
  wire   [26:0] boothout8;
  wire   [26:0] boothout9;
  wire   [26:0] boothout10;
  wire   [26:0] boothout11;
  wire   [25:0] boothout12;
  wire   [22:0] boothout13;
  wire   [29:2] cout1;
  wire   [31:3] mulout1;
  wire   [35:8] cout2;
  wire   [37:6] mulout2;
  wire   [41:14] cout3;
  wire   [42:12] mulout3;
  wire   [46:20] cout4;
  wire   [47:18] mulout4;
  wire   [31:3] cout5;
  wire   [46:4] mulout5;
  wire   [37:9] cout6;
  wire   [42:6] mulout6;
  wire   [46:18] cout7;
  wire   [47:12] mulout7;
  wire   [38:4] cout8;
  wire   [46:5] mulout8;
  wire   [46:12] cout9;
  wire   [47:6] mulout9;
  wire   [46:5] cout10;
  wire   [47:6] mulout10;
  wire   [46:6] cout11;
  wire   [47:7] mulout11;
  wire   [47:0] a;
  wire   [47:8] b;

  booth27_39 booth1 ( .out1({boothout1, SYNOPSYS_UNCONNECTED_1, 
        SYNOPSYS_UNCONNECTED_2}), .in1({in1[1:0], 1'b0}), .in2({1'b0, 1'b0, 
        1'b1, in2[22:19], n25, in2[17:16], n24, in2[14:13], n23, n22, in2[10], 
        n21, in2[8:4], n20, in2[2], n19, n18}) );
  booth27_38 booth2 ( .out1(boothout2), .in1(in1[3:1]), .in2({1'b0, 1'b0, 1'b1, 
        in2[22:19], n25, in2[17:16], n24, in2[14:13], n23, n22, in2[10], n21, 
        in2[8:4], n20, in2[2], n19, n18}) );
  booth27_37 booth3 ( .out1(boothout3), .in1(in1[5:3]), .in2({1'b0, 1'b0, 1'b1, 
        in2[22:19], n25, in2[17:16], n24, in2[14:13], n23, n22, in2[10], n21, 
        in2[8:4], n20, in2[2], n19, n18}) );
  booth27_36 booth4 ( .out1(boothout4), .in1({in1[7], 1'b0, in1[5]}), .in2({
        1'b0, 1'b0, 1'b1, in2[22:19], n25, in2[17:16], n24, in2[14:13], n23, 
        n22, in2[10], n21, in2[8:4], n20, in2[2], n19, n18}) );
  booth27_35 booth5 ( .out1(boothout5), .in1(in1[9:7]), .in2({1'b0, 1'b0, 1'b1, 
        in2[22:19], n25, in2[17:16], n24, in2[14:13], n23, n22, in2[10], n21, 
        in2[8:4], n20, in2[2], n19, n18}) );
  booth27_34 booth6 ( .out1(boothout6), .in1(in1[11:9]), .in2({1'b0, 1'b0, 
        1'b1, in2[22:19], n25, in2[17:16], n24, in2[14:13], n23, n22, in2[10], 
        n21, in2[8:4], n20, in2[2], n19, n18}) );
  booth27_33 booth7 ( .out1({SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4, 
        boothout7}), .in1({1'b0, in1[12:11]}), .in2({1'b0, 1'b0, 1'b1, 
        in2[22:19], n25, in2[17:16], n24, in2[14:13], n23, n22, in2[10], n21, 
        in2[8:4], n20, in2[2], n19, n18}) );
  booth27_32 booth8 ( .out1(boothout8), .in1({in1[15:14], 1'b0}), .in2({1'b0, 
        1'b0, 1'b1, in2[22:19], n25, in2[17:16], n24, in2[14:13], n23, n22, 
        in2[10], n21, in2[8:4], n20, in2[2], n19, n18}) );
  booth27_31 booth9 ( .out1(boothout9), .in1(in1[17:15]), .in2({1'b0, 1'b0, 
        1'b1, in2[22:19], n25, in2[17:16], n24, in2[14:13], n23, n22, in2[10], 
        n21, in2[8:4], n20, in2[2], n19, n18}) );
  booth27_30 booth10 ( .out1(boothout10), .in1(in1[19:17]), .in2({1'b0, 1'b0, 
        1'b1, in2[22:19], n25, in2[17:16], n24, in2[14:13], n23, n22, in2[10], 
        n21, in2[8:4], n20, in2[2], n19, n18}) );
  booth27_29 booth11 ( .out1(boothout11), .in1(in1[21:19]), .in2({1'b0, 1'b0, 
        1'b1, in2[22:19], n25, in2[17:16], n24, in2[14:13], n23, n22, in2[10], 
        n21, in2[8:4], n20, in2[2], n19, n18}) );
  booth27_28 booth12 ( .out1({SYNOPSYS_UNCONNECTED_5, boothout12}), .in1({1'b1, 
        in1[22:21]}), .in2({1'b0, 1'b0, 1'b1, in2[22:19], n25, in2[17:16], n24, 
        in2[14:13], n23, n22, in2[10], n21, in2[8:4], n20, in2[2], n19, n18})
         );
  booth27_27 booth13 ( .out1({SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, 
        SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, boothout13}), .in1({
        1'b0, 1'b0, 1'b1}), .in2({1'b0, 1'b0, 1'b1, in2[22:19], n25, 
        in2[17:16], n24, in2[14:13], n23, n22, in2[10], n21, in2[8:4], n20, 
        in2[2], n19, n18}) );
  csa51squ_36 csa51squ1 ( .cout({SYNOPSYS_UNCONNECTED_10, 
        SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12, 
        SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14, 
        SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16, 
        SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18, 
        SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20, 
        SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22, 
        SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24, 
        SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26, 
        SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28, 
        SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30, cout1, 
        SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32}), .sumout({
        SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34, 
        SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36, 
        SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38, 
        SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40, 
        SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42, 
        SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44, 
        SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46, 
        SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48, 
        SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50, 
        SYNOPSYS_UNCONNECTED_51, mulout1[31], SYNOPSYS_UNCONNECTED_52, 
        mulout1[29:3], SYNOPSYS_UNCONNECTED_53, SYNOPSYS_UNCONNECTED_54, 
        SYNOPSYS_UNCONNECTED_55}), .in1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, boothout1, 1'b0, 1'b0}), .in2({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, boothout2, 
        1'b0, 1'b0}), .in3({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n125, 
        1'b0, boothout3[25:0], 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_35 csa51squ2 ( .cout({SYNOPSYS_UNCONNECTED_56, 
        SYNOPSYS_UNCONNECTED_57, SYNOPSYS_UNCONNECTED_58, 
        SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_60, 
        SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_62, 
        SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_64, 
        SYNOPSYS_UNCONNECTED_65, SYNOPSYS_UNCONNECTED_66, 
        SYNOPSYS_UNCONNECTED_67, SYNOPSYS_UNCONNECTED_68, 
        SYNOPSYS_UNCONNECTED_69, SYNOPSYS_UNCONNECTED_70, cout2, 
        SYNOPSYS_UNCONNECTED_71, SYNOPSYS_UNCONNECTED_72, 
        SYNOPSYS_UNCONNECTED_73, SYNOPSYS_UNCONNECTED_74, 
        SYNOPSYS_UNCONNECTED_75, SYNOPSYS_UNCONNECTED_76, 
        SYNOPSYS_UNCONNECTED_77, SYNOPSYS_UNCONNECTED_78}), .sumout({
        SYNOPSYS_UNCONNECTED_79, SYNOPSYS_UNCONNECTED_80, 
        SYNOPSYS_UNCONNECTED_81, SYNOPSYS_UNCONNECTED_82, 
        SYNOPSYS_UNCONNECTED_83, SYNOPSYS_UNCONNECTED_84, 
        SYNOPSYS_UNCONNECTED_85, SYNOPSYS_UNCONNECTED_86, 
        SYNOPSYS_UNCONNECTED_87, SYNOPSYS_UNCONNECTED_88, 
        SYNOPSYS_UNCONNECTED_89, SYNOPSYS_UNCONNECTED_90, 
        SYNOPSYS_UNCONNECTED_91, mulout2[37], SYNOPSYS_UNCONNECTED_92, 
        mulout2[35:6], SYNOPSYS_UNCONNECTED_93, SYNOPSYS_UNCONNECTED_94, 
        SYNOPSYS_UNCONNECTED_95, SYNOPSYS_UNCONNECTED_96, 
        SYNOPSYS_UNCONNECTED_97, SYNOPSYS_UNCONNECTED_98}), .in1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, boothout4, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, boothout5, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .in3({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n124, 1'b0, boothout6[25:0], 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_34 csa51squ3 ( .cout({SYNOPSYS_UNCONNECTED_99, 
        SYNOPSYS_UNCONNECTED_100, SYNOPSYS_UNCONNECTED_101, 
        SYNOPSYS_UNCONNECTED_102, SYNOPSYS_UNCONNECTED_103, 
        SYNOPSYS_UNCONNECTED_104, SYNOPSYS_UNCONNECTED_105, 
        SYNOPSYS_UNCONNECTED_106, SYNOPSYS_UNCONNECTED_107, cout3, 
        SYNOPSYS_UNCONNECTED_108, SYNOPSYS_UNCONNECTED_109, 
        SYNOPSYS_UNCONNECTED_110, SYNOPSYS_UNCONNECTED_111, 
        SYNOPSYS_UNCONNECTED_112, SYNOPSYS_UNCONNECTED_113, 
        SYNOPSYS_UNCONNECTED_114, SYNOPSYS_UNCONNECTED_115, 
        SYNOPSYS_UNCONNECTED_116, SYNOPSYS_UNCONNECTED_117, 
        SYNOPSYS_UNCONNECTED_118, SYNOPSYS_UNCONNECTED_119, 
        SYNOPSYS_UNCONNECTED_120, SYNOPSYS_UNCONNECTED_121}), .sumout({
        SYNOPSYS_UNCONNECTED_122, SYNOPSYS_UNCONNECTED_123, 
        SYNOPSYS_UNCONNECTED_124, SYNOPSYS_UNCONNECTED_125, 
        SYNOPSYS_UNCONNECTED_126, SYNOPSYS_UNCONNECTED_127, 
        SYNOPSYS_UNCONNECTED_128, SYNOPSYS_UNCONNECTED_129, mulout3, 
        SYNOPSYS_UNCONNECTED_130, SYNOPSYS_UNCONNECTED_131, 
        SYNOPSYS_UNCONNECTED_132, SYNOPSYS_UNCONNECTED_133, 
        SYNOPSYS_UNCONNECTED_134, SYNOPSYS_UNCONNECTED_135, 
        SYNOPSYS_UNCONNECTED_136, SYNOPSYS_UNCONNECTED_137, 
        SYNOPSYS_UNCONNECTED_138, SYNOPSYS_UNCONNECTED_139, 
        SYNOPSYS_UNCONNECTED_140, SYNOPSYS_UNCONNECTED_141}), .in1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 
        boothout7, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .in2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, boothout8, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in3({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, boothout9, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_33 csa51squ4 ( .cout({SYNOPSYS_UNCONNECTED_142, 
        SYNOPSYS_UNCONNECTED_143, SYNOPSYS_UNCONNECTED_144, 
        SYNOPSYS_UNCONNECTED_145, cout4, SYNOPSYS_UNCONNECTED_146, 
        SYNOPSYS_UNCONNECTED_147, SYNOPSYS_UNCONNECTED_148, 
        SYNOPSYS_UNCONNECTED_149, SYNOPSYS_UNCONNECTED_150, 
        SYNOPSYS_UNCONNECTED_151, SYNOPSYS_UNCONNECTED_152, 
        SYNOPSYS_UNCONNECTED_153, SYNOPSYS_UNCONNECTED_154, 
        SYNOPSYS_UNCONNECTED_155, SYNOPSYS_UNCONNECTED_156, 
        SYNOPSYS_UNCONNECTED_157, SYNOPSYS_UNCONNECTED_158, 
        SYNOPSYS_UNCONNECTED_159, SYNOPSYS_UNCONNECTED_160, 
        SYNOPSYS_UNCONNECTED_161, SYNOPSYS_UNCONNECTED_162, 
        SYNOPSYS_UNCONNECTED_163, SYNOPSYS_UNCONNECTED_164, 
        SYNOPSYS_UNCONNECTED_165}), .sumout({SYNOPSYS_UNCONNECTED_166, 
        SYNOPSYS_UNCONNECTED_167, SYNOPSYS_UNCONNECTED_168, mulout4, 
        SYNOPSYS_UNCONNECTED_169, SYNOPSYS_UNCONNECTED_170, 
        SYNOPSYS_UNCONNECTED_171, SYNOPSYS_UNCONNECTED_172, 
        SYNOPSYS_UNCONNECTED_173, SYNOPSYS_UNCONNECTED_174, 
        SYNOPSYS_UNCONNECTED_175, SYNOPSYS_UNCONNECTED_176, 
        SYNOPSYS_UNCONNECTED_177, SYNOPSYS_UNCONNECTED_178, 
        SYNOPSYS_UNCONNECTED_179, SYNOPSYS_UNCONNECTED_180, 
        SYNOPSYS_UNCONNECTED_181, SYNOPSYS_UNCONNECTED_182, 
        SYNOPSYS_UNCONNECTED_183, SYNOPSYS_UNCONNECTED_184, 
        SYNOPSYS_UNCONNECTED_185, SYNOPSYS_UNCONNECTED_186}), .in1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, boothout10, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 1'b0, 1'b0, 1'b0, boothout11, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .in3({1'b0, 1'b0, 1'b0, boothout12, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_32 csa51squ5 ( .cout({SYNOPSYS_UNCONNECTED_187, 
        SYNOPSYS_UNCONNECTED_188, SYNOPSYS_UNCONNECTED_189, 
        SYNOPSYS_UNCONNECTED_190, SYNOPSYS_UNCONNECTED_191, 
        SYNOPSYS_UNCONNECTED_192, SYNOPSYS_UNCONNECTED_193, 
        SYNOPSYS_UNCONNECTED_194, SYNOPSYS_UNCONNECTED_195, 
        SYNOPSYS_UNCONNECTED_196, SYNOPSYS_UNCONNECTED_197, 
        SYNOPSYS_UNCONNECTED_198, SYNOPSYS_UNCONNECTED_199, 
        SYNOPSYS_UNCONNECTED_200, SYNOPSYS_UNCONNECTED_201, 
        SYNOPSYS_UNCONNECTED_202, SYNOPSYS_UNCONNECTED_203, 
        SYNOPSYS_UNCONNECTED_204, SYNOPSYS_UNCONNECTED_205, cout5, 
        SYNOPSYS_UNCONNECTED_206, SYNOPSYS_UNCONNECTED_207, 
        SYNOPSYS_UNCONNECTED_208}), .sumout({SYNOPSYS_UNCONNECTED_209, 
        SYNOPSYS_UNCONNECTED_210, SYNOPSYS_UNCONNECTED_211, 
        SYNOPSYS_UNCONNECTED_212, mulout5, SYNOPSYS_UNCONNECTED_213, 
        SYNOPSYS_UNCONNECTED_214, SYNOPSYS_UNCONNECTED_215, 
        SYNOPSYS_UNCONNECTED_216}), .in1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, cout1, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, mulout1[31], 1'b0, mulout1[29:3], 1'b0, 1'b0, 1'b0}), 
        .in3({1'b0, 1'b0, 1'b0, 1'b1, boothout13, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_31 csa51squ6 ( .cout({SYNOPSYS_UNCONNECTED_217, 
        SYNOPSYS_UNCONNECTED_218, SYNOPSYS_UNCONNECTED_219, 
        SYNOPSYS_UNCONNECTED_220, SYNOPSYS_UNCONNECTED_221, 
        SYNOPSYS_UNCONNECTED_222, SYNOPSYS_UNCONNECTED_223, 
        SYNOPSYS_UNCONNECTED_224, SYNOPSYS_UNCONNECTED_225, 
        SYNOPSYS_UNCONNECTED_226, SYNOPSYS_UNCONNECTED_227, 
        SYNOPSYS_UNCONNECTED_228, SYNOPSYS_UNCONNECTED_229, cout6, 
        SYNOPSYS_UNCONNECTED_230, SYNOPSYS_UNCONNECTED_231, 
        SYNOPSYS_UNCONNECTED_232, SYNOPSYS_UNCONNECTED_233, 
        SYNOPSYS_UNCONNECTED_234, SYNOPSYS_UNCONNECTED_235, 
        SYNOPSYS_UNCONNECTED_236, SYNOPSYS_UNCONNECTED_237, 
        SYNOPSYS_UNCONNECTED_238}), .sumout({SYNOPSYS_UNCONNECTED_239, 
        SYNOPSYS_UNCONNECTED_240, SYNOPSYS_UNCONNECTED_241, 
        SYNOPSYS_UNCONNECTED_242, SYNOPSYS_UNCONNECTED_243, 
        SYNOPSYS_UNCONNECTED_244, SYNOPSYS_UNCONNECTED_245, 
        SYNOPSYS_UNCONNECTED_246, mulout6, SYNOPSYS_UNCONNECTED_247, 
        SYNOPSYS_UNCONNECTED_248, SYNOPSYS_UNCONNECTED_249, 
        SYNOPSYS_UNCONNECTED_250, SYNOPSYS_UNCONNECTED_251, 
        SYNOPSYS_UNCONNECTED_252}), .in1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, cout2, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        mulout2[37], 1'b0, mulout2[35:6], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .in3({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, cout3, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  csa51squ_30 csa51squ7 ( .cout({SYNOPSYS_UNCONNECTED_253, 
        SYNOPSYS_UNCONNECTED_254, SYNOPSYS_UNCONNECTED_255, 
        SYNOPSYS_UNCONNECTED_256, cout7, SYNOPSYS_UNCONNECTED_257, 
        SYNOPSYS_UNCONNECTED_258, SYNOPSYS_UNCONNECTED_259, 
        SYNOPSYS_UNCONNECTED_260, SYNOPSYS_UNCONNECTED_261, 
        SYNOPSYS_UNCONNECTED_262, SYNOPSYS_UNCONNECTED_263, 
        SYNOPSYS_UNCONNECTED_264, SYNOPSYS_UNCONNECTED_265, 
        SYNOPSYS_UNCONNECTED_266, SYNOPSYS_UNCONNECTED_267, 
        SYNOPSYS_UNCONNECTED_268, SYNOPSYS_UNCONNECTED_269, 
        SYNOPSYS_UNCONNECTED_270, SYNOPSYS_UNCONNECTED_271, 
        SYNOPSYS_UNCONNECTED_272, SYNOPSYS_UNCONNECTED_273, 
        SYNOPSYS_UNCONNECTED_274}), .sumout({SYNOPSYS_UNCONNECTED_275, 
        SYNOPSYS_UNCONNECTED_276, SYNOPSYS_UNCONNECTED_277, mulout7, 
        SYNOPSYS_UNCONNECTED_278, SYNOPSYS_UNCONNECTED_279, 
        SYNOPSYS_UNCONNECTED_280, SYNOPSYS_UNCONNECTED_281, 
        SYNOPSYS_UNCONNECTED_282, SYNOPSYS_UNCONNECTED_283, 
        SYNOPSYS_UNCONNECTED_284, SYNOPSYS_UNCONNECTED_285, 
        SYNOPSYS_UNCONNECTED_286, SYNOPSYS_UNCONNECTED_287, 
        SYNOPSYS_UNCONNECTED_288, SYNOPSYS_UNCONNECTED_289}), .in1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mulout3, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 1'b0, 
        1'b0, cout4, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in3({1'b0, 1'b0, 1'b0, mulout4, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_29 csa51squ8 ( .cout({SYNOPSYS_UNCONNECTED_290, 
        SYNOPSYS_UNCONNECTED_291, SYNOPSYS_UNCONNECTED_292, 
        SYNOPSYS_UNCONNECTED_293, SYNOPSYS_UNCONNECTED_294, 
        SYNOPSYS_UNCONNECTED_295, SYNOPSYS_UNCONNECTED_296, 
        SYNOPSYS_UNCONNECTED_297, SYNOPSYS_UNCONNECTED_298, 
        SYNOPSYS_UNCONNECTED_299, SYNOPSYS_UNCONNECTED_300, 
        SYNOPSYS_UNCONNECTED_301, cout8, SYNOPSYS_UNCONNECTED_302, 
        SYNOPSYS_UNCONNECTED_303, SYNOPSYS_UNCONNECTED_304, 
        SYNOPSYS_UNCONNECTED_305}), .sumout({SYNOPSYS_UNCONNECTED_306, 
        SYNOPSYS_UNCONNECTED_307, SYNOPSYS_UNCONNECTED_308, 
        SYNOPSYS_UNCONNECTED_309, mulout8, SYNOPSYS_UNCONNECTED_310, 
        SYNOPSYS_UNCONNECTED_311, SYNOPSYS_UNCONNECTED_312, 
        SYNOPSYS_UNCONNECTED_313, SYNOPSYS_UNCONNECTED_314}), .in1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, cout5, 1'b0, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 
        1'b0, 1'b0, 1'b1, mulout5, 1'b0, 1'b0, 1'b0, 1'b0}), .in3({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, cout6, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_28 csa51squ9 ( .cout({SYNOPSYS_UNCONNECTED_315, 
        SYNOPSYS_UNCONNECTED_316, SYNOPSYS_UNCONNECTED_317, 
        SYNOPSYS_UNCONNECTED_318, cout9, SYNOPSYS_UNCONNECTED_319, 
        SYNOPSYS_UNCONNECTED_320, SYNOPSYS_UNCONNECTED_321, 
        SYNOPSYS_UNCONNECTED_322, SYNOPSYS_UNCONNECTED_323, 
        SYNOPSYS_UNCONNECTED_324, SYNOPSYS_UNCONNECTED_325, 
        SYNOPSYS_UNCONNECTED_326, SYNOPSYS_UNCONNECTED_327, 
        SYNOPSYS_UNCONNECTED_328, SYNOPSYS_UNCONNECTED_329, 
        SYNOPSYS_UNCONNECTED_330}), .sumout({SYNOPSYS_UNCONNECTED_331, 
        SYNOPSYS_UNCONNECTED_332, SYNOPSYS_UNCONNECTED_333, mulout9, 
        SYNOPSYS_UNCONNECTED_334, SYNOPSYS_UNCONNECTED_335, 
        SYNOPSYS_UNCONNECTED_336, SYNOPSYS_UNCONNECTED_337, 
        SYNOPSYS_UNCONNECTED_338, SYNOPSYS_UNCONNECTED_339}), .in1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mulout6, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .in2({1'b0, 1'b0, 1'b0, cout7, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .in3({1'b0, 1'b0, 1'b0, mulout7, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_27 csa51squ10 ( .cout({SYNOPSYS_UNCONNECTED_340, 
        SYNOPSYS_UNCONNECTED_341, SYNOPSYS_UNCONNECTED_342, 
        SYNOPSYS_UNCONNECTED_343, cout10, SYNOPSYS_UNCONNECTED_344, 
        SYNOPSYS_UNCONNECTED_345, SYNOPSYS_UNCONNECTED_346, 
        SYNOPSYS_UNCONNECTED_347, SYNOPSYS_UNCONNECTED_348}), .sumout({
        SYNOPSYS_UNCONNECTED_349, SYNOPSYS_UNCONNECTED_350, 
        SYNOPSYS_UNCONNECTED_351, mulout10, SYNOPSYS_UNCONNECTED_352, 
        SYNOPSYS_UNCONNECTED_353, SYNOPSYS_UNCONNECTED_354, 
        SYNOPSYS_UNCONNECTED_355, SYNOPSYS_UNCONNECTED_356, 
        SYNOPSYS_UNCONNECTED_357}), .in1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, cout8, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .in2({1'b0, 1'b0, 1'b0, 1'b1, mulout8, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .in3({1'b0, 1'b0, 1'b0, cout9, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_26 csa51squ11 ( .cout({SYNOPSYS_UNCONNECTED_358, 
        SYNOPSYS_UNCONNECTED_359, SYNOPSYS_UNCONNECTED_360, 
        SYNOPSYS_UNCONNECTED_361, cout11, SYNOPSYS_UNCONNECTED_362, 
        SYNOPSYS_UNCONNECTED_363, SYNOPSYS_UNCONNECTED_364, 
        SYNOPSYS_UNCONNECTED_365, SYNOPSYS_UNCONNECTED_366, 
        SYNOPSYS_UNCONNECTED_367}), .sumout({SYNOPSYS_UNCONNECTED_368, 
        SYNOPSYS_UNCONNECTED_369, SYNOPSYS_UNCONNECTED_370, mulout11, 
        SYNOPSYS_UNCONNECTED_371, SYNOPSYS_UNCONNECTED_372, 
        SYNOPSYS_UNCONNECTED_373, SYNOPSYS_UNCONNECTED_374, 
        SYNOPSYS_UNCONNECTED_375, SYNOPSYS_UNCONNECTED_376, 
        SYNOPSYS_UNCONNECTED_377}), .in1({1'b0, 1'b0, 1'b0, mulout9, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 1'b0, 1'b0, cout10, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in3({1'b0, 1'b0, 1'b0, mulout10, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  csa51squ_25 csa51squ12 ( .sumout({SYNOPSYS_UNCONNECTED_378, 
        SYNOPSYS_UNCONNECTED_379, SYNOPSYS_UNCONNECTED_380, N101, N100, N99, 
        N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, 
        N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, 
        N70, N69, N68, N67, N66, N65, N64, N63, N62, SYNOPSYS_UNCONNECTED_381, 
        SYNOPSYS_UNCONNECTED_382, SYNOPSYS_UNCONNECTED_383, 
        SYNOPSYS_UNCONNECTED_384, SYNOPSYS_UNCONNECTED_385, 
        SYNOPSYS_UNCONNECTED_386, SYNOPSYS_UNCONNECTED_387, 
        SYNOPSYS_UNCONNECTED_388}), .in1({1'b0, 1'b0, 1'b0, mulout11, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 1'b0, 1'b0, cout11, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in3({1'b1, 1'b0, 1'b1, 
        1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 
        1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .cout_46_(N50), .cout_44_(N48), .cout_42_(N46), .cout_40_(N44), .cout_38_(
        N42), .cout_36_(N40), .cout_34_(N38), .cout_32_(N36), .cout_30_(N34), 
        .cout_28_(N32), .cout_27_(N31), .cout_7__BAR(N11), .cout_8__BAR(N12), 
        .cout_9__BAR(N13), .cout_10__BAR(N14), .cout_11__BAR(N15), 
        .cout_12__BAR(N16), .cout_13__BAR(N17), .cout_14__BAR(N18), 
        .cout_15__BAR(N19), .cout_16__BAR(N20), .cout_17__BAR(N21), 
        .cout_18__BAR(N22), .cout_19__BAR(N23), .cout_20__BAR(N24), 
        .cout_21__BAR(N25), .cout_22__BAR(N26), .cout_23__BAR(N27), 
        .cout_24__BAR(N28), .cout_25__BAR(N29), .cout_26__BAR(N30), 
        .cout_29__BAR(N33), .cout_31__BAR(N35), .cout_33__BAR(N37), 
        .cout_35__BAR(N39), .cout_37__BAR(N41), .cout_39__BAR(N43), 
        .cout_41__BAR(N45), .cout_43__BAR(N47), .cout_45__BAR(N49) );
  cla51squ_3 cla51squ ( .out({SYNOPSYS_UNCONNECTED_389, 
        SYNOPSYS_UNCONNECTED_390, SYNOPSYS_UNCONNECTED_391, mulout[47:23], 
        SYNOPSYS_UNCONNECTED_392, SYNOPSYS_UNCONNECTED_393, 
        SYNOPSYS_UNCONNECTED_394, SYNOPSYS_UNCONNECTED_395, 
        SYNOPSYS_UNCONNECTED_396, SYNOPSYS_UNCONNECTED_397, 
        SYNOPSYS_UNCONNECTED_398, SYNOPSYS_UNCONNECTED_399, 
        SYNOPSYS_UNCONNECTED_400, SYNOPSYS_UNCONNECTED_401, 
        SYNOPSYS_UNCONNECTED_402, SYNOPSYS_UNCONNECTED_403, 
        SYNOPSYS_UNCONNECTED_404, SYNOPSYS_UNCONNECTED_405, 
        SYNOPSYS_UNCONNECTED_406, SYNOPSYS_UNCONNECTED_407, 
        SYNOPSYS_UNCONNECTED_408, SYNOPSYS_UNCONNECTED_409, 
        SYNOPSYS_UNCONNECTED_410, SYNOPSYS_UNCONNECTED_411, 
        SYNOPSYS_UNCONNECTED_412, SYNOPSYS_UNCONNECTED_413, 
        SYNOPSYS_UNCONNECTED_414}), .a({1'b0, 1'b0, 1'b0, a[47:8], 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({1'b0, 1'b0, 1'b0, b, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  DFFARX1 b_reg_47_ ( .D(N101), .CLK(clk), .RSTB(rst_n), .Q(b[47]) );
  DFFARX1 b_reg_46_ ( .D(N100), .CLK(clk), .RSTB(rst_n), .Q(b[46]) );
  DFFARX1 b_reg_45_ ( .D(N99), .CLK(clk), .RSTB(rst_n), .Q(b[45]) );
  DFFARX1 b_reg_44_ ( .D(N98), .CLK(clk), .RSTB(rst_n), .Q(b[44]) );
  DFFARX1 b_reg_43_ ( .D(N97), .CLK(clk), .RSTB(rst_n), .Q(b[43]) );
  DFFARX1 b_reg_42_ ( .D(N96), .CLK(clk), .RSTB(rst_n), .Q(b[42]) );
  DFFARX1 b_reg_41_ ( .D(N95), .CLK(clk), .RSTB(rst_n), .Q(b[41]) );
  DFFARX1 b_reg_40_ ( .D(N94), .CLK(clk), .RSTB(rst_n), .Q(b[40]) );
  DFFARX1 b_reg_39_ ( .D(N93), .CLK(clk), .RSTB(rst_n), .Q(b[39]) );
  DFFARX1 b_reg_38_ ( .D(N92), .CLK(clk), .RSTB(rst_n), .Q(b[38]) );
  DFFARX1 b_reg_37_ ( .D(N91), .CLK(clk), .RSTB(rst_n), .Q(b[37]) );
  DFFARX1 b_reg_36_ ( .D(N90), .CLK(clk), .RSTB(rst_n), .Q(b[36]) );
  DFFARX1 b_reg_35_ ( .D(N89), .CLK(clk), .RSTB(rst_n), .Q(b[35]) );
  DFFARX1 b_reg_34_ ( .D(N88), .CLK(clk), .RSTB(rst_n), .Q(b[34]) );
  DFFARX1 b_reg_33_ ( .D(N87), .CLK(clk), .RSTB(rst_n), .Q(b[33]) );
  DFFARX1 b_reg_32_ ( .D(N86), .CLK(clk), .RSTB(rst_n), .Q(b[32]) );
  DFFARX1 b_reg_31_ ( .D(N85), .CLK(clk), .RSTB(rst_n), .Q(b[31]) );
  DFFARX1 b_reg_30_ ( .D(N84), .CLK(clk), .RSTB(rst_n), .Q(b[30]) );
  DFFARX1 b_reg_29_ ( .D(N83), .CLK(clk), .RSTB(rst_n), .Q(b[29]) );
  DFFARX1 b_reg_28_ ( .D(N82), .CLK(clk), .RSTB(rst_n), .Q(b[28]) );
  DFFARX1 b_reg_27_ ( .D(N81), .CLK(clk), .RSTB(rst_n), .Q(b[27]) );
  DFFARX1 b_reg_26_ ( .D(N80), .CLK(clk), .RSTB(rst_n), .Q(b[26]) );
  DFFARX1 b_reg_25_ ( .D(N79), .CLK(clk), .RSTB(rst_n), .Q(b[25]) );
  DFFARX1 b_reg_24_ ( .D(N78), .CLK(clk), .RSTB(rst_n), .Q(b[24]) );
  DFFARX1 b_reg_23_ ( .D(N77), .CLK(clk), .RSTB(rst_n), .Q(b[23]) );
  DFFARX1 b_reg_22_ ( .D(N76), .CLK(clk), .RSTB(rst_n), .Q(b[22]) );
  DFFARX1 b_reg_21_ ( .D(N75), .CLK(clk), .RSTB(rst_n), .Q(b[21]) );
  DFFARX1 b_reg_20_ ( .D(N74), .CLK(clk), .RSTB(rst_n), .Q(b[20]) );
  DFFARX1 b_reg_19_ ( .D(N73), .CLK(clk), .RSTB(rst_n), .Q(b[19]) );
  DFFARX1 b_reg_18_ ( .D(N72), .CLK(clk), .RSTB(rst_n), .Q(b[18]) );
  DFFARX1 b_reg_17_ ( .D(N71), .CLK(clk), .RSTB(rst_n), .Q(b[17]) );
  DFFARX1 b_reg_16_ ( .D(N70), .CLK(clk), .RSTB(rst_n), .Q(b[16]) );
  DFFARX1 b_reg_15_ ( .D(N69), .CLK(clk), .RSTB(rst_n), .Q(b[15]) );
  DFFARX1 b_reg_14_ ( .D(N68), .CLK(clk), .RSTB(rst_n), .Q(b[14]) );
  DFFARX1 b_reg_13_ ( .D(N67), .CLK(clk), .RSTB(rst_n), .Q(b[13]) );
  DFFARX1 b_reg_12_ ( .D(N66), .CLK(clk), .RSTB(rst_n), .Q(b[12]) );
  DFFARX1 b_reg_11_ ( .D(N65), .CLK(clk), .RSTB(rst_n), .Q(b[11]) );
  DFFARX1 b_reg_10_ ( .D(N64), .CLK(clk), .RSTB(rst_n), .Q(b[10]) );
  DFFARX1 b_reg_9_ ( .D(N63), .CLK(clk), .RSTB(rst_n), .Q(b[9]) );
  DFFARX1 b_reg_8_ ( .D(N62), .CLK(clk), .RSTB(rst_n), .Q(b[8]) );
  DFFARX1 a_reg_47_ ( .D(N50), .CLK(clk), .RSTB(rst_n), .Q(a[47]) );
  DFFARX1 a_reg_46_ ( .D(n55), .CLK(clk), .RSTB(rst_n), .Q(a[46]) );
  DFFARX1 a_reg_45_ ( .D(N48), .CLK(clk), .RSTB(rst_n), .Q(a[45]) );
  DFFARX1 a_reg_44_ ( .D(n56), .CLK(clk), .RSTB(rst_n), .Q(a[44]) );
  DFFARX1 a_reg_43_ ( .D(N46), .CLK(clk), .RSTB(rst_n), .Q(a[43]) );
  DFFARX1 a_reg_42_ ( .D(n57), .CLK(clk), .RSTB(rst_n), .Q(a[42]) );
  DFFARX1 a_reg_41_ ( .D(N44), .CLK(clk), .RSTB(rst_n), .Q(a[41]) );
  DFFARX1 a_reg_40_ ( .D(n58), .CLK(clk), .RSTB(rst_n), .Q(a[40]) );
  DFFARX1 a_reg_39_ ( .D(N42), .CLK(clk), .RSTB(rst_n), .Q(a[39]) );
  DFFARX1 a_reg_38_ ( .D(n59), .CLK(clk), .RSTB(rst_n), .Q(a[38]) );
  DFFARX1 a_reg_37_ ( .D(N40), .CLK(clk), .RSTB(rst_n), .Q(a[37]) );
  DFFARX1 a_reg_36_ ( .D(n60), .CLK(clk), .RSTB(rst_n), .Q(a[36]) );
  DFFARX1 a_reg_35_ ( .D(N38), .CLK(clk), .RSTB(rst_n), .Q(a[35]) );
  DFFARX1 a_reg_34_ ( .D(n61), .CLK(clk), .RSTB(rst_n), .Q(a[34]) );
  DFFARX1 a_reg_33_ ( .D(N36), .CLK(clk), .RSTB(rst_n), .Q(a[33]) );
  DFFARX1 a_reg_32_ ( .D(n62), .CLK(clk), .RSTB(rst_n), .Q(a[32]) );
  DFFARX1 a_reg_31_ ( .D(N34), .CLK(clk), .RSTB(rst_n), .Q(a[31]) );
  DFFARX1 a_reg_30_ ( .D(n63), .CLK(clk), .RSTB(rst_n), .Q(a[30]) );
  DFFARX1 a_reg_29_ ( .D(N32), .CLK(clk), .RSTB(rst_n), .Q(a[29]) );
  DFFARX1 a_reg_28_ ( .D(N31), .CLK(clk), .RSTB(rst_n), .Q(a[28]) );
  DFFARX1 a_reg_27_ ( .D(n64), .CLK(clk), .RSTB(rst_n), .Q(a[27]) );
  DFFARX1 a_reg_26_ ( .D(n65), .CLK(clk), .RSTB(rst_n), .Q(a[26]) );
  DFFARX1 a_reg_25_ ( .D(n66), .CLK(clk), .RSTB(rst_n), .Q(a[25]) );
  DFFARX1 a_reg_24_ ( .D(n67), .CLK(clk), .RSTB(rst_n), .Q(a[24]) );
  DFFARX1 a_reg_23_ ( .D(n68), .CLK(clk), .RSTB(rst_n), .Q(a[23]) );
  DFFARX1 a_reg_22_ ( .D(n69), .CLK(clk), .RSTB(rst_n), .Q(a[22]) );
  DFFARX1 a_reg_21_ ( .D(n70), .CLK(clk), .RSTB(rst_n), .Q(a[21]) );
  DFFARX1 a_reg_20_ ( .D(n71), .CLK(clk), .RSTB(rst_n), .Q(a[20]) );
  DFFARX1 a_reg_19_ ( .D(n72), .CLK(clk), .RSTB(rst_n), .Q(a[19]) );
  DFFARX1 a_reg_18_ ( .D(n73), .CLK(clk), .RSTB(rst_n), .Q(a[18]) );
  DFFARX1 a_reg_17_ ( .D(n74), .CLK(clk), .RSTB(rst_n), .Q(a[17]) );
  DFFARX1 a_reg_16_ ( .D(n75), .CLK(clk), .RSTB(rst_n), .Q(a[16]) );
  DFFARX1 a_reg_15_ ( .D(n76), .CLK(clk), .RSTB(rst_n), .Q(a[15]) );
  DFFARX1 a_reg_14_ ( .D(n77), .CLK(clk), .RSTB(rst_n), .Q(a[14]) );
  DFFARX1 a_reg_13_ ( .D(n78), .CLK(clk), .RSTB(rst_n), .Q(a[13]) );
  DFFARX1 a_reg_12_ ( .D(n79), .CLK(clk), .RSTB(rst_n), .Q(a[12]) );
  DFFARX1 a_reg_11_ ( .D(n80), .CLK(clk), .RSTB(rst_n), .Q(a[11]) );
  DFFARX1 a_reg_10_ ( .D(n81), .CLK(clk), .RSTB(rst_n), .Q(a[10]) );
  DFFARX1 a_reg_9_ ( .D(n82), .CLK(clk), .RSTB(rst_n), .Q(a[9]) );
  DFFARX1 a_reg_8_ ( .D(n83), .CLK(clk), .RSTB(rst_n), .Q(a[8]) );
  INVX0 U5 ( .INP(boothout3[26]), .ZN(n125) );
  INVX0 U8 ( .INP(boothout6[26]), .ZN(n124) );
  NBUFFX8 U3 ( .INP(in2[18]), .Z(n25) );
  NBUFFX8 U4 ( .INP(in2[3]), .Z(n20) );
  NBUFFX8 U6 ( .INP(in2[9]), .Z(n21) );
  NBUFFX8 U7 ( .INP(in2[11]), .Z(n22) );
  NBUFFX8 U9 ( .INP(in2[15]), .Z(n24) );
  NBUFFX2 U10 ( .INP(in2[12]), .Z(n23) );
  NBUFFX8 U11 ( .INP(in2[1]), .Z(n19) );
  NBUFFX8 U12 ( .INP(in2[0]), .Z(n18) );
  INVX0 U64 ( .INP(N49), .ZN(n55) );
  INVX0 U65 ( .INP(N47), .ZN(n56) );
  INVX0 U66 ( .INP(N45), .ZN(n57) );
  INVX0 U67 ( .INP(N43), .ZN(n58) );
  INVX0 U68 ( .INP(N41), .ZN(n59) );
  INVX0 U69 ( .INP(N39), .ZN(n60) );
  INVX0 U70 ( .INP(N37), .ZN(n61) );
  INVX0 U71 ( .INP(N35), .ZN(n62) );
  INVX0 U72 ( .INP(N33), .ZN(n63) );
  INVX0 U73 ( .INP(N30), .ZN(n64) );
  INVX0 U74 ( .INP(N29), .ZN(n65) );
  INVX0 U75 ( .INP(N28), .ZN(n66) );
  INVX0 U76 ( .INP(N27), .ZN(n67) );
  INVX0 U77 ( .INP(N26), .ZN(n68) );
  INVX0 U78 ( .INP(N25), .ZN(n69) );
  INVX0 U79 ( .INP(N24), .ZN(n70) );
  INVX0 U80 ( .INP(N23), .ZN(n71) );
  INVX0 U81 ( .INP(N22), .ZN(n72) );
  INVX0 U82 ( .INP(N21), .ZN(n73) );
  INVX0 U83 ( .INP(N20), .ZN(n74) );
  INVX0 U84 ( .INP(N19), .ZN(n75) );
  INVX0 U85 ( .INP(N18), .ZN(n76) );
  INVX0 U86 ( .INP(N17), .ZN(n77) );
  INVX0 U87 ( .INP(N16), .ZN(n78) );
  INVX0 U88 ( .INP(N15), .ZN(n79) );
  INVX0 U89 ( .INP(N14), .ZN(n80) );
  INVX0 U90 ( .INP(N13), .ZN(n81) );
  INVX0 U91 ( .INP(N12), .ZN(n82) );
  INVX0 U92 ( .INP(N11), .ZN(n83) );
endmodule


module add_321 ( s, a, b, co, ci_BAR );
  input a, b, ci_BAR;
  output s, co;


  XOR2X1 U1 ( .IN1(a), .IN2(ci_BAR), .Q(s) );
endmodule


module add_322 ( s, a, b, ci, co_BAR );
  input a, b, ci;
  output s, co_BAR;


  NAND2X0 U1 ( .IN1(ci), .IN2(a), .QN(co_BAR) );
  OA21X1 U2 ( .IN1(ci), .IN2(a), .IN3(co_BAR), .Q(s) );
endmodule


module add_323 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_324 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_325 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_326 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(ci), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(ci), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module add_327 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  INVX0 U1 ( .INP(a), .ZN(s) );
  NBUFFX2 U2 ( .INP(a), .Z(co) );
endmodule


module add_328 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  NBUFFX2 U1 ( .INP(a), .Z(s) );
endmodule


module adder8_23 ( out, a, b, cin );
  output [7:0] out;
  input [7:0] a;
  input [7:0] b;
  input cin;

  wire   [6:1] c;

  add_328 add_01 ( .s(out[0]), .a(a[0]), .b(1'b1), .ci(1'b1) );
  add_327 add_02 ( .s(out[1]), .a(a[1]), .b(1'b0), .ci(1'b1), .co(c[1]) );
  add_326 add_03 ( .s(out[2]), .a(a[2]), .b(1'b0), .ci(c[1]), .co(c[2]) );
  add_325 add_04 ( .s(out[3]), .a(a[3]), .b(1'b0), .ci(c[2]), .co(c[3]) );
  add_324 add_05 ( .s(out[4]), .a(a[4]), .b(1'b0), .ci(c[3]), .co(c[4]) );
  add_323 add_06 ( .s(out[5]), .a(a[5]), .b(1'b0), .ci(c[4]), .co(c[5]) );
  add_322 add_07 ( .s(out[6]), .a(a[6]), .b(1'b0), .ci(c[5]), .co_BAR(c[6]) );
  add_321 add_08 ( .s(out[7]), .a(a[7]), .b(1'b1), .ci_BAR(c[6]) );
endmodule


module add_329 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  XOR2X1 U1 ( .IN1(ci), .IN2(b), .Q(s) );
endmodule


module add_330 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_331 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_332 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_333 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_334 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_335 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;


  FADDX1 U1 ( .A(a), .B(b), .CI(ci), .CO(co), .S(s) );
endmodule


module add_336 ( s, a, b, ci, co );
  input a, b, ci;
  output s, co;
  wire   n1;

  AND2X1 U1 ( .IN1(b), .IN2(a), .Q(co) );
  NOR2X0 U2 ( .IN1(b), .IN2(a), .QN(n1) );
  NOR2X0 U3 ( .IN1(n1), .IN2(co), .QN(s) );
endmodule


module adder8_24 ( out, a, b, cin );
  output [7:0] out;
  input [7:0] a;
  input [7:0] b;
  input cin;

  wire   [6:0] c;

  add_336 add_01 ( .s(out[0]), .a(a[0]), .b(b[0]), .ci(1'b0), .co(c[0]) );
  add_335 add_02 ( .s(out[1]), .a(a[1]), .b(b[1]), .ci(c[0]), .co(c[1]) );
  add_334 add_03 ( .s(out[2]), .a(a[2]), .b(b[2]), .ci(c[1]), .co(c[2]) );
  add_333 add_04 ( .s(out[3]), .a(a[3]), .b(b[3]), .ci(c[2]), .co(c[3]) );
  add_332 add_05 ( .s(out[4]), .a(a[4]), .b(b[4]), .ci(c[3]), .co(c[4]) );
  add_331 add_06 ( .s(out[5]), .a(a[5]), .b(b[5]), .ci(c[4]), .co(c[5]) );
  add_330 add_07 ( .s(out[6]), .a(a[6]), .b(b[6]), .ci(c[5]), .co(c[6]) );
  add_329 add_08 ( .s(out[7]), .a(1'b0), .b(b[7]), .ci(c[6]) );
endmodule


module floating_point_multiple_3 ( clk, rst_n, input_factor_01, 
        input_factor_02, output_multiply );
  input [31:0] input_factor_01;
  input [31:0] input_factor_02;
  output [31:0] output_multiply;
  input clk, rst_n;
  wire   N5, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22,
         N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N48, N49, N50, N51,
         N52, N53, N54, N55, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22,
         SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24,
         SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26;
  wire   [47:23] base_multiply_result;
  wire   [47:23] mulout;
  wire   [7:0] exponent_factor_12;
  wire   [7:0] pre_mul_output_exponent;

  mul26_3 mul26_01 ( .clk(clk), .rst_n(rst_n), .in1({1'b0, 1'b0, 1'b1, 
        input_factor_01[22:14], 1'b0, input_factor_01[12:7], 1'b0, 
        input_factor_01[5:0]}), .in2({1'b0, 1'b0, 1'b1, input_factor_02[22:7], 
        n3, input_factor_02[5:0]}), .en(1'b1), .mulout({SYNOPSYS_UNCONNECTED_1, 
        SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, mulout, 
        SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, 
        SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, 
        SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11, 
        SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13, 
        SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, 
        SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17, 
        SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19, 
        SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21, 
        SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_23, 
        SYNOPSYS_UNCONNECTED_24, SYNOPSYS_UNCONNECTED_25, 
        SYNOPSYS_UNCONNECTED_26}) );
  adder8_24 adder8_01 ( .out(exponent_factor_12), .a({1'b0, 
        input_factor_01[29:23]}), .b(input_factor_02[30:23]), .cin(1'b0) );
  adder8_23 adder8_02 ( .out(pre_mul_output_exponent), .a(exponent_factor_12), 
        .b({1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0}), .cin(1'b1) );
  DFFARX1 mul_output_sign_reg ( .D(N5), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[31]) );
  DFFARX1 base_multiply_result_reg_47_ ( .D(mulout[47]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[47]) );
  DFFARX1 base_multiply_result_reg_46_ ( .D(mulout[46]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[46]) );
  DFFARX1 base_multiply_result_reg_45_ ( .D(mulout[45]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[45]) );
  DFFARX1 base_multiply_result_reg_44_ ( .D(mulout[44]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[44]) );
  DFFARX1 base_multiply_result_reg_43_ ( .D(mulout[43]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[43]) );
  DFFARX1 base_multiply_result_reg_42_ ( .D(mulout[42]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[42]) );
  DFFARX1 base_multiply_result_reg_41_ ( .D(mulout[41]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[41]) );
  DFFARX1 base_multiply_result_reg_40_ ( .D(mulout[40]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[40]) );
  DFFARX1 base_multiply_result_reg_39_ ( .D(mulout[39]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[39]) );
  DFFARX1 base_multiply_result_reg_38_ ( .D(mulout[38]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[38]) );
  DFFARX1 base_multiply_result_reg_37_ ( .D(mulout[37]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[37]) );
  DFFARX1 base_multiply_result_reg_36_ ( .D(mulout[36]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[36]) );
  DFFARX1 base_multiply_result_reg_35_ ( .D(mulout[35]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[35]) );
  DFFARX1 base_multiply_result_reg_34_ ( .D(mulout[34]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[34]) );
  DFFARX1 base_multiply_result_reg_33_ ( .D(mulout[33]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[33]) );
  DFFARX1 base_multiply_result_reg_32_ ( .D(mulout[32]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[32]) );
  DFFARX1 base_multiply_result_reg_31_ ( .D(mulout[31]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[31]) );
  DFFARX1 base_multiply_result_reg_30_ ( .D(mulout[30]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[30]) );
  DFFARX1 base_multiply_result_reg_29_ ( .D(mulout[29]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[29]) );
  DFFARX1 base_multiply_result_reg_28_ ( .D(mulout[28]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[28]) );
  DFFARX1 base_multiply_result_reg_27_ ( .D(mulout[27]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[27]) );
  DFFARX1 base_multiply_result_reg_26_ ( .D(mulout[26]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[26]) );
  DFFARX1 base_multiply_result_reg_25_ ( .D(mulout[25]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[25]) );
  DFFARX1 base_multiply_result_reg_24_ ( .D(mulout[24]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[24]) );
  DFFARX1 base_multiply_result_reg_23_ ( .D(mulout[23]), .CLK(clk), .RSTB(
        rst_n), .Q(base_multiply_result[23]) );
  DFFARX1 mul_output_significand_reg_22_ ( .D(N32), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[22]) );
  DFFARX1 mul_output_significand_reg_21_ ( .D(N31), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[21]) );
  DFFARX1 mul_output_significand_reg_20_ ( .D(N30), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[20]) );
  DFFARX1 mul_output_significand_reg_19_ ( .D(N29), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[19]) );
  DFFARX1 mul_output_significand_reg_18_ ( .D(N28), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[18]) );
  DFFARX1 mul_output_significand_reg_17_ ( .D(N27), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[17]) );
  DFFARX1 mul_output_significand_reg_16_ ( .D(N26), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[16]) );
  DFFARX1 mul_output_significand_reg_15_ ( .D(N25), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[15]) );
  DFFARX1 mul_output_significand_reg_14_ ( .D(N24), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[14]) );
  DFFARX1 mul_output_significand_reg_13_ ( .D(N23), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[13]) );
  DFFARX1 mul_output_significand_reg_12_ ( .D(N22), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[12]) );
  DFFARX1 mul_output_significand_reg_11_ ( .D(N21), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[11]) );
  DFFARX1 mul_output_significand_reg_10_ ( .D(N20), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[10]) );
  DFFARX1 mul_output_significand_reg_9_ ( .D(N19), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[9]) );
  DFFARX1 mul_output_significand_reg_8_ ( .D(N18), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[8]) );
  DFFARX1 mul_output_significand_reg_7_ ( .D(N17), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[7]) );
  DFFARX1 mul_output_significand_reg_6_ ( .D(N16), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[6]) );
  DFFARX1 mul_output_significand_reg_5_ ( .D(N15), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[5]) );
  DFFARX1 mul_output_significand_reg_4_ ( .D(N14), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[4]) );
  DFFARX1 mul_output_significand_reg_3_ ( .D(N13), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[3]) );
  DFFARX1 mul_output_significand_reg_2_ ( .D(N12), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[2]) );
  DFFARX1 mul_output_significand_reg_1_ ( .D(N11), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[1]) );
  DFFARX1 mul_output_significand_reg_0_ ( .D(N10), .CLK(clk), .RSTB(rst_n), 
        .Q(output_multiply[0]) );
  DFFARX1 mul_output_exponent_reg_7_ ( .D(N55), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[30]) );
  DFFARX1 mul_output_exponent_reg_6_ ( .D(N54), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[29]) );
  DFFARX1 mul_output_exponent_reg_5_ ( .D(N53), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[28]) );
  DFFARX1 mul_output_exponent_reg_4_ ( .D(N52), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[27]) );
  DFFARX1 mul_output_exponent_reg_3_ ( .D(N51), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[26]) );
  DFFARX1 mul_output_exponent_reg_2_ ( .D(N50), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[25]) );
  DFFARX1 mul_output_exponent_reg_1_ ( .D(N49), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[24]) );
  DFFARX1 mul_output_exponent_reg_0_ ( .D(N48), .CLK(clk), .RSTB(rst_n), .Q(
        output_multiply[23]) );
  AND2X1 U3 ( .IN1(base_multiply_result[47]), .IN2(n36), .Q(n33) );
  INVX0 U4 ( .INP(n1), .ZN(n2) );
  OR2X1 U5 ( .IN1(base_multiply_result[47]), .IN2(n25), .Q(n1) );
  NBUFFX2 U6 ( .INP(input_factor_02[6]), .Z(n3) );
  INVX0 U7 ( .INP(input_factor_02[31]), .ZN(n4) );
  NOR4X0 U9 ( .IN1(input_factor_01[21]), .IN2(input_factor_01[23]), .IN3(
        input_factor_01[17]), .IN4(input_factor_01[18]), .QN(n8) );
  NOR4X0 U10 ( .IN1(input_factor_01[11]), .IN2(input_factor_01[12]), .IN3(
        input_factor_01[22]), .IN4(input_factor_01[20]), .QN(n7) );
  NOR4X0 U11 ( .IN1(input_factor_01[28]), .IN2(input_factor_01[15]), .IN3(
        input_factor_01[16]), .IN4(input_factor_01[14]), .QN(n6) );
  NOR4X0 U12 ( .IN1(input_factor_01[19]), .IN2(input_factor_01[2]), .IN3(
        input_factor_01[1]), .IN4(input_factor_01[29]), .QN(n5) );
  NAND4X0 U13 ( .IN1(n8), .IN2(n7), .IN3(n6), .IN4(n5), .QN(n24) );
  NOR4X0 U14 ( .IN1(input_factor_01[8]), .IN2(input_factor_01[9]), .IN3(
        input_factor_01[24]), .IN4(input_factor_01[25]), .QN(n12) );
  NOR4X0 U15 ( .IN1(input_factor_01[4]), .IN2(input_factor_01[5]), .IN3(
        input_factor_01[0]), .IN4(input_factor_01[10]), .QN(n11) );
  NOR4X0 U16 ( .IN1(input_factor_01[26]), .IN2(input_factor_01[27]), .IN3(
        input_factor_01[31]), .IN4(input_factor_01[3]), .QN(n10) );
  INVX0 U17 ( .INP(input_factor_01[7]), .ZN(n9) );
  NAND4X0 U18 ( .IN1(n12), .IN2(n11), .IN3(n10), .IN4(n9), .QN(n23) );
  NOR4X0 U19 ( .IN1(input_factor_02[0]), .IN2(input_factor_02[10]), .IN3(
        input_factor_02[11]), .IN4(input_factor_02[12]), .QN(n16) );
  NOR4X0 U20 ( .IN1(input_factor_02[13]), .IN2(input_factor_02[14]), .IN3(
        input_factor_02[15]), .IN4(input_factor_02[16]), .QN(n15) );
  NOR4X0 U21 ( .IN1(input_factor_02[17]), .IN2(input_factor_02[18]), .IN3(
        input_factor_02[19]), .IN4(input_factor_02[1]), .QN(n14) );
  NOR4X0 U22 ( .IN1(input_factor_02[20]), .IN2(input_factor_02[21]), .IN3(
        input_factor_02[22]), .IN4(input_factor_02[23]), .QN(n13) );
  NAND4X0 U23 ( .IN1(n16), .IN2(n15), .IN3(n14), .IN4(n13), .QN(n22) );
  NOR4X0 U24 ( .IN1(input_factor_02[24]), .IN2(input_factor_02[25]), .IN3(
        input_factor_02[26]), .IN4(input_factor_02[27]), .QN(n20) );
  NOR4X0 U25 ( .IN1(input_factor_02[28]), .IN2(input_factor_02[29]), .IN3(
        input_factor_02[2]), .IN4(input_factor_02[30]), .QN(n19) );
  NOR4X0 U26 ( .IN1(input_factor_02[31]), .IN2(input_factor_02[3]), .IN3(
        input_factor_02[4]), .IN4(input_factor_02[5]), .QN(n18) );
  NOR4X0 U27 ( .IN1(n3), .IN2(input_factor_02[7]), .IN3(input_factor_02[8]), 
        .IN4(input_factor_02[9]), .QN(n17) );
  NAND4X0 U28 ( .IN1(n20), .IN2(n19), .IN3(n18), .IN4(n17), .QN(n21) );
  OA22X1 U29 ( .IN1(n24), .IN2(n23), .IN3(n22), .IN4(n21), .Q(n36) );
  INVX0 U30 ( .INP(n36), .ZN(n25) );
  AO22X1 U31 ( .IN1(n2), .IN2(base_multiply_result[23]), .IN3(n33), .IN4(
        base_multiply_result[24]), .Q(N10) );
  AO22X1 U32 ( .IN1(n2), .IN2(base_multiply_result[24]), .IN3(n33), .IN4(
        base_multiply_result[25]), .Q(N11) );
  AO22X1 U33 ( .IN1(n2), .IN2(base_multiply_result[25]), .IN3(n33), .IN4(
        base_multiply_result[26]), .Q(N12) );
  AO22X1 U34 ( .IN1(n2), .IN2(base_multiply_result[26]), .IN3(n33), .IN4(
        base_multiply_result[27]), .Q(N13) );
  AO22X1 U35 ( .IN1(n2), .IN2(base_multiply_result[27]), .IN3(n33), .IN4(
        base_multiply_result[28]), .Q(N14) );
  AO22X1 U36 ( .IN1(n2), .IN2(base_multiply_result[28]), .IN3(n33), .IN4(
        base_multiply_result[29]), .Q(N15) );
  AO22X1 U37 ( .IN1(n2), .IN2(base_multiply_result[29]), .IN3(n33), .IN4(
        base_multiply_result[30]), .Q(N16) );
  AO22X1 U38 ( .IN1(n2), .IN2(base_multiply_result[30]), .IN3(n33), .IN4(
        base_multiply_result[31]), .Q(N17) );
  AO22X1 U39 ( .IN1(n2), .IN2(base_multiply_result[31]), .IN3(n33), .IN4(
        base_multiply_result[32]), .Q(N18) );
  AO22X1 U40 ( .IN1(n2), .IN2(base_multiply_result[32]), .IN3(n33), .IN4(
        base_multiply_result[33]), .Q(N19) );
  AO22X1 U41 ( .IN1(n2), .IN2(base_multiply_result[33]), .IN3(n33), .IN4(
        base_multiply_result[34]), .Q(N20) );
  AO22X1 U42 ( .IN1(n2), .IN2(base_multiply_result[34]), .IN3(n33), .IN4(
        base_multiply_result[35]), .Q(N21) );
  AO22X1 U43 ( .IN1(n2), .IN2(base_multiply_result[35]), .IN3(n33), .IN4(
        base_multiply_result[36]), .Q(N22) );
  AO22X1 U44 ( .IN1(n2), .IN2(base_multiply_result[36]), .IN3(n33), .IN4(
        base_multiply_result[37]), .Q(N23) );
  AO22X1 U45 ( .IN1(n2), .IN2(base_multiply_result[37]), .IN3(n33), .IN4(
        base_multiply_result[38]), .Q(N24) );
  AO22X1 U46 ( .IN1(n2), .IN2(base_multiply_result[38]), .IN3(n33), .IN4(
        base_multiply_result[39]), .Q(N25) );
  AO22X1 U47 ( .IN1(n2), .IN2(base_multiply_result[39]), .IN3(n33), .IN4(
        base_multiply_result[40]), .Q(N26) );
  AO22X1 U48 ( .IN1(n2), .IN2(base_multiply_result[40]), .IN3(n33), .IN4(
        base_multiply_result[41]), .Q(N27) );
  AO22X1 U49 ( .IN1(n2), .IN2(base_multiply_result[41]), .IN3(n33), .IN4(
        base_multiply_result[42]), .Q(N28) );
  AO22X1 U50 ( .IN1(n2), .IN2(base_multiply_result[42]), .IN3(n33), .IN4(
        base_multiply_result[43]), .Q(N29) );
  AO22X1 U51 ( .IN1(n2), .IN2(base_multiply_result[43]), .IN3(n33), .IN4(
        base_multiply_result[44]), .Q(N30) );
  AO22X1 U52 ( .IN1(n2), .IN2(base_multiply_result[44]), .IN3(n33), .IN4(
        base_multiply_result[45]), .Q(N31) );
  AO22X1 U53 ( .IN1(n2), .IN2(base_multiply_result[45]), .IN3(n33), .IN4(
        base_multiply_result[46]), .Q(N32) );
  MUX21X1 U54 ( .IN1(n2), .IN2(n33), .S(pre_mul_output_exponent[0]), .Q(N48)
         );
  AO21X1 U55 ( .IN1(pre_mul_output_exponent[0]), .IN2(n2), .IN3(n33), .Q(n26)
         );
  NOR3X0 U56 ( .IN1(pre_mul_output_exponent[1]), .IN2(
        pre_mul_output_exponent[0]), .IN3(n1), .QN(n28) );
  AO21X1 U57 ( .IN1(pre_mul_output_exponent[1]), .IN2(n26), .IN3(n28), .Q(N49)
         );
  INVX0 U58 ( .INP(input_factor_01[31]), .ZN(n27) );
  OA221X1 U59 ( .IN1(input_factor_01[31]), .IN2(input_factor_02[31]), .IN3(n27), .IN4(n4), .IN5(n36), .Q(N5) );
  AO221X1 U60 ( .IN1(n2), .IN2(pre_mul_output_exponent[1]), .IN3(n2), .IN4(
        pre_mul_output_exponent[0]), .IN5(n33), .Q(n29) );
  MUX21X1 U61 ( .IN1(n28), .IN2(n29), .S(pre_mul_output_exponent[2]), .Q(N50)
         );
  AND2X1 U62 ( .IN1(n2), .IN2(pre_mul_output_exponent[2]), .Q(n30) );
  OR4X1 U63 ( .IN1(pre_mul_output_exponent[1]), .IN2(
        pre_mul_output_exponent[0]), .IN3(pre_mul_output_exponent[3]), .IN4(
        pre_mul_output_exponent[2]), .Q(n35) );
  NOR2X0 U64 ( .IN1(n1), .IN2(n35), .QN(n32) );
  AO221X1 U65 ( .IN1(pre_mul_output_exponent[3]), .IN2(n30), .IN3(
        pre_mul_output_exponent[3]), .IN4(n29), .IN5(n32), .Q(N51) );
  OA21X1 U66 ( .IN1(base_multiply_result[47]), .IN2(n35), .IN3(n36), .Q(n31)
         );
  MUX21X1 U67 ( .IN1(n32), .IN2(n31), .S(pre_mul_output_exponent[4]), .Q(N52)
         );
  AO221X1 U68 ( .IN1(n2), .IN2(pre_mul_output_exponent[4]), .IN3(n2), .IN4(n35), .IN5(n33), .Q(n34) );
  NOR4X0 U69 ( .IN1(pre_mul_output_exponent[5]), .IN2(
        pre_mul_output_exponent[4]), .IN3(n35), .IN4(n1), .QN(n38) );
  AO21X1 U70 ( .IN1(pre_mul_output_exponent[5]), .IN2(n34), .IN3(n38), .Q(N53)
         );
  OR3X1 U71 ( .IN1(pre_mul_output_exponent[5]), .IN2(
        pre_mul_output_exponent[4]), .IN3(n35), .Q(n37) );
  OA21X1 U72 ( .IN1(base_multiply_result[47]), .IN2(n37), .IN3(n36), .Q(n40)
         );
  INVX0 U73 ( .INP(n38), .ZN(n39) );
  NOR2X0 U74 ( .IN1(pre_mul_output_exponent[6]), .IN2(n39), .QN(n42) );
  AO21X1 U75 ( .IN1(pre_mul_output_exponent[6]), .IN2(n40), .IN3(n42), .Q(N54)
         );
  AO21X1 U76 ( .IN1(n2), .IN2(pre_mul_output_exponent[6]), .IN3(n40), .Q(n41)
         );
  MUX21X1 U77 ( .IN1(n42), .IN2(n41), .S(pre_mul_output_exponent[7]), .Q(N55)
         );
endmodule


module tansigmoid_function ( clk, rst_n, tansigmoid_input, tansigmoid_output
 );
  input [31:0] tansigmoid_input;
  output [31:0] tansigmoid_output;
  input clk, rst_n;
  wire   n1, n2, n3, n4, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16;
  wire   [31:0] factor_a;
  wire   [31:0] factor_b;
  wire   [31:0] factor_c;
  wire   [31:0] factor_d;
  wire   [31:0] next_factor_a;
  wire   [31:0] next_factor_b;
  wire   [31:0] next_factor_c;
  wire   [31:0] next_factor_d;
  wire   [31:0] result_mult_b;
  wire   [31:0] next_result_mult_b;
  wire   [31:0] result_adder_b;
  wire   [31:0] next_result_adder_b;
  wire   [31:0] result_mult_c;
  wire   [31:0] next_result_mult_c;
  wire   [31:0] result_adder_c;
  wire   [31:0] next_result_adder_c;
  wire   [31:0] result_mult_d;
  wire   [31:0] next_result_mult_d;
  wire   [31:0] result_adder_d;

  tansigmoid_floating_point_compare floating_point_compare_01 ( .clk(clk), 
        .rst_n(rst_n), .factor_input({tansigmoid_input[31:11], n4, 
        tansigmoid_input[9], n3, tansigmoid_input[7:5], n2, 
        tansigmoid_input[3], n1, tansigmoid_input[1:0]}), .factor_a({
        factor_a[31], SYNOPSYS_UNCONNECTED_1, factor_a[29:14], 
        SYNOPSYS_UNCONNECTED_2, factor_a[12:7], SYNOPSYS_UNCONNECTED_3, 
        factor_a[5:0]}), .factor_b({factor_b[31], SYNOPSYS_UNCONNECTED_4, 
        factor_b[29:23], SYNOPSYS_UNCONNECTED_5, factor_b[21:20], 
        SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, factor_b[17:0]}), 
        .factor_c({factor_c[31], SYNOPSYS_UNCONNECTED_8, factor_c[29:21], 
        SYNOPSYS_UNCONNECTED_9, factor_c[19:13], SYNOPSYS_UNCONNECTED_10, 
        factor_c[11:2], SYNOPSYS_UNCONNECTED_11, factor_c[0]}), .factor_d({
        factor_d[31], SYNOPSYS_UNCONNECTED_12, factor_d[29], 
        SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14, 
        SYNOPSYS_UNCONNECTED_15, factor_d[25:24], SYNOPSYS_UNCONNECTED_16, 
        factor_d[22:0]}) );
  floating_point_multiple_3 multiple_01 ( .clk(clk), .rst_n(rst_n), 
        .input_factor_01({next_factor_a[31], 1'b0, next_factor_a[29:14], 1'b0, 
        next_factor_a[12:7], 1'b0, next_factor_a[5:0]}), .input_factor_02({
        tansigmoid_input[31:11], n4, tansigmoid_input[9], n3, 
        tansigmoid_input[7:5], n2, tansigmoid_input[3], n1, 
        tansigmoid_input[1:0]}), .output_multiply(result_mult_b) );
  floating_point_adder_3 adder_01 ( .clk(clk), .rst_n(rst_n), 
        .input_factor_01(next_result_mult_b), .input_factor_02({
        next_factor_b[31], 1'b0, next_factor_b[29:23], 1'b0, 
        next_factor_b[21:20], 1'b0, 1'b0, next_factor_b[17:0]}), 
        .output_adder(result_adder_b) );
  floating_point_multiple_2 multiple_02 ( .clk(clk), .rst_n(rst_n), 
        .input_factor_01(next_result_adder_b), .input_factor_02({
        tansigmoid_input[31:11], n4, tansigmoid_input[9], n3, 
        tansigmoid_input[7:5], n2, tansigmoid_input[3], n1, 
        tansigmoid_input[1:0]}), .output_multiply(result_mult_c) );
  floating_point_adder_2 adder_02 ( .clk(clk), .rst_n(rst_n), 
        .input_factor_01(next_result_mult_c), .input_factor_02({
        next_factor_c[31], 1'b0, next_factor_c[29:21], 1'b0, 
        next_factor_c[19:13], 1'b0, next_factor_c[11:2], 1'b0, 
        next_factor_c[0]}), .output_adder(result_adder_c) );
  floating_point_multiple_1 multiple_03 ( .clk(clk), .rst_n(rst_n), 
        .input_factor_01(next_result_adder_c), .input_factor_02({
        tansigmoid_input[31:11], n4, tansigmoid_input[9], n3, 
        tansigmoid_input[7:5], n2, tansigmoid_input[3], n1, 
        tansigmoid_input[1:0]}), .output_multiply(result_mult_d) );
  floating_point_adder_1 adder_03 ( .clk(clk), .rst_n(rst_n), 
        .input_factor_01(next_result_mult_d), .input_factor_02({
        next_factor_d[31], 1'b0, next_factor_d[29], next_factor_d[29], 
        next_factor_d[29], next_factor_d[29], next_factor_d[25:24], 
        next_factor_d[25], next_factor_d[22:0]}), .output_adder(result_adder_d) );
  DFFARX1 next_factor_a_reg_31_ ( .D(factor_a[31]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_a[31]) );
  DFFARX1 next_factor_a_reg_29_ ( .D(factor_a[29]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_a[29]) );
  DFFARX1 next_factor_a_reg_28_ ( .D(factor_a[28]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_a[28]) );
  DFFARX1 next_factor_a_reg_27_ ( .D(factor_a[27]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_a[27]) );
  DFFARX1 next_factor_a_reg_26_ ( .D(factor_a[26]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_a[26]) );
  DFFARX1 next_factor_a_reg_25_ ( .D(factor_a[25]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_a[25]) );
  DFFARX1 next_factor_a_reg_24_ ( .D(factor_a[24]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_a[24]) );
  DFFARX1 next_factor_a_reg_23_ ( .D(factor_a[23]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_a[23]) );
  DFFARX1 next_factor_a_reg_22_ ( .D(factor_a[22]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_a[22]) );
  DFFARX1 next_factor_a_reg_21_ ( .D(factor_a[21]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_a[21]) );
  DFFARX1 next_factor_a_reg_20_ ( .D(factor_a[20]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_a[20]) );
  DFFARX1 next_factor_a_reg_19_ ( .D(factor_a[19]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_a[19]) );
  DFFARX1 next_factor_a_reg_18_ ( .D(factor_a[18]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_a[18]) );
  DFFARX1 next_factor_a_reg_17_ ( .D(factor_a[17]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_a[17]) );
  DFFARX1 next_factor_a_reg_16_ ( .D(factor_a[16]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_a[16]) );
  DFFARX1 next_factor_a_reg_15_ ( .D(factor_a[15]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_a[15]) );
  DFFARX1 next_factor_a_reg_14_ ( .D(factor_a[14]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_a[14]) );
  DFFARX1 next_factor_a_reg_12_ ( .D(factor_a[12]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_a[12]) );
  DFFARX1 next_factor_a_reg_11_ ( .D(factor_a[11]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_a[11]) );
  DFFARX1 next_factor_a_reg_10_ ( .D(factor_a[10]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_a[10]) );
  DFFARX1 next_factor_a_reg_9_ ( .D(factor_a[9]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_a[9]) );
  DFFARX1 next_factor_a_reg_8_ ( .D(factor_a[8]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_a[8]) );
  DFFARX1 next_factor_a_reg_7_ ( .D(factor_a[7]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_a[7]) );
  DFFARX1 next_factor_a_reg_5_ ( .D(factor_a[5]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_a[5]) );
  DFFARX1 next_factor_a_reg_4_ ( .D(factor_a[4]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_a[4]) );
  DFFARX1 next_factor_a_reg_3_ ( .D(factor_a[3]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_a[3]) );
  DFFARX1 next_factor_a_reg_2_ ( .D(factor_a[2]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_a[2]) );
  DFFARX1 next_factor_a_reg_1_ ( .D(factor_a[1]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_a[1]) );
  DFFARX1 next_factor_a_reg_0_ ( .D(factor_a[0]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_a[0]) );
  DFFARX1 next_factor_b_reg_31_ ( .D(factor_b[31]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_b[31]) );
  DFFARX1 next_factor_b_reg_29_ ( .D(factor_b[29]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_b[29]) );
  DFFARX1 next_factor_b_reg_28_ ( .D(factor_b[28]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_b[28]) );
  DFFARX1 next_factor_b_reg_27_ ( .D(factor_b[27]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_b[27]) );
  DFFARX1 next_factor_b_reg_26_ ( .D(factor_b[26]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_b[26]) );
  DFFARX1 next_factor_b_reg_25_ ( .D(factor_b[25]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_b[25]) );
  DFFARX1 next_factor_b_reg_24_ ( .D(factor_b[24]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_b[24]) );
  DFFARX1 next_factor_b_reg_23_ ( .D(factor_b[23]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_b[23]) );
  DFFARX1 next_factor_b_reg_21_ ( .D(factor_b[21]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_b[21]) );
  DFFARX1 next_factor_b_reg_20_ ( .D(factor_b[20]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_b[20]) );
  DFFARX1 next_factor_b_reg_17_ ( .D(factor_b[17]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_b[17]) );
  DFFARX1 next_factor_b_reg_16_ ( .D(factor_b[16]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_b[16]) );
  DFFARX1 next_factor_b_reg_15_ ( .D(factor_b[15]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_b[15]) );
  DFFARX1 next_factor_b_reg_14_ ( .D(factor_b[14]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_b[14]) );
  DFFARX1 next_factor_b_reg_13_ ( .D(factor_b[13]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_b[13]) );
  DFFARX1 next_factor_b_reg_12_ ( .D(factor_b[12]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_b[12]) );
  DFFARX1 next_factor_b_reg_11_ ( .D(factor_b[11]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_b[11]) );
  DFFARX1 next_factor_b_reg_10_ ( .D(factor_b[10]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_b[10]) );
  DFFARX1 next_factor_b_reg_9_ ( .D(factor_b[9]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_b[9]) );
  DFFARX1 next_factor_b_reg_8_ ( .D(factor_b[8]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_b[8]) );
  DFFARX1 next_factor_b_reg_7_ ( .D(factor_b[7]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_b[7]) );
  DFFARX1 next_factor_b_reg_6_ ( .D(factor_b[6]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_b[6]) );
  DFFARX1 next_factor_b_reg_5_ ( .D(factor_b[5]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_b[5]) );
  DFFARX1 next_factor_b_reg_4_ ( .D(factor_b[4]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_b[4]) );
  DFFARX1 next_factor_b_reg_3_ ( .D(factor_b[3]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_b[3]) );
  DFFARX1 next_factor_b_reg_2_ ( .D(factor_b[2]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_b[2]) );
  DFFARX1 next_factor_b_reg_1_ ( .D(factor_b[1]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_b[1]) );
  DFFARX1 next_factor_b_reg_0_ ( .D(factor_b[0]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_b[0]) );
  DFFARX1 next_factor_c_reg_31_ ( .D(factor_c[31]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_c[31]) );
  DFFARX1 next_factor_c_reg_29_ ( .D(factor_c[29]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_c[29]) );
  DFFARX1 next_factor_c_reg_28_ ( .D(factor_c[28]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_c[28]) );
  DFFARX1 next_factor_c_reg_27_ ( .D(factor_c[27]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_c[27]) );
  DFFARX1 next_factor_c_reg_26_ ( .D(factor_c[26]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_c[26]) );
  DFFARX1 next_factor_c_reg_25_ ( .D(factor_c[25]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_c[25]) );
  DFFARX1 next_factor_c_reg_24_ ( .D(factor_c[24]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_c[24]) );
  DFFARX1 next_factor_c_reg_23_ ( .D(factor_c[23]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_c[23]) );
  DFFARX1 next_factor_c_reg_22_ ( .D(factor_c[22]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_c[22]) );
  DFFARX1 next_factor_c_reg_21_ ( .D(factor_c[21]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_c[21]) );
  DFFARX1 next_factor_c_reg_19_ ( .D(factor_c[19]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_c[19]) );
  DFFARX1 next_factor_c_reg_18_ ( .D(factor_c[18]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_c[18]) );
  DFFARX1 next_factor_c_reg_17_ ( .D(factor_c[17]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_c[17]) );
  DFFARX1 next_factor_c_reg_16_ ( .D(factor_c[16]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_c[16]) );
  DFFARX1 next_factor_c_reg_15_ ( .D(factor_c[15]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_c[15]) );
  DFFARX1 next_factor_c_reg_14_ ( .D(factor_c[14]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_c[14]) );
  DFFARX1 next_factor_c_reg_13_ ( .D(factor_c[13]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_c[13]) );
  DFFARX1 next_factor_c_reg_11_ ( .D(factor_c[11]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_c[11]) );
  DFFARX1 next_factor_c_reg_10_ ( .D(factor_c[10]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_c[10]) );
  DFFARX1 next_factor_c_reg_9_ ( .D(factor_c[9]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_c[9]) );
  DFFARX1 next_factor_c_reg_8_ ( .D(factor_c[8]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_c[8]) );
  DFFARX1 next_factor_c_reg_7_ ( .D(factor_c[7]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_c[7]) );
  DFFARX1 next_factor_c_reg_6_ ( .D(factor_c[6]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_c[6]) );
  DFFARX1 next_factor_c_reg_5_ ( .D(factor_c[5]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_c[5]) );
  DFFARX1 next_factor_c_reg_4_ ( .D(factor_c[4]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_c[4]) );
  DFFARX1 next_factor_c_reg_3_ ( .D(factor_c[3]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_c[3]) );
  DFFARX1 next_factor_c_reg_2_ ( .D(factor_c[2]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_c[2]) );
  DFFARX1 next_factor_c_reg_0_ ( .D(factor_c[0]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_c[0]) );
  DFFARX1 next_factor_d_reg_31_ ( .D(factor_d[31]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_d[31]) );
  DFFARX1 next_factor_d_reg_29_ ( .D(factor_d[29]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_d[29]) );
  DFFARX1 next_factor_d_reg_25_ ( .D(factor_d[25]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_d[25]) );
  DFFARX1 next_factor_d_reg_24_ ( .D(factor_d[24]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_d[24]) );
  DFFARX1 next_factor_d_reg_22_ ( .D(factor_d[22]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_d[22]) );
  DFFARX1 next_factor_d_reg_21_ ( .D(factor_d[21]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_d[21]) );
  DFFARX1 next_factor_d_reg_20_ ( .D(factor_d[20]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_d[20]) );
  DFFARX1 next_factor_d_reg_19_ ( .D(factor_d[19]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_d[19]) );
  DFFARX1 next_factor_d_reg_18_ ( .D(factor_d[18]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_d[18]) );
  DFFARX1 next_factor_d_reg_17_ ( .D(factor_d[17]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_d[17]) );
  DFFARX1 next_factor_d_reg_16_ ( .D(factor_d[16]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_d[16]) );
  DFFARX1 next_factor_d_reg_15_ ( .D(factor_d[15]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_d[15]) );
  DFFARX1 next_factor_d_reg_14_ ( .D(factor_d[14]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_d[14]) );
  DFFARX1 next_factor_d_reg_13_ ( .D(factor_d[13]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_d[13]) );
  DFFARX1 next_factor_d_reg_12_ ( .D(factor_d[12]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_d[12]) );
  DFFARX1 next_factor_d_reg_11_ ( .D(factor_d[11]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_d[11]) );
  DFFARX1 next_factor_d_reg_10_ ( .D(factor_d[10]), .CLK(clk), .RSTB(rst_n), 
        .Q(next_factor_d[10]) );
  DFFARX1 next_factor_d_reg_9_ ( .D(factor_d[9]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_d[9]) );
  DFFARX1 next_factor_d_reg_8_ ( .D(factor_d[8]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_d[8]) );
  DFFARX1 next_factor_d_reg_7_ ( .D(factor_d[7]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_d[7]) );
  DFFARX1 next_factor_d_reg_6_ ( .D(factor_d[6]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_d[6]) );
  DFFARX1 next_factor_d_reg_5_ ( .D(factor_d[5]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_d[5]) );
  DFFARX1 next_factor_d_reg_4_ ( .D(factor_d[4]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_d[4]) );
  DFFARX1 next_factor_d_reg_3_ ( .D(factor_d[3]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_d[3]) );
  DFFARX1 next_factor_d_reg_2_ ( .D(factor_d[2]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_d[2]) );
  DFFARX1 next_factor_d_reg_1_ ( .D(factor_d[1]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_d[1]) );
  DFFARX1 next_factor_d_reg_0_ ( .D(factor_d[0]), .CLK(clk), .RSTB(rst_n), .Q(
        next_factor_d[0]) );
  DFFARX1 next_result_mult_b_reg_31_ ( .D(result_mult_b[31]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_b[31]) );
  DFFARX1 next_result_mult_b_reg_30_ ( .D(result_mult_b[30]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_b[30]) );
  DFFARX1 next_result_mult_b_reg_29_ ( .D(result_mult_b[29]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_b[29]) );
  DFFARX1 next_result_mult_b_reg_28_ ( .D(result_mult_b[28]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_b[28]) );
  DFFARX1 next_result_mult_b_reg_27_ ( .D(result_mult_b[27]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_b[27]) );
  DFFARX1 next_result_mult_b_reg_26_ ( .D(result_mult_b[26]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_b[26]) );
  DFFARX1 next_result_mult_b_reg_25_ ( .D(result_mult_b[25]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_b[25]) );
  DFFARX1 next_result_mult_b_reg_24_ ( .D(result_mult_b[24]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_b[24]) );
  DFFARX1 next_result_mult_b_reg_23_ ( .D(result_mult_b[23]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_b[23]) );
  DFFARX1 next_result_mult_b_reg_22_ ( .D(result_mult_b[22]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_b[22]) );
  DFFARX1 next_result_mult_b_reg_21_ ( .D(result_mult_b[21]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_b[21]) );
  DFFARX1 next_result_mult_b_reg_20_ ( .D(result_mult_b[20]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_b[20]) );
  DFFARX1 next_result_mult_b_reg_19_ ( .D(result_mult_b[19]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_b[19]) );
  DFFARX1 next_result_mult_b_reg_18_ ( .D(result_mult_b[18]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_b[18]) );
  DFFARX1 next_result_mult_b_reg_17_ ( .D(result_mult_b[17]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_b[17]) );
  DFFARX1 next_result_mult_b_reg_16_ ( .D(result_mult_b[16]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_b[16]) );
  DFFARX1 next_result_mult_b_reg_15_ ( .D(result_mult_b[15]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_b[15]) );
  DFFARX1 next_result_mult_b_reg_14_ ( .D(result_mult_b[14]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_b[14]) );
  DFFARX1 next_result_mult_b_reg_13_ ( .D(result_mult_b[13]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_b[13]) );
  DFFARX1 next_result_mult_b_reg_12_ ( .D(result_mult_b[12]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_b[12]) );
  DFFARX1 next_result_mult_b_reg_11_ ( .D(result_mult_b[11]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_b[11]) );
  DFFARX1 next_result_mult_b_reg_10_ ( .D(result_mult_b[10]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_b[10]) );
  DFFARX1 next_result_mult_b_reg_9_ ( .D(result_mult_b[9]), .CLK(clk), .RSTB(
        rst_n), .Q(next_result_mult_b[9]) );
  DFFARX1 next_result_mult_b_reg_8_ ( .D(result_mult_b[8]), .CLK(clk), .RSTB(
        rst_n), .Q(next_result_mult_b[8]) );
  DFFARX1 next_result_mult_b_reg_7_ ( .D(result_mult_b[7]), .CLK(clk), .RSTB(
        rst_n), .Q(next_result_mult_b[7]) );
  DFFARX1 next_result_mult_b_reg_6_ ( .D(result_mult_b[6]), .CLK(clk), .RSTB(
        rst_n), .Q(next_result_mult_b[6]) );
  DFFARX1 next_result_mult_b_reg_5_ ( .D(result_mult_b[5]), .CLK(clk), .RSTB(
        rst_n), .Q(next_result_mult_b[5]) );
  DFFARX1 next_result_mult_b_reg_4_ ( .D(result_mult_b[4]), .CLK(clk), .RSTB(
        rst_n), .Q(next_result_mult_b[4]) );
  DFFARX1 next_result_mult_b_reg_3_ ( .D(result_mult_b[3]), .CLK(clk), .RSTB(
        rst_n), .Q(next_result_mult_b[3]) );
  DFFARX1 next_result_mult_b_reg_2_ ( .D(result_mult_b[2]), .CLK(clk), .RSTB(
        rst_n), .Q(next_result_mult_b[2]) );
  DFFARX1 next_result_mult_b_reg_1_ ( .D(result_mult_b[1]), .CLK(clk), .RSTB(
        rst_n), .Q(next_result_mult_b[1]) );
  DFFARX1 next_result_mult_b_reg_0_ ( .D(result_mult_b[0]), .CLK(clk), .RSTB(
        rst_n), .Q(next_result_mult_b[0]) );
  DFFARX1 next_result_adder_b_reg_31_ ( .D(result_adder_b[31]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[31]) );
  DFFARX1 next_result_adder_b_reg_30_ ( .D(result_adder_b[30]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[30]) );
  DFFARX1 next_result_adder_b_reg_29_ ( .D(result_adder_b[29]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[29]) );
  DFFARX1 next_result_adder_b_reg_28_ ( .D(result_adder_b[28]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[28]) );
  DFFARX1 next_result_adder_b_reg_27_ ( .D(result_adder_b[27]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[27]) );
  DFFARX1 next_result_adder_b_reg_26_ ( .D(result_adder_b[26]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[26]) );
  DFFARX1 next_result_adder_b_reg_25_ ( .D(result_adder_b[25]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[25]) );
  DFFARX1 next_result_adder_b_reg_24_ ( .D(result_adder_b[24]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[24]) );
  DFFARX1 next_result_adder_b_reg_23_ ( .D(result_adder_b[23]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[23]) );
  DFFARX1 next_result_adder_b_reg_22_ ( .D(result_adder_b[22]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[22]) );
  DFFARX1 next_result_adder_b_reg_21_ ( .D(result_adder_b[21]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[21]) );
  DFFARX1 next_result_adder_b_reg_20_ ( .D(result_adder_b[20]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[20]) );
  DFFARX1 next_result_adder_b_reg_19_ ( .D(result_adder_b[19]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[19]) );
  DFFARX1 next_result_adder_b_reg_18_ ( .D(result_adder_b[18]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[18]) );
  DFFARX1 next_result_adder_b_reg_17_ ( .D(result_adder_b[17]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[17]) );
  DFFARX1 next_result_adder_b_reg_16_ ( .D(result_adder_b[16]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[16]) );
  DFFARX1 next_result_adder_b_reg_15_ ( .D(result_adder_b[15]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[15]) );
  DFFARX1 next_result_adder_b_reg_14_ ( .D(result_adder_b[14]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[14]) );
  DFFARX1 next_result_adder_b_reg_13_ ( .D(result_adder_b[13]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[13]) );
  DFFARX1 next_result_adder_b_reg_12_ ( .D(result_adder_b[12]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[12]) );
  DFFARX1 next_result_adder_b_reg_11_ ( .D(result_adder_b[11]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[11]) );
  DFFARX1 next_result_adder_b_reg_10_ ( .D(result_adder_b[10]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[10]) );
  DFFARX1 next_result_adder_b_reg_9_ ( .D(result_adder_b[9]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[9]) );
  DFFARX1 next_result_adder_b_reg_8_ ( .D(result_adder_b[8]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[8]) );
  DFFARX1 next_result_adder_b_reg_7_ ( .D(result_adder_b[7]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[7]) );
  DFFARX1 next_result_adder_b_reg_6_ ( .D(result_adder_b[6]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[6]) );
  DFFARX1 next_result_adder_b_reg_5_ ( .D(result_adder_b[5]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[5]) );
  DFFARX1 next_result_adder_b_reg_4_ ( .D(result_adder_b[4]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[4]) );
  DFFARX1 next_result_adder_b_reg_3_ ( .D(result_adder_b[3]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[3]) );
  DFFARX1 next_result_adder_b_reg_2_ ( .D(result_adder_b[2]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[2]) );
  DFFARX1 next_result_adder_b_reg_1_ ( .D(result_adder_b[1]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[1]) );
  DFFARX1 next_result_adder_b_reg_0_ ( .D(result_adder_b[0]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_b[0]) );
  DFFARX1 next_result_mult_c_reg_31_ ( .D(result_mult_c[31]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_c[31]) );
  DFFARX1 next_result_mult_c_reg_30_ ( .D(result_mult_c[30]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_c[30]) );
  DFFARX1 next_result_mult_c_reg_29_ ( .D(result_mult_c[29]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_c[29]) );
  DFFARX1 next_result_mult_c_reg_28_ ( .D(result_mult_c[28]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_c[28]) );
  DFFARX1 next_result_mult_c_reg_27_ ( .D(result_mult_c[27]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_c[27]) );
  DFFARX1 next_result_mult_c_reg_26_ ( .D(result_mult_c[26]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_c[26]) );
  DFFARX1 next_result_mult_c_reg_25_ ( .D(result_mult_c[25]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_c[25]) );
  DFFARX1 next_result_mult_c_reg_24_ ( .D(result_mult_c[24]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_c[24]) );
  DFFARX1 next_result_mult_c_reg_23_ ( .D(result_mult_c[23]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_c[23]) );
  DFFARX1 next_result_mult_c_reg_22_ ( .D(result_mult_c[22]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_c[22]) );
  DFFARX1 next_result_mult_c_reg_21_ ( .D(result_mult_c[21]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_c[21]) );
  DFFARX1 next_result_mult_c_reg_20_ ( .D(result_mult_c[20]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_c[20]) );
  DFFARX1 next_result_mult_c_reg_19_ ( .D(result_mult_c[19]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_c[19]) );
  DFFARX1 next_result_mult_c_reg_18_ ( .D(result_mult_c[18]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_c[18]) );
  DFFARX1 next_result_mult_c_reg_17_ ( .D(result_mult_c[17]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_c[17]) );
  DFFARX1 next_result_mult_c_reg_16_ ( .D(result_mult_c[16]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_c[16]) );
  DFFARX1 next_result_mult_c_reg_15_ ( .D(result_mult_c[15]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_c[15]) );
  DFFARX1 next_result_mult_c_reg_14_ ( .D(result_mult_c[14]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_c[14]) );
  DFFARX1 next_result_mult_c_reg_13_ ( .D(result_mult_c[13]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_c[13]) );
  DFFARX1 next_result_mult_c_reg_12_ ( .D(result_mult_c[12]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_c[12]) );
  DFFARX1 next_result_mult_c_reg_11_ ( .D(result_mult_c[11]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_c[11]) );
  DFFARX1 next_result_mult_c_reg_10_ ( .D(result_mult_c[10]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_c[10]) );
  DFFARX1 next_result_mult_c_reg_9_ ( .D(result_mult_c[9]), .CLK(clk), .RSTB(
        rst_n), .Q(next_result_mult_c[9]) );
  DFFARX1 next_result_mult_c_reg_8_ ( .D(result_mult_c[8]), .CLK(clk), .RSTB(
        rst_n), .Q(next_result_mult_c[8]) );
  DFFARX1 next_result_mult_c_reg_7_ ( .D(result_mult_c[7]), .CLK(clk), .RSTB(
        rst_n), .Q(next_result_mult_c[7]) );
  DFFARX1 next_result_mult_c_reg_6_ ( .D(result_mult_c[6]), .CLK(clk), .RSTB(
        rst_n), .Q(next_result_mult_c[6]) );
  DFFARX1 next_result_mult_c_reg_5_ ( .D(result_mult_c[5]), .CLK(clk), .RSTB(
        rst_n), .Q(next_result_mult_c[5]) );
  DFFARX1 next_result_mult_c_reg_4_ ( .D(result_mult_c[4]), .CLK(clk), .RSTB(
        rst_n), .Q(next_result_mult_c[4]) );
  DFFARX1 next_result_mult_c_reg_3_ ( .D(result_mult_c[3]), .CLK(clk), .RSTB(
        rst_n), .Q(next_result_mult_c[3]) );
  DFFARX1 next_result_mult_c_reg_2_ ( .D(result_mult_c[2]), .CLK(clk), .RSTB(
        rst_n), .Q(next_result_mult_c[2]) );
  DFFARX1 next_result_mult_c_reg_1_ ( .D(result_mult_c[1]), .CLK(clk), .RSTB(
        rst_n), .Q(next_result_mult_c[1]) );
  DFFARX1 next_result_mult_c_reg_0_ ( .D(result_mult_c[0]), .CLK(clk), .RSTB(
        rst_n), .Q(next_result_mult_c[0]) );
  DFFARX1 next_result_adder_c_reg_31_ ( .D(result_adder_c[31]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[31]) );
  DFFARX1 next_result_adder_c_reg_30_ ( .D(result_adder_c[30]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[30]) );
  DFFARX1 next_result_adder_c_reg_29_ ( .D(result_adder_c[29]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[29]) );
  DFFARX1 next_result_adder_c_reg_28_ ( .D(result_adder_c[28]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[28]) );
  DFFARX1 next_result_adder_c_reg_27_ ( .D(result_adder_c[27]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[27]) );
  DFFARX1 next_result_adder_c_reg_26_ ( .D(result_adder_c[26]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[26]) );
  DFFARX1 next_result_adder_c_reg_25_ ( .D(result_adder_c[25]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[25]) );
  DFFARX1 next_result_adder_c_reg_24_ ( .D(result_adder_c[24]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[24]) );
  DFFARX1 next_result_adder_c_reg_23_ ( .D(result_adder_c[23]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[23]) );
  DFFARX1 next_result_adder_c_reg_22_ ( .D(result_adder_c[22]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[22]) );
  DFFARX1 next_result_adder_c_reg_21_ ( .D(result_adder_c[21]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[21]) );
  DFFARX1 next_result_adder_c_reg_20_ ( .D(result_adder_c[20]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[20]) );
  DFFARX1 next_result_adder_c_reg_19_ ( .D(result_adder_c[19]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[19]) );
  DFFARX1 next_result_adder_c_reg_18_ ( .D(result_adder_c[18]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[18]) );
  DFFARX1 next_result_adder_c_reg_17_ ( .D(result_adder_c[17]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[17]) );
  DFFARX1 next_result_adder_c_reg_16_ ( .D(result_adder_c[16]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[16]) );
  DFFARX1 next_result_adder_c_reg_15_ ( .D(result_adder_c[15]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[15]) );
  DFFARX1 next_result_adder_c_reg_14_ ( .D(result_adder_c[14]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[14]) );
  DFFARX1 next_result_adder_c_reg_13_ ( .D(result_adder_c[13]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[13]) );
  DFFARX1 next_result_adder_c_reg_12_ ( .D(result_adder_c[12]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[12]) );
  DFFARX1 next_result_adder_c_reg_11_ ( .D(result_adder_c[11]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[11]) );
  DFFARX1 next_result_adder_c_reg_10_ ( .D(result_adder_c[10]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[10]) );
  DFFARX1 next_result_adder_c_reg_9_ ( .D(result_adder_c[9]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[9]) );
  DFFARX1 next_result_adder_c_reg_8_ ( .D(result_adder_c[8]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[8]) );
  DFFARX1 next_result_adder_c_reg_7_ ( .D(result_adder_c[7]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[7]) );
  DFFARX1 next_result_adder_c_reg_6_ ( .D(result_adder_c[6]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[6]) );
  DFFARX1 next_result_adder_c_reg_5_ ( .D(result_adder_c[5]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[5]) );
  DFFARX1 next_result_adder_c_reg_4_ ( .D(result_adder_c[4]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[4]) );
  DFFARX1 next_result_adder_c_reg_3_ ( .D(result_adder_c[3]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[3]) );
  DFFARX1 next_result_adder_c_reg_2_ ( .D(result_adder_c[2]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[2]) );
  DFFARX1 next_result_adder_c_reg_1_ ( .D(result_adder_c[1]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[1]) );
  DFFARX1 next_result_adder_c_reg_0_ ( .D(result_adder_c[0]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_adder_c[0]) );
  DFFARX1 next_result_mult_d_reg_31_ ( .D(result_mult_d[31]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_d[31]) );
  DFFARX1 next_result_mult_d_reg_30_ ( .D(result_mult_d[30]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_d[30]) );
  DFFARX1 next_result_mult_d_reg_29_ ( .D(result_mult_d[29]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_d[29]) );
  DFFARX1 next_result_mult_d_reg_28_ ( .D(result_mult_d[28]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_d[28]) );
  DFFARX1 next_result_mult_d_reg_27_ ( .D(result_mult_d[27]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_d[27]) );
  DFFARX1 next_result_mult_d_reg_26_ ( .D(result_mult_d[26]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_d[26]) );
  DFFARX1 next_result_mult_d_reg_25_ ( .D(result_mult_d[25]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_d[25]) );
  DFFARX1 next_result_mult_d_reg_24_ ( .D(result_mult_d[24]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_d[24]) );
  DFFARX1 next_result_mult_d_reg_23_ ( .D(result_mult_d[23]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_d[23]) );
  DFFARX1 next_result_mult_d_reg_22_ ( .D(result_mult_d[22]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_d[22]) );
  DFFARX1 next_result_mult_d_reg_21_ ( .D(result_mult_d[21]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_d[21]) );
  DFFARX1 next_result_mult_d_reg_20_ ( .D(result_mult_d[20]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_d[20]) );
  DFFARX1 next_result_mult_d_reg_19_ ( .D(result_mult_d[19]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_d[19]) );
  DFFARX1 next_result_mult_d_reg_18_ ( .D(result_mult_d[18]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_d[18]) );
  DFFARX1 next_result_mult_d_reg_17_ ( .D(result_mult_d[17]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_d[17]) );
  DFFARX1 next_result_mult_d_reg_16_ ( .D(result_mult_d[16]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_d[16]) );
  DFFARX1 next_result_mult_d_reg_15_ ( .D(result_mult_d[15]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_d[15]) );
  DFFARX1 next_result_mult_d_reg_14_ ( .D(result_mult_d[14]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_d[14]) );
  DFFARX1 next_result_mult_d_reg_13_ ( .D(result_mult_d[13]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_d[13]) );
  DFFARX1 next_result_mult_d_reg_12_ ( .D(result_mult_d[12]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_d[12]) );
  DFFARX1 next_result_mult_d_reg_11_ ( .D(result_mult_d[11]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_d[11]) );
  DFFARX1 next_result_mult_d_reg_10_ ( .D(result_mult_d[10]), .CLK(clk), 
        .RSTB(rst_n), .Q(next_result_mult_d[10]) );
  DFFARX1 next_result_mult_d_reg_9_ ( .D(result_mult_d[9]), .CLK(clk), .RSTB(
        rst_n), .Q(next_result_mult_d[9]) );
  DFFARX1 next_result_mult_d_reg_8_ ( .D(result_mult_d[8]), .CLK(clk), .RSTB(
        rst_n), .Q(next_result_mult_d[8]) );
  DFFARX1 next_result_mult_d_reg_7_ ( .D(result_mult_d[7]), .CLK(clk), .RSTB(
        rst_n), .Q(next_result_mult_d[7]) );
  DFFARX1 next_result_mult_d_reg_6_ ( .D(result_mult_d[6]), .CLK(clk), .RSTB(
        rst_n), .Q(next_result_mult_d[6]) );
  DFFARX1 next_result_mult_d_reg_5_ ( .D(result_mult_d[5]), .CLK(clk), .RSTB(
        rst_n), .Q(next_result_mult_d[5]) );
  DFFARX1 next_result_mult_d_reg_4_ ( .D(result_mult_d[4]), .CLK(clk), .RSTB(
        rst_n), .Q(next_result_mult_d[4]) );
  DFFARX1 next_result_mult_d_reg_3_ ( .D(result_mult_d[3]), .CLK(clk), .RSTB(
        rst_n), .Q(next_result_mult_d[3]) );
  DFFARX1 next_result_mult_d_reg_2_ ( .D(result_mult_d[2]), .CLK(clk), .RSTB(
        rst_n), .Q(next_result_mult_d[2]) );
  DFFARX1 next_result_mult_d_reg_1_ ( .D(result_mult_d[1]), .CLK(clk), .RSTB(
        rst_n), .Q(next_result_mult_d[1]) );
  DFFARX1 next_result_mult_d_reg_0_ ( .D(result_mult_d[0]), .CLK(clk), .RSTB(
        rst_n), .Q(next_result_mult_d[0]) );
  DFFARX1 tansigmoid_output_reg_31_ ( .D(result_adder_d[31]), .CLK(clk), 
        .RSTB(rst_n), .Q(tansigmoid_output[31]) );
  DFFARX1 tansigmoid_output_reg_30_ ( .D(result_adder_d[30]), .CLK(clk), 
        .RSTB(rst_n), .Q(tansigmoid_output[30]) );
  DFFARX1 tansigmoid_output_reg_29_ ( .D(result_adder_d[29]), .CLK(clk), 
        .RSTB(rst_n), .Q(tansigmoid_output[29]) );
  DFFARX1 tansigmoid_output_reg_28_ ( .D(result_adder_d[28]), .CLK(clk), 
        .RSTB(rst_n), .Q(tansigmoid_output[28]) );
  DFFARX1 tansigmoid_output_reg_27_ ( .D(result_adder_d[27]), .CLK(clk), 
        .RSTB(rst_n), .Q(tansigmoid_output[27]) );
  DFFARX1 tansigmoid_output_reg_26_ ( .D(result_adder_d[26]), .CLK(clk), 
        .RSTB(rst_n), .Q(tansigmoid_output[26]) );
  DFFARX1 tansigmoid_output_reg_25_ ( .D(result_adder_d[25]), .CLK(clk), 
        .RSTB(rst_n), .Q(tansigmoid_output[25]) );
  DFFARX1 tansigmoid_output_reg_24_ ( .D(result_adder_d[24]), .CLK(clk), 
        .RSTB(rst_n), .Q(tansigmoid_output[24]) );
  DFFARX1 tansigmoid_output_reg_23_ ( .D(result_adder_d[23]), .CLK(clk), 
        .RSTB(rst_n), .Q(tansigmoid_output[23]) );
  DFFARX1 tansigmoid_output_reg_22_ ( .D(result_adder_d[22]), .CLK(clk), 
        .RSTB(rst_n), .Q(tansigmoid_output[22]) );
  DFFARX1 tansigmoid_output_reg_21_ ( .D(result_adder_d[21]), .CLK(clk), 
        .RSTB(rst_n), .Q(tansigmoid_output[21]) );
  DFFARX1 tansigmoid_output_reg_20_ ( .D(result_adder_d[20]), .CLK(clk), 
        .RSTB(rst_n), .Q(tansigmoid_output[20]) );
  DFFARX1 tansigmoid_output_reg_19_ ( .D(result_adder_d[19]), .CLK(clk), 
        .RSTB(rst_n), .Q(tansigmoid_output[19]) );
  DFFARX1 tansigmoid_output_reg_18_ ( .D(result_adder_d[18]), .CLK(clk), 
        .RSTB(rst_n), .Q(tansigmoid_output[18]) );
  DFFARX1 tansigmoid_output_reg_17_ ( .D(result_adder_d[17]), .CLK(clk), 
        .RSTB(rst_n), .Q(tansigmoid_output[17]) );
  DFFARX1 tansigmoid_output_reg_16_ ( .D(result_adder_d[16]), .CLK(clk), 
        .RSTB(rst_n), .Q(tansigmoid_output[16]) );
  DFFARX1 tansigmoid_output_reg_15_ ( .D(result_adder_d[15]), .CLK(clk), 
        .RSTB(rst_n), .Q(tansigmoid_output[15]) );
  DFFARX1 tansigmoid_output_reg_14_ ( .D(result_adder_d[14]), .CLK(clk), 
        .RSTB(rst_n), .Q(tansigmoid_output[14]) );
  DFFARX1 tansigmoid_output_reg_13_ ( .D(result_adder_d[13]), .CLK(clk), 
        .RSTB(rst_n), .Q(tansigmoid_output[13]) );
  DFFARX1 tansigmoid_output_reg_12_ ( .D(result_adder_d[12]), .CLK(clk), 
        .RSTB(rst_n), .Q(tansigmoid_output[12]) );
  DFFARX1 tansigmoid_output_reg_11_ ( .D(result_adder_d[11]), .CLK(clk), 
        .RSTB(rst_n), .Q(tansigmoid_output[11]) );
  DFFARX1 tansigmoid_output_reg_10_ ( .D(result_adder_d[10]), .CLK(clk), 
        .RSTB(rst_n), .Q(tansigmoid_output[10]) );
  DFFARX1 tansigmoid_output_reg_9_ ( .D(result_adder_d[9]), .CLK(clk), .RSTB(
        rst_n), .Q(tansigmoid_output[9]) );
  DFFARX1 tansigmoid_output_reg_8_ ( .D(result_adder_d[8]), .CLK(clk), .RSTB(
        rst_n), .Q(tansigmoid_output[8]) );
  DFFARX1 tansigmoid_output_reg_7_ ( .D(result_adder_d[7]), .CLK(clk), .RSTB(
        rst_n), .Q(tansigmoid_output[7]) );
  DFFARX1 tansigmoid_output_reg_6_ ( .D(result_adder_d[6]), .CLK(clk), .RSTB(
        rst_n), .Q(tansigmoid_output[6]) );
  DFFARX1 tansigmoid_output_reg_5_ ( .D(result_adder_d[5]), .CLK(clk), .RSTB(
        rst_n), .Q(tansigmoid_output[5]) );
  DFFARX1 tansigmoid_output_reg_4_ ( .D(result_adder_d[4]), .CLK(clk), .RSTB(
        rst_n), .Q(tansigmoid_output[4]) );
  DFFARX1 tansigmoid_output_reg_3_ ( .D(result_adder_d[3]), .CLK(clk), .RSTB(
        rst_n), .Q(tansigmoid_output[3]) );
  DFFARX1 tansigmoid_output_reg_2_ ( .D(result_adder_d[2]), .CLK(clk), .RSTB(
        rst_n), .Q(tansigmoid_output[2]) );
  DFFARX1 tansigmoid_output_reg_1_ ( .D(result_adder_d[1]), .CLK(clk), .RSTB(
        rst_n), .Q(tansigmoid_output[1]) );
  DFFARX1 tansigmoid_output_reg_0_ ( .D(result_adder_d[0]), .CLK(clk), .RSTB(
        rst_n), .Q(tansigmoid_output[0]) );
  NBUFFX8 U3 ( .INP(tansigmoid_input[10]), .Z(n4) );
  NBUFFX8 U4 ( .INP(tansigmoid_input[8]), .Z(n3) );
  NBUFFX8 U5 ( .INP(tansigmoid_input[4]), .Z(n2) );
  NBUFFX8 U6 ( .INP(tansigmoid_input[2]), .Z(n1) );
endmodule


module wr_int_mem_controller ( clk, rst_n, ena_wr_output_mem, is_odd_layer, 
        is_first_layer, change_layer, int_mem_addr_wr, output_mem_addr, 
        ena_wr_int_mem_BAR );
  output [19:0] int_mem_addr_wr;
  output [19:0] output_mem_addr;
  input clk, rst_n, ena_wr_output_mem, is_odd_layer, is_first_layer,
         change_layer, ena_wr_int_mem_BAR;
  wire   n3, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n1, n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123;
  wire   [9:0] addr_mem_back;
  wire   [9:0] addr_mem_front;

  DFFASX1 addr_mem_back_reg_9_ ( .D(n60), .CLK(clk), .SETB(rst_n), .Q(
        addr_mem_back[9]), .QN(n13) );
  DFFARX1 addr_mem_back_reg_8_ ( .D(n61), .CLK(clk), .RSTB(rst_n), .Q(
        addr_mem_back[8]), .QN(n7) );
  DFFARX1 addr_mem_back_reg_7_ ( .D(n62), .CLK(clk), .RSTB(rst_n), .Q(
        addr_mem_back[7]) );
  DFFARX1 addr_mem_back_reg_6_ ( .D(n63), .CLK(clk), .RSTB(rst_n), .Q(
        addr_mem_back[6]), .QN(n6) );
  DFFARX1 addr_mem_back_reg_5_ ( .D(n64), .CLK(clk), .RSTB(rst_n), .Q(
        addr_mem_back[5]) );
  DFFARX1 addr_mem_back_reg_4_ ( .D(n65), .CLK(clk), .RSTB(rst_n), .Q(
        addr_mem_back[4]), .QN(n5) );
  DFFARX1 addr_mem_back_reg_3_ ( .D(n66), .CLK(clk), .RSTB(rst_n), .Q(
        addr_mem_back[3]) );
  DFFARX1 addr_mem_back_reg_2_ ( .D(n67), .CLK(clk), .RSTB(rst_n), .Q(
        addr_mem_back[2]) );
  DFFARX1 addr_mem_back_reg_1_ ( .D(n68), .CLK(clk), .RSTB(rst_n), .Q(
        addr_mem_back[1]) );
  DFFARX1 addr_mem_back_reg_0_ ( .D(n69), .CLK(clk), .RSTB(rst_n), .Q(
        addr_mem_back[0]), .QN(n1) );
  DFFARX1 addr_mem_front_reg_9_ ( .D(n40), .CLK(clk), .RSTB(rst_n), .Q(
        addr_mem_front[9]) );
  DFFARX1 addr_mem_front_reg_8_ ( .D(n41), .CLK(clk), .RSTB(rst_n), .Q(
        addr_mem_front[8]), .QN(n10) );
  DFFARX1 addr_mem_front_reg_7_ ( .D(n42), .CLK(clk), .RSTB(rst_n), .Q(
        addr_mem_front[7]) );
  DFFARX1 addr_mem_front_reg_6_ ( .D(n43), .CLK(clk), .RSTB(rst_n), .Q(
        addr_mem_front[6]), .QN(n9) );
  DFFARX1 addr_mem_front_reg_5_ ( .D(n44), .CLK(clk), .RSTB(rst_n), .Q(
        addr_mem_front[5]) );
  DFFARX1 addr_mem_front_reg_4_ ( .D(n45), .CLK(clk), .RSTB(rst_n), .Q(
        addr_mem_front[4]), .QN(n8) );
  DFFARX1 addr_mem_front_reg_3_ ( .D(n46), .CLK(clk), .RSTB(rst_n), .Q(
        addr_mem_front[3]) );
  DFFARX1 addr_mem_front_reg_2_ ( .D(n47), .CLK(clk), .RSTB(rst_n), .Q(
        addr_mem_front[2]) );
  DFFARX1 addr_mem_front_reg_1_ ( .D(n48), .CLK(clk), .RSTB(rst_n), .Q(
        addr_mem_front[1]) );
  DFFARX1 addr_mem_front_reg_0_ ( .D(n49), .CLK(clk), .RSTB(rst_n), .Q(
        addr_mem_front[0]), .QN(n2) );
  DFFARX1 output_mem_addr_reg_9_ ( .D(n20), .CLK(clk), .RSTB(rst_n), .Q(
        output_mem_addr[9]), .QN(n4) );
  DFFARX1 output_mem_addr_reg_8_ ( .D(n21), .CLK(clk), .RSTB(rst_n), .Q(
        output_mem_addr[8]) );
  DFFARX1 output_mem_addr_reg_7_ ( .D(n22), .CLK(clk), .RSTB(rst_n), .Q(
        output_mem_addr[7]) );
  DFFARX1 output_mem_addr_reg_6_ ( .D(n23), .CLK(clk), .RSTB(rst_n), .Q(
        output_mem_addr[6]), .QN(n11) );
  DFFARX1 output_mem_addr_reg_5_ ( .D(n24), .CLK(clk), .RSTB(rst_n), .Q(
        output_mem_addr[5]) );
  DFFARX1 output_mem_addr_reg_4_ ( .D(n25), .CLK(clk), .RSTB(rst_n), .Q(
        output_mem_addr[4]), .QN(n12) );
  DFFARX1 output_mem_addr_reg_3_ ( .D(n26), .CLK(clk), .RSTB(rst_n), .Q(
        output_mem_addr[3]) );
  DFFARX1 output_mem_addr_reg_2_ ( .D(n27), .CLK(clk), .RSTB(rst_n), .Q(
        output_mem_addr[2]) );
  DFFARX1 output_mem_addr_reg_1_ ( .D(n28), .CLK(clk), .RSTB(rst_n), .Q(
        output_mem_addr[1]) );
  DFFARX1 output_mem_addr_reg_0_ ( .D(n29), .CLK(clk), .RSTB(rst_n), .Q(
        output_mem_addr[0]) );
  DFFASX1 ena_wr_int_mem_w1_reg ( .D(ena_wr_int_mem_BAR), .CLK(clk), .SETB(
        rst_n), .Q(n3) );
  NAND2X0 U3 ( .IN1(n120), .IN2(n117), .QN(n122) );
  NAND2X0 U4 ( .IN1(n117), .IN2(n95), .QN(n98) );
  NAND2X0 U5 ( .IN1(output_mem_addr[8]), .IN2(output_mem_addr[7]), .QN(n112)
         );
  NAND2X0 U6 ( .IN1(n120), .IN2(n2), .QN(n58) );
  NAND2X0 U7 ( .IN1(n94), .IN2(n58), .QN(n71) );
  NAND2X0 U8 ( .IN1(n92), .IN2(n93), .QN(n94) );
  NAND2X0 U9 ( .IN1(n120), .IN2(n1), .QN(n15) );
  NAND2X0 U10 ( .IN1(n94), .IN2(n15), .QN(n18) );
  NAND2X0 U11 ( .IN1(output_mem_addr[1]), .IN2(output_mem_addr[0]), .QN(n96)
         );
  NAND2X0 U12 ( .IN1(n121), .IN2(n4), .QN(n114) );
  NAND2X0 U13 ( .IN1(addr_mem_front[1]), .IN2(addr_mem_front[0]), .QN(n59) );
  NAND2X0 U14 ( .IN1(addr_mem_back[1]), .IN2(addr_mem_back[0]), .QN(n16) );
  NAND2X0 U15 ( .IN1(n56), .IN2(n92), .QN(n60) );
  NOR2X0 U16 ( .IN1(is_odd_layer), .IN2(is_first_layer), .QN(n14) );
  NAND2X0 U17 ( .IN1(n3), .IN2(n123), .QN(n93) );
  INVX0 U18 ( .INP(n118), .ZN(n120) );
  INVX0 U19 ( .INP(change_layer), .ZN(n92) );
  NAND3X0 U20 ( .IN1(n3), .IN2(n92), .IN3(n123), .QN(n118) );
  INVX0 U21 ( .INP(ena_wr_int_mem_BAR), .ZN(n123) );
  MUX21X1 U22 ( .IN1(addr_mem_front[0]), .IN2(addr_mem_back[0]), .S(n14), .Q(
        int_mem_addr_wr[0]) );
  MUX21X1 U23 ( .IN1(addr_mem_front[1]), .IN2(addr_mem_back[1]), .S(n14), .Q(
        int_mem_addr_wr[1]) );
  MUX21X1 U24 ( .IN1(addr_mem_front[2]), .IN2(addr_mem_back[2]), .S(n14), .Q(
        int_mem_addr_wr[2]) );
  MUX21X1 U25 ( .IN1(addr_mem_front[3]), .IN2(addr_mem_back[3]), .S(n14), .Q(
        int_mem_addr_wr[3]) );
  MUX21X1 U26 ( .IN1(addr_mem_front[4]), .IN2(addr_mem_back[4]), .S(n14), .Q(
        int_mem_addr_wr[4]) );
  MUX21X1 U27 ( .IN1(addr_mem_front[5]), .IN2(addr_mem_back[5]), .S(n14), .Q(
        int_mem_addr_wr[5]) );
  MUX21X1 U28 ( .IN1(addr_mem_front[6]), .IN2(addr_mem_back[6]), .S(n14), .Q(
        int_mem_addr_wr[6]) );
  MUX21X1 U29 ( .IN1(addr_mem_front[7]), .IN2(addr_mem_back[7]), .S(n14), .Q(
        int_mem_addr_wr[7]) );
  MUX21X1 U30 ( .IN1(addr_mem_front[8]), .IN2(addr_mem_back[8]), .S(n14), .Q(
        int_mem_addr_wr[8]) );
  MUX21X1 U31 ( .IN1(addr_mem_front[9]), .IN2(addr_mem_back[9]), .S(n14), .Q(
        int_mem_addr_wr[9]) );
  OAI21X1 U32 ( .IN1(n1), .IN2(n94), .IN3(n15), .QN(n69) );
  NOR2X0 U33 ( .IN1(addr_mem_back[1]), .IN2(n118), .QN(n19) );
  AO22X1 U34 ( .IN1(addr_mem_back[1]), .IN2(n18), .IN3(addr_mem_back[0]), 
        .IN4(n19), .Q(n68) );
  NOR3X0 U35 ( .IN1(addr_mem_back[2]), .IN2(n16), .IN3(n118), .QN(n17) );
  AO221X1 U36 ( .IN1(addr_mem_back[2]), .IN2(n19), .IN3(addr_mem_back[2]), 
        .IN4(n18), .IN5(n17), .Q(n67) );
  NAND3X0 U37 ( .IN1(addr_mem_back[1]), .IN2(addr_mem_back[0]), .IN3(
        addr_mem_back[2]), .QN(n30) );
  INVX0 U38 ( .INP(n30), .ZN(n34) );
  NOR2X0 U39 ( .IN1(addr_mem_back[3]), .IN2(n118), .QN(n33) );
  OA21X1 U40 ( .IN1(n93), .IN2(n30), .IN3(n92), .Q(n32) );
  AO22X1 U41 ( .IN1(n34), .IN2(n33), .IN3(addr_mem_back[3]), .IN4(n32), .Q(n66) );
  AND3X1 U42 ( .IN1(n120), .IN2(n34), .IN3(addr_mem_back[3]), .Q(n31) );
  AO222X1 U43 ( .IN1(addr_mem_back[4]), .IN2(n33), .IN3(addr_mem_back[4]), 
        .IN4(n32), .IN5(n31), .IN6(n5), .Q(n65) );
  NAND3X0 U44 ( .IN1(n34), .IN2(addr_mem_back[4]), .IN3(addr_mem_back[3]), 
        .QN(n35) );
  INVX0 U45 ( .INP(n35), .ZN(n39) );
  NOR2X0 U46 ( .IN1(addr_mem_back[5]), .IN2(n118), .QN(n38) );
  OA21X1 U47 ( .IN1(n93), .IN2(n35), .IN3(n92), .Q(n37) );
  AO22X1 U48 ( .IN1(n39), .IN2(n38), .IN3(addr_mem_back[5]), .IN4(n37), .Q(n64) );
  AND3X1 U49 ( .IN1(n120), .IN2(n39), .IN3(addr_mem_back[5]), .Q(n36) );
  AO222X1 U50 ( .IN1(addr_mem_back[6]), .IN2(n38), .IN3(addr_mem_back[6]), 
        .IN4(n37), .IN5(n36), .IN6(n6), .Q(n63) );
  NAND3X0 U51 ( .IN1(n39), .IN2(addr_mem_back[6]), .IN3(addr_mem_back[5]), 
        .QN(n50) );
  INVX0 U52 ( .INP(n50), .ZN(n54) );
  NOR2X0 U53 ( .IN1(addr_mem_back[7]), .IN2(n118), .QN(n53) );
  OA21X1 U54 ( .IN1(n93), .IN2(n50), .IN3(n92), .Q(n52) );
  AO22X1 U55 ( .IN1(n54), .IN2(n53), .IN3(addr_mem_back[7]), .IN4(n52), .Q(n62) );
  AND3X1 U56 ( .IN1(n120), .IN2(n54), .IN3(addr_mem_back[7]), .Q(n51) );
  AO222X1 U57 ( .IN1(addr_mem_back[8]), .IN2(n53), .IN3(addr_mem_back[8]), 
        .IN4(n52), .IN5(n51), .IN6(n7), .Q(n61) );
  NAND3X0 U58 ( .IN1(n54), .IN2(addr_mem_back[8]), .IN3(addr_mem_back[7]), 
        .QN(n57) );
  NOR2X0 U59 ( .IN1(n93), .IN2(n57), .QN(n55) );
  MUX21X1 U60 ( .IN1(n13), .IN2(addr_mem_back[9]), .S(n55), .Q(n56) );
  OAI21X1 U61 ( .IN1(n2), .IN2(n94), .IN3(n58), .QN(n49) );
  NOR2X0 U62 ( .IN1(addr_mem_front[1]), .IN2(n118), .QN(n72) );
  AO22X1 U63 ( .IN1(addr_mem_front[1]), .IN2(n71), .IN3(addr_mem_front[0]), 
        .IN4(n72), .Q(n48) );
  NOR3X0 U64 ( .IN1(addr_mem_front[2]), .IN2(n59), .IN3(n118), .QN(n70) );
  AO221X1 U65 ( .IN1(addr_mem_front[2]), .IN2(n72), .IN3(addr_mem_front[2]), 
        .IN4(n71), .IN5(n70), .Q(n47) );
  NAND3X0 U66 ( .IN1(addr_mem_front[1]), .IN2(addr_mem_front[0]), .IN3(
        addr_mem_front[2]), .QN(n73) );
  INVX0 U67 ( .INP(n73), .ZN(n77) );
  NOR2X0 U68 ( .IN1(addr_mem_front[3]), .IN2(n118), .QN(n76) );
  OA21X1 U69 ( .IN1(n93), .IN2(n73), .IN3(n92), .Q(n75) );
  AO22X1 U70 ( .IN1(n77), .IN2(n76), .IN3(addr_mem_front[3]), .IN4(n75), .Q(
        n46) );
  AND3X1 U71 ( .IN1(n120), .IN2(n77), .IN3(addr_mem_front[3]), .Q(n74) );
  AO222X1 U72 ( .IN1(addr_mem_front[4]), .IN2(n76), .IN3(addr_mem_front[4]), 
        .IN4(n75), .IN5(n74), .IN6(n8), .Q(n45) );
  NAND3X0 U73 ( .IN1(n77), .IN2(addr_mem_front[4]), .IN3(addr_mem_front[3]), 
        .QN(n78) );
  INVX0 U74 ( .INP(n78), .ZN(n82) );
  NOR2X0 U75 ( .IN1(addr_mem_front[5]), .IN2(n118), .QN(n81) );
  OA21X1 U76 ( .IN1(n93), .IN2(n78), .IN3(n92), .Q(n80) );
  AO22X1 U77 ( .IN1(n82), .IN2(n81), .IN3(addr_mem_front[5]), .IN4(n80), .Q(
        n44) );
  AND3X1 U78 ( .IN1(n120), .IN2(n82), .IN3(addr_mem_front[5]), .Q(n79) );
  AO222X1 U79 ( .IN1(addr_mem_front[6]), .IN2(n81), .IN3(addr_mem_front[6]), 
        .IN4(n80), .IN5(n79), .IN6(n9), .Q(n43) );
  NAND3X0 U80 ( .IN1(n82), .IN2(addr_mem_front[6]), .IN3(addr_mem_front[5]), 
        .QN(n83) );
  INVX0 U81 ( .INP(n83), .ZN(n87) );
  NOR2X0 U82 ( .IN1(addr_mem_front[7]), .IN2(n118), .QN(n86) );
  OA21X1 U83 ( .IN1(n93), .IN2(n83), .IN3(n92), .Q(n85) );
  AO22X1 U84 ( .IN1(n87), .IN2(n86), .IN3(addr_mem_front[7]), .IN4(n85), .Q(
        n42) );
  AND3X1 U85 ( .IN1(n120), .IN2(n87), .IN3(addr_mem_front[7]), .Q(n84) );
  AO222X1 U86 ( .IN1(addr_mem_front[8]), .IN2(n86), .IN3(addr_mem_front[8]), 
        .IN4(n85), .IN5(n84), .IN6(n10), .Q(n41) );
  NAND3X0 U87 ( .IN1(n87), .IN2(addr_mem_front[8]), .IN3(addr_mem_front[7]), 
        .QN(n88) );
  INVX0 U88 ( .INP(n88), .ZN(n91) );
  NOR2X0 U89 ( .IN1(addr_mem_front[9]), .IN2(n118), .QN(n90) );
  OA21X1 U90 ( .IN1(n93), .IN2(n88), .IN3(n92), .Q(n89) );
  AO22X1 U91 ( .IN1(n91), .IN2(n90), .IN3(addr_mem_front[9]), .IN4(n89), .Q(
        n40) );
  OA21X1 U92 ( .IN1(change_layer), .IN2(ena_wr_output_mem), .IN3(n94), .Q(n117) );
  INVX0 U93 ( .INP(n122), .ZN(n121) );
  INVX0 U94 ( .INP(n117), .ZN(n119) );
  MUX21X1 U95 ( .IN1(n121), .IN2(n119), .S(output_mem_addr[0]), .Q(n29) );
  OR2X1 U96 ( .IN1(n122), .IN2(output_mem_addr[0]), .Q(n95) );
  NOR2X0 U97 ( .IN1(output_mem_addr[1]), .IN2(n122), .QN(n99) );
  AO22X1 U98 ( .IN1(output_mem_addr[1]), .IN2(n98), .IN3(output_mem_addr[0]), 
        .IN4(n99), .Q(n28) );
  NOR3X0 U99 ( .IN1(output_mem_addr[2]), .IN2(n96), .IN3(n122), .QN(n97) );
  AO221X1 U100 ( .IN1(output_mem_addr[2]), .IN2(n99), .IN3(output_mem_addr[2]), 
        .IN4(n98), .IN5(n97), .Q(n27) );
  AND3X1 U101 ( .IN1(output_mem_addr[1]), .IN2(output_mem_addr[0]), .IN3(
        output_mem_addr[2]), .Q(n103) );
  NOR2X0 U102 ( .IN1(output_mem_addr[3]), .IN2(n122), .QN(n102) );
  OAI21X1 U103 ( .IN1(n103), .IN2(n118), .IN3(n117), .QN(n101) );
  AO22X1 U104 ( .IN1(n103), .IN2(n102), .IN3(output_mem_addr[3]), .IN4(n101), 
        .Q(n26) );
  AND3X1 U105 ( .IN1(n121), .IN2(n103), .IN3(output_mem_addr[3]), .Q(n100) );
  AO222X1 U106 ( .IN1(output_mem_addr[4]), .IN2(n102), .IN3(output_mem_addr[4]), .IN4(n101), .IN5(n100), .IN6(n12), .Q(n25) );
  AND3X1 U107 ( .IN1(n103), .IN2(output_mem_addr[4]), .IN3(output_mem_addr[3]), 
        .Q(n107) );
  NOR2X0 U108 ( .IN1(output_mem_addr[5]), .IN2(n122), .QN(n106) );
  OAI21X1 U109 ( .IN1(n107), .IN2(n118), .IN3(n117), .QN(n105) );
  AO22X1 U110 ( .IN1(n107), .IN2(n106), .IN3(output_mem_addr[5]), .IN4(n105), 
        .Q(n24) );
  AND3X1 U111 ( .IN1(n121), .IN2(n107), .IN3(output_mem_addr[5]), .Q(n104) );
  AO222X1 U112 ( .IN1(output_mem_addr[6]), .IN2(n106), .IN3(output_mem_addr[6]), .IN4(n105), .IN5(n104), .IN6(n11), .Q(n23) );
  NAND3X0 U113 ( .IN1(n107), .IN2(output_mem_addr[6]), .IN3(output_mem_addr[5]), .QN(n111) );
  NOR2X0 U114 ( .IN1(n122), .IN2(n111), .QN(n108) );
  AO21X1 U115 ( .IN1(n120), .IN2(n111), .IN3(n119), .Q(n109) );
  MUX21X1 U116 ( .IN1(n108), .IN2(n109), .S(output_mem_addr[7]), .Q(n22) );
  AO21X1 U117 ( .IN1(output_mem_addr[7]), .IN2(n108), .IN3(output_mem_addr[8]), 
        .Q(n110) );
  AO221X1 U118 ( .IN1(n110), .IN2(n112), .IN3(n110), .IN4(n109), .IN5(
        change_layer), .Q(n21) );
  NOR2X0 U119 ( .IN1(n112), .IN2(n111), .QN(n116) );
  OA21X1 U120 ( .IN1(n116), .IN2(n118), .IN3(n117), .Q(n115) );
  INVX0 U121 ( .INP(n116), .ZN(n113) );
  OAI22X1 U122 ( .IN1(n115), .IN2(n4), .IN3(n113), .IN4(n114), .QN(n20) );
endmodule


module network_control ( clk, rst_n, ena_neural, mac_time, num_of_layer, 
        num_of_node_for_each_layer, ena_rd_user_para, ena_mac, ena_mac_wait, 
        ena_act_func, input_or_int_mem_sel, is_first_layer, is_odd_layer, 
        refresh_mac, change_layer, ena_wr_output_mem, end_neural, 
        ena_wr_int_mem_BAR );
  input [11:0] mac_time;
  input [3:0] num_of_layer;
  input [7:0] num_of_node_for_each_layer;
  input clk, rst_n, ena_neural;
  output ena_rd_user_para, ena_mac, ena_mac_wait, ena_act_func,
         input_or_int_mem_sel, is_first_layer, is_odd_layer, refresh_mac,
         change_layer, ena_wr_output_mem, end_neural, ena_wr_int_mem_BAR;
  wire   N146, N147, N148, N149, N150, N151, N152, N153, N172, N173, N174,
         N175, N176, N177, N178, N179, N208, N209, N210, N211, N212, N213,
         N214, N215, N216, N217, N218, N219, N239, N240, N241, N242, N243,
         N244, N245, N246, N265, N266, N267, N268, N269, N270, N271, N272,
         N291, N292, N293, N294, N295, N296, N297, N298, ena_setup_w4, N320,
         is_last_layer, N334, n1, n2, n3, n4, n13, n14, n21, n29, n42, n43,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n5, n6, n7, n8, n9, n10, n11, n12, n15,
         n16, n17, n18, n19, n20, n22, n23, n24, n25, n26, n27, n28, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n44, n45, n46, n47,
         n48, n50, n51, n52, n53, n54, n55, n56, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278;
  wire   [2:1] state;
  wire   [7:0] counter_rd_user_para;
  wire   [7:0] counter_setup;
  wire   [11:0] counter_mac;
  wire   [7:0] counter_mac_wait;
  wire   [7:0] counter_act_func;
  wire   [7:0] counter_wr_int_mem;
  wire   [7:0] node_counter;
  wire   [3:0] layer_counter;

  DFFARX1 is_last_layer_reg ( .D(N334), .CLK(clk), .RSTB(rst_n), .Q(
        is_last_layer), .QN(n51) );
  DFFARX1 state_reg_1_ ( .D(n123), .CLK(clk), .RSTB(rst_n), .Q(state[1]), .QN(
        n9) );
  DFFARX1 state_reg_0_ ( .D(n122), .CLK(clk), .RSTB(rst_n), .Q(n5), .QN(n13)
         );
  DFFARX1 counter_mac_wait_reg_7_ ( .D(N246), .CLK(clk), .RSTB(rst_n), .Q(
        counter_mac_wait[7]), .QN(n53) );
  DFFARX1 counter_mac_wait_reg_6_ ( .D(N245), .CLK(clk), .RSTB(rst_n), .Q(
        counter_mac_wait[6]), .QN(n33) );
  DFFARX1 counter_mac_wait_reg_5_ ( .D(N244), .CLK(clk), .RSTB(rst_n), .Q(
        counter_mac_wait[5]) );
  DFFARX1 counter_mac_wait_reg_4_ ( .D(N243), .CLK(clk), .RSTB(rst_n), .Q(
        counter_mac_wait[4]), .QN(n30) );
  DFFARX1 counter_mac_wait_reg_3_ ( .D(N242), .CLK(clk), .RSTB(rst_n), .Q(
        counter_mac_wait[3]) );
  DFFARX1 counter_mac_wait_reg_2_ ( .D(N241), .CLK(clk), .RSTB(rst_n), .Q(
        counter_mac_wait[2]) );
  DFFARX1 counter_mac_wait_reg_1_ ( .D(N240), .CLK(clk), .RSTB(rst_n), .Q(
        counter_mac_wait[1]) );
  DFFARX1 counter_mac_wait_reg_0_ ( .D(N239), .CLK(clk), .RSTB(rst_n), .Q(
        counter_mac_wait[0]) );
  DFFARX1 state_reg_2_ ( .D(n124), .CLK(clk), .RSTB(rst_n), .Q(state[2]) );
  DFFARX1 counter_rd_user_para_reg_7_ ( .D(N153), .CLK(clk), .RSTB(rst_n), .Q(
        counter_rd_user_para[7]), .QN(n54) );
  DFFARX1 counter_rd_user_para_reg_6_ ( .D(N152), .CLK(clk), .RSTB(rst_n), .Q(
        counter_rd_user_para[6]), .QN(n36) );
  DFFARX1 counter_rd_user_para_reg_5_ ( .D(N151), .CLK(clk), .RSTB(rst_n), .Q(
        counter_rd_user_para[5]) );
  DFFARX1 counter_rd_user_para_reg_4_ ( .D(N150), .CLK(clk), .RSTB(rst_n), .Q(
        counter_rd_user_para[4]), .QN(n26) );
  DFFARX1 counter_rd_user_para_reg_3_ ( .D(N149), .CLK(clk), .RSTB(rst_n), .Q(
        counter_rd_user_para[3]) );
  DFFARX1 counter_rd_user_para_reg_2_ ( .D(N148), .CLK(clk), .RSTB(rst_n), .Q(
        counter_rd_user_para[2]), .QN(n23) );
  DFFARX1 counter_rd_user_para_reg_1_ ( .D(N147), .CLK(clk), .RSTB(rst_n), .Q(
        counter_rd_user_para[1]) );
  DFFARX1 counter_rd_user_para_reg_0_ ( .D(N146), .CLK(clk), .RSTB(rst_n), .Q(
        counter_rd_user_para[0]) );
  DFFARX1 counter_setup_reg_7_ ( .D(N179), .CLK(clk), .RSTB(rst_n), .Q(
        counter_setup[7]), .QN(n55) );
  DFFARX1 counter_setup_reg_6_ ( .D(N178), .CLK(clk), .RSTB(rst_n), .Q(
        counter_setup[6]), .QN(n35) );
  DFFARX1 counter_setup_reg_5_ ( .D(N177), .CLK(clk), .RSTB(rst_n), .Q(
        counter_setup[5]) );
  DFFARX1 counter_setup_reg_4_ ( .D(N176), .CLK(clk), .RSTB(rst_n), .Q(
        counter_setup[4]) );
  DFFARX1 counter_setup_reg_3_ ( .D(N175), .CLK(clk), .RSTB(rst_n), .Q(
        counter_setup[3]), .QN(n25) );
  DFFARX1 counter_setup_reg_2_ ( .D(N174), .CLK(clk), .RSTB(rst_n), .Q(
        counter_setup[2]) );
  DFFARX1 counter_setup_reg_1_ ( .D(N173), .CLK(clk), .RSTB(rst_n), .Q(
        counter_setup[1]) );
  DFFARX1 counter_setup_reg_0_ ( .D(N172), .CLK(clk), .RSTB(rst_n), .Q(
        counter_setup[0]) );
  DFFASX1 ena_setup_w1_reg ( .D(n43), .CLK(clk), .SETB(rst_n), .Q(n4) );
  DFFASX1 ena_setup_w2_reg ( .D(n4), .CLK(clk), .SETB(rst_n), .Q(n3) );
  DFFASX1 ena_setup_w3_reg ( .D(n3), .CLK(clk), .SETB(rst_n), .Q(n2) );
  DFFASX1 ena_setup_w4_reg ( .D(n2), .CLK(clk), .SETB(rst_n), .Q(n1), .QN(
        ena_setup_w4) );
  DFFASX1 ena_setup_w5_reg ( .D(n1), .CLK(clk), .SETB(rst_n), .Q(n14) );
  DFFARX1 node_counter_reg_7_ ( .D(n114), .CLK(clk), .RSTB(rst_n), .Q(
        node_counter[7]), .QN(n31) );
  DFFARX1 node_counter_reg_6_ ( .D(n115), .CLK(clk), .RSTB(rst_n), .Q(
        node_counter[6]), .QN(n8) );
  DFFARX1 node_counter_reg_5_ ( .D(n116), .CLK(clk), .RSTB(rst_n), .Q(
        node_counter[5]), .QN(n38) );
  DFFARX1 node_counter_reg_4_ ( .D(n117), .CLK(clk), .RSTB(rst_n), .Q(
        node_counter[4]), .QN(n20) );
  DFFARX1 node_counter_reg_3_ ( .D(n118), .CLK(clk), .RSTB(rst_n), .Q(
        node_counter[3]), .QN(n41) );
  DFFARX1 node_counter_reg_2_ ( .D(n119), .CLK(clk), .RSTB(rst_n), .Q(
        node_counter[2]), .QN(n40) );
  DFFARX1 node_counter_reg_1_ ( .D(n120), .CLK(clk), .RSTB(rst_n), .Q(
        node_counter[1]), .QN(n17) );
  DFFARX1 node_counter_reg_0_ ( .D(n121), .CLK(clk), .RSTB(rst_n), .Q(
        node_counter[0]), .QN(n6) );
  DFFARX1 change_layer_reg ( .D(N320), .CLK(clk), .RSTB(rst_n), .Q(
        change_layer), .QN(n18) );
  DFFARX1 layer_counter_reg_0_ ( .D(n113), .CLK(clk), .RSTB(rst_n), .Q(
        layer_counter[0]), .QN(n44) );
  DFFASX1 layer_counter_reg_1_ ( .D(n29), .CLK(clk), .SETB(rst_n), .Q(n19), 
        .QN(layer_counter[1]) );
  DFFARX1 layer_counter_reg_2_ ( .D(n112), .CLK(clk), .RSTB(rst_n), .Q(
        layer_counter[2]), .QN(n7) );
  DFFARX1 layer_counter_reg_3_ ( .D(n111), .CLK(clk), .RSTB(rst_n), .Q(
        layer_counter[3]), .QN(n24) );
  DFFARX1 counter_mac_reg_11_ ( .D(N219), .CLK(clk), .RSTB(rst_n), .Q(
        counter_mac[11]), .QN(n32) );
  DFFARX1 counter_mac_reg_10_ ( .D(N218), .CLK(clk), .RSTB(rst_n), .Q(
        counter_mac[10]), .QN(n16) );
  DFFARX1 counter_mac_reg_9_ ( .D(N217), .CLK(clk), .RSTB(rst_n), .Q(
        counter_mac[9]), .QN(n45) );
  DFFARX1 counter_mac_reg_8_ ( .D(N216), .CLK(clk), .RSTB(rst_n), .Q(
        counter_mac[8]), .QN(n15) );
  DFFARX1 counter_mac_reg_7_ ( .D(N215), .CLK(clk), .RSTB(rst_n), .Q(
        counter_mac[7]), .QN(n47) );
  DFFARX1 counter_mac_reg_6_ ( .D(N214), .CLK(clk), .RSTB(rst_n), .Q(
        counter_mac[6]), .QN(n12) );
  DFFARX1 counter_mac_reg_5_ ( .D(N213), .CLK(clk), .RSTB(rst_n), .Q(
        counter_mac[5]), .QN(n46) );
  DFFARX1 counter_mac_reg_4_ ( .D(N212), .CLK(clk), .RSTB(rst_n), .Q(
        counter_mac[4]), .QN(n11) );
  DFFARX1 counter_mac_reg_3_ ( .D(N211), .CLK(clk), .RSTB(rst_n), .Q(
        counter_mac[3]), .QN(n48) );
  DFFARX1 counter_mac_reg_2_ ( .D(N210), .CLK(clk), .RSTB(rst_n), .Q(
        counter_mac[2]), .QN(n10) );
  DFFARX1 counter_mac_reg_1_ ( .D(N209), .CLK(clk), .RSTB(rst_n), .Q(
        counter_mac[1]), .QN(n50) );
  DFFARX1 counter_mac_reg_0_ ( .D(N208), .CLK(clk), .RSTB(rst_n), .Q(
        counter_mac[0]), .QN(n22) );
  DFFARX1 counter_wr_int_mem_reg_7_ ( .D(N298), .CLK(clk), .RSTB(rst_n), .Q(
        counter_wr_int_mem[7]), .QN(n56) );
  DFFARX1 counter_wr_int_mem_reg_6_ ( .D(N297), .CLK(clk), .RSTB(rst_n), .Q(
        counter_wr_int_mem[6]), .QN(n34) );
  DFFARX1 counter_wr_int_mem_reg_5_ ( .D(N296), .CLK(clk), .RSTB(rst_n), .Q(
        counter_wr_int_mem[5]) );
  DFFARX1 counter_wr_int_mem_reg_4_ ( .D(N295), .CLK(clk), .RSTB(rst_n), .Q(
        counter_wr_int_mem[4]), .QN(n27) );
  DFFARX1 counter_wr_int_mem_reg_3_ ( .D(N294), .CLK(clk), .RSTB(rst_n), .Q(
        counter_wr_int_mem[3]) );
  DFFARX1 counter_wr_int_mem_reg_2_ ( .D(N293), .CLK(clk), .RSTB(rst_n), .Q(
        counter_wr_int_mem[2]) );
  DFFARX1 counter_wr_int_mem_reg_1_ ( .D(N292), .CLK(clk), .RSTB(rst_n), .Q(
        counter_wr_int_mem[1]), .QN(n39) );
  DFFARX1 counter_wr_int_mem_reg_0_ ( .D(N291), .CLK(clk), .RSTB(rst_n), .Q(
        counter_wr_int_mem[0]) );
  DFFARX1 counter_act_func_reg_7_ ( .D(N272), .CLK(clk), .RSTB(rst_n), .Q(
        counter_act_func[7]), .QN(n52) );
  DFFARX1 counter_act_func_reg_6_ ( .D(N271), .CLK(clk), .RSTB(rst_n), .Q(
        counter_act_func[6]), .QN(n37) );
  DFFARX1 counter_act_func_reg_5_ ( .D(N270), .CLK(clk), .RSTB(rst_n), .Q(
        counter_act_func[5]) );
  DFFARX1 counter_act_func_reg_4_ ( .D(N269), .CLK(clk), .RSTB(rst_n), .Q(
        counter_act_func[4]), .QN(n28) );
  DFFARX1 counter_act_func_reg_3_ ( .D(N268), .CLK(clk), .RSTB(rst_n), .Q(
        counter_act_func[3]) );
  DFFARX1 counter_act_func_reg_2_ ( .D(N267), .CLK(clk), .RSTB(rst_n), .Q(
        counter_act_func[2]) );
  DFFARX1 counter_act_func_reg_1_ ( .D(N266), .CLK(clk), .RSTB(rst_n), .Q(
        counter_act_func[1]) );
  DFFARX1 counter_act_func_reg_0_ ( .D(N265), .CLK(clk), .RSTB(rst_n), .Q(
        counter_act_func[0]) );
  DFFARX1 is_first_layer_reg ( .D(n110), .CLK(clk), .RSTB(rst_n), .Q(
        is_first_layer) );
  DFFARX1 is_odd_layer_reg ( .D(n109), .CLK(clk), .RSTB(rst_n), .Q(
        is_odd_layer), .QN(n21) );
  DFFASX1 end_neural_reg ( .D(n42), .CLK(clk), .SETB(rst_n), .QN(end_neural)
         );
  NAND2X0 U3 ( .IN1(counter_wr_int_mem[0]), .IN2(n39), .QN(n202) );
  NAND3X0 U4 ( .IN1(state[2]), .IN2(n9), .IN3(n5), .QN(n176) );
  NAND2X0 U5 ( .IN1(ena_act_func), .IN2(n231), .QN(n191) );
  NAND2X0 U6 ( .IN1(counter_act_func[3]), .IN2(n192), .QN(n194) );
  NAND2X0 U7 ( .IN1(counter_act_func[5]), .IN2(n195), .QN(n196) );
  NAND2X0 U8 ( .IN1(counter_wr_int_mem[3]), .IN2(n206), .QN(n208) );
  NAND2X0 U9 ( .IN1(counter_wr_int_mem[5]), .IN2(n209), .QN(n210) );
  NAND2X0 U10 ( .IN1(counter_mac[0]), .IN2(counter_mac[1]), .QN(n155) );
  NAND2X0 U11 ( .IN1(counter_mac[3]), .IN2(n156), .QN(n158) );
  NAND2X0 U12 ( .IN1(counter_mac[5]), .IN2(n159), .QN(n161) );
  NAND2X0 U13 ( .IN1(counter_mac[7]), .IN2(n162), .QN(n164) );
  NAND2X0 U14 ( .IN1(counter_mac[9]), .IN2(n165), .QN(n166) );
  NAND2X0 U15 ( .IN1(n256), .IN2(n252), .QN(n254) );
  NAND2X0 U16 ( .IN1(n269), .IN2(n6), .QN(n252) );
  NAND2X0 U17 ( .IN1(counter_setup[1]), .IN2(counter_setup[0]), .QN(n125) );
  NAND2X0 U18 ( .IN1(counter_setup[5]), .IN2(n132), .QN(n133) );
  NAND2X0 U19 ( .IN1(counter_rd_user_para[1]), .IN2(counter_rd_user_para[0]), 
        .QN(n98) );
  NAND2X0 U20 ( .IN1(counter_rd_user_para[5]), .IN2(n102), .QN(n103) );
  NAND2X0 U21 ( .IN1(counter_mac_wait[1]), .IN2(counter_mac_wait[0]), .QN(n172) );
  NAND2X0 U22 ( .IN1(n177), .IN2(counter_mac_wait[3]), .QN(n179) );
  NAND2X0 U23 ( .IN1(counter_mac_wait[5]), .IN2(n180), .QN(n181) );
  NAND2X0 U24 ( .IN1(n18), .IN2(n247), .QN(n240) );
  NAND2X0 U25 ( .IN1(ena_mac), .IN2(n229), .QN(n233) );
  NAND2X0 U26 ( .IN1(n194), .IN2(n198), .QN(n65) );
  NAND2X0 U27 ( .IN1(n196), .IN2(n198), .QN(n63) );
  NAND2X0 U28 ( .IN1(n37), .IN2(n196), .QN(n197) );
  NAND2X0 U29 ( .IN1(n208), .IN2(n212), .QN(n61) );
  NAND2X0 U30 ( .IN1(n210), .IN2(n212), .QN(n59) );
  NAND2X0 U31 ( .IN1(n34), .IN2(n210), .QN(n211) );
  NAND2X0 U32 ( .IN1(n155), .IN2(n168), .QN(n81) );
  NAND2X0 U33 ( .IN1(n158), .IN2(n168), .QN(n79) );
  NAND2X0 U34 ( .IN1(n161), .IN2(n168), .QN(n77) );
  NAND2X0 U35 ( .IN1(n164), .IN2(n168), .QN(n75) );
  NAND2X0 U36 ( .IN1(n166), .IN2(n168), .QN(n73) );
  NAND2X0 U37 ( .IN1(n16), .IN2(n166), .QN(n167) );
  NAND2X0 U38 ( .IN1(n272), .IN2(n19), .QN(n273) );
  NAND2X0 U39 ( .IN1(n125), .IN2(n135), .QN(n87) );
  NAND2X0 U40 ( .IN1(n127), .IN2(n135), .QN(n85) );
  NAND2X0 U41 ( .IN1(n133), .IN2(n135), .QN(n83) );
  NAND2X0 U42 ( .IN1(n35), .IN2(n133), .QN(n134) );
  NAND2X0 U43 ( .IN1(n98), .IN2(n105), .QN(n93) );
  NAND2X0 U44 ( .IN1(n101), .IN2(n105), .QN(n91) );
  NAND2X0 U45 ( .IN1(n103), .IN2(n105), .QN(n89) );
  NAND2X0 U46 ( .IN1(n36), .IN2(n103), .QN(n104) );
  NAND2X0 U47 ( .IN1(n172), .IN2(n183), .QN(n71) );
  NAND2X0 U48 ( .IN1(n179), .IN2(ena_mac_wait), .QN(n69) );
  NAND2X0 U49 ( .IN1(n181), .IN2(n183), .QN(n67) );
  NAND2X0 U50 ( .IN1(n33), .IN2(n181), .QN(n182) );
  NAND2X0 U51 ( .IN1(n245), .IN2(ena_mac_wait), .QN(n250) );
  NAND2X0 U52 ( .IN1(n42), .IN2(n240), .QN(n241) );
  NAND3X0 U53 ( .IN1(state[1]), .IN2(state[2]), .IN3(n5), .QN(
        ena_wr_int_mem_BAR) );
  NAND2X0 U54 ( .IN1(ena_setup_w4), .IN2(n14), .QN(n262) );
  NAND2X0 U55 ( .IN1(refresh_mac), .IN2(n5), .QN(n43) );
  NAND2X0 U56 ( .IN1(change_layer), .IN2(is_last_layer), .QN(n42) );
  NOR2X0 U57 ( .IN1(n229), .IN2(n153), .QN(n168) );
  NOR2X0 U58 ( .IN1(state[2]), .IN2(n9), .QN(refresh_mac) );
  NOR2X0 U59 ( .IN1(n9), .IN2(n186), .QN(ena_act_func) );
  NOR2X0 U60 ( .IN1(state[1]), .IN2(n186), .QN(ena_mac) );
  NAND2X0 U61 ( .IN1(n13), .IN2(state[2]), .QN(n186) );
  INVX0 U62 ( .INP(n176), .ZN(ena_mac_wait) );
  NBUFFX2 U63 ( .INP(is_first_layer), .Z(input_or_int_mem_sel) );
  NOR2X0 U64 ( .IN1(ena_wr_int_mem_BAR), .IN2(n51), .QN(ena_wr_output_mem) );
  NOR2X0 U65 ( .IN1(n68), .IN2(n69), .QN(N242) );
  NOR2X0 U66 ( .IN1(counter_mac_wait[3]), .IN2(n177), .QN(n68) );
  NOR2X0 U67 ( .IN1(n60), .IN2(n61), .QN(N294) );
  NOR2X0 U68 ( .IN1(n206), .IN2(counter_wr_int_mem[3]), .QN(n60) );
  NOR2X0 U69 ( .IN1(n84), .IN2(n85), .QN(N174) );
  NOR2X0 U70 ( .IN1(counter_setup[2]), .IN2(n126), .QN(n84) );
  NOR2X0 U71 ( .IN1(n82), .IN2(n83), .QN(N177) );
  NOR2X0 U72 ( .IN1(n132), .IN2(counter_setup[5]), .QN(n82) );
  NOR2X0 U73 ( .IN1(n86), .IN2(n87), .QN(N173) );
  NOR2X0 U74 ( .IN1(counter_setup[0]), .IN2(counter_setup[1]), .QN(n86) );
  NOR2X0 U75 ( .IN1(n92), .IN2(n93), .QN(N147) );
  NOR2X0 U76 ( .IN1(counter_rd_user_para[0]), .IN2(counter_rd_user_para[1]), 
        .QN(n92) );
  NOR2X0 U77 ( .IN1(n90), .IN2(n91), .QN(N149) );
  NOR2X0 U78 ( .IN1(n99), .IN2(counter_rd_user_para[3]), .QN(n90) );
  NOR2X0 U79 ( .IN1(n88), .IN2(n89), .QN(N151) );
  NOR2X0 U80 ( .IN1(n102), .IN2(counter_rd_user_para[5]), .QN(n88) );
  NOR2X0 U81 ( .IN1(n58), .IN2(n59), .QN(N296) );
  NOR2X0 U82 ( .IN1(n209), .IN2(counter_wr_int_mem[5]), .QN(n58) );
  NOR2X0 U83 ( .IN1(n70), .IN2(n71), .QN(N240) );
  NOR2X0 U84 ( .IN1(counter_mac_wait[0]), .IN2(counter_mac_wait[1]), .QN(n70)
         );
  NOR2X0 U85 ( .IN1(n66), .IN2(n67), .QN(N244) );
  NOR2X0 U86 ( .IN1(n180), .IN2(counter_mac_wait[5]), .QN(n66) );
  NOR2X0 U87 ( .IN1(n80), .IN2(n81), .QN(N209) );
  NOR2X0 U88 ( .IN1(counter_mac[1]), .IN2(counter_mac[0]), .QN(n80) );
  NOR2X0 U89 ( .IN1(n78), .IN2(n79), .QN(N211) );
  NOR2X0 U90 ( .IN1(n156), .IN2(counter_mac[3]), .QN(n78) );
  NOR2X0 U91 ( .IN1(n76), .IN2(n77), .QN(N213) );
  NOR2X0 U92 ( .IN1(n159), .IN2(counter_mac[5]), .QN(n76) );
  NOR2X0 U93 ( .IN1(n74), .IN2(n75), .QN(N215) );
  NOR2X0 U94 ( .IN1(n162), .IN2(counter_mac[7]), .QN(n74) );
  NOR2X0 U95 ( .IN1(n62), .IN2(n63), .QN(N270) );
  NOR2X0 U96 ( .IN1(n195), .IN2(counter_act_func[5]), .QN(n62) );
  NOR2X0 U97 ( .IN1(n64), .IN2(n65), .QN(N268) );
  NOR2X0 U98 ( .IN1(n192), .IN2(counter_act_func[3]), .QN(n64) );
  NOR2X0 U99 ( .IN1(n72), .IN2(n73), .QN(N217) );
  NOR2X0 U100 ( .IN1(n165), .IN2(counter_mac[9]), .QN(n72) );
  NAND2X0 U101 ( .IN1(n13), .IN2(refresh_mac), .QN(n95) );
  INVX0 U102 ( .INP(n95), .ZN(ena_rd_user_para) );
  OR4X1 U103 ( .IN1(counter_rd_user_para[4]), .IN2(counter_rd_user_para[7]), 
        .IN3(counter_rd_user_para[3]), .IN4(counter_rd_user_para[5]), .Q(n94)
         );
  NOR4X0 U104 ( .IN1(counter_rd_user_para[2]), .IN2(counter_rd_user_para[6]), 
        .IN3(n98), .IN4(n94), .QN(n237) );
  NOR2X0 U105 ( .IN1(n237), .IN2(n95), .QN(n105) );
  INVX0 U106 ( .INP(n105), .ZN(n96) );
  NOR2X0 U107 ( .IN1(counter_rd_user_para[0]), .IN2(n96), .QN(N146) );
  INVX0 U108 ( .INP(n98), .ZN(n97) );
  OA221X1 U109 ( .IN1(counter_rd_user_para[2]), .IN2(n97), .IN3(n23), .IN4(n98), .IN5(n105), .Q(N148) );
  NOR2X0 U110 ( .IN1(n23), .IN2(n98), .QN(n99) );
  NAND4X0 U111 ( .IN1(counter_rd_user_para[2]), .IN2(counter_rd_user_para[1]), 
        .IN3(counter_rd_user_para[0]), .IN4(counter_rd_user_para[3]), .QN(n101) );
  INVX0 U112 ( .INP(n101), .ZN(n100) );
  OA221X1 U113 ( .IN1(counter_rd_user_para[4]), .IN2(n100), .IN3(n26), .IN4(
        n101), .IN5(n105), .Q(N150) );
  NOR2X0 U114 ( .IN1(n26), .IN2(n101), .QN(n102) );
  NOR2X0 U115 ( .IN1(n36), .IN2(n103), .QN(n107) );
  INVX0 U116 ( .INP(n107), .ZN(n106) );
  AND3X1 U117 ( .IN1(n106), .IN2(n105), .IN3(n104), .Q(N152) );
  OA221X1 U118 ( .IN1(counter_rd_user_para[7]), .IN2(n107), .IN3(n54), .IN4(
        n106), .IN5(n105), .Q(N153) );
  NAND3X0 U119 ( .IN1(counter_setup[1]), .IN2(counter_setup[0]), .IN3(
        counter_setup[2]), .QN(n127) );
  OR4X1 U120 ( .IN1(counter_setup[4]), .IN2(counter_setup[7]), .IN3(
        counter_setup[3]), .IN4(counter_setup[5]), .Q(n108) );
  NOR3X0 U121 ( .IN1(counter_setup[6]), .IN2(n127), .IN3(n108), .QN(n235) );
  NOR2X0 U122 ( .IN1(n235), .IN2(n43), .QN(n135) );
  INVX0 U123 ( .INP(n135), .ZN(n130) );
  NOR2X0 U124 ( .IN1(counter_setup[0]), .IN2(n130), .QN(N172) );
  INVX0 U125 ( .INP(n125), .ZN(n126) );
  INVX0 U126 ( .INP(n127), .ZN(n129) );
  OA221X1 U127 ( .IN1(n129), .IN2(counter_setup[3]), .IN3(n127), .IN4(n25), 
        .IN5(n135), .Q(N175) );
  NOR2X0 U128 ( .IN1(n127), .IN2(n25), .QN(n128) );
  NOR2X0 U129 ( .IN1(n128), .IN2(counter_setup[4]), .QN(n131) );
  AND3X1 U130 ( .IN1(n129), .IN2(counter_setup[4]), .IN3(counter_setup[3]), 
        .Q(n132) );
  NOR3X0 U131 ( .IN1(n131), .IN2(n132), .IN3(n130), .QN(N176) );
  NOR2X0 U132 ( .IN1(n35), .IN2(n133), .QN(n137) );
  INVX0 U133 ( .INP(n137), .ZN(n136) );
  AND3X1 U134 ( .IN1(n136), .IN2(n135), .IN3(n134), .Q(N178) );
  OA221X1 U135 ( .IN1(counter_setup[7]), .IN2(n137), .IN3(n55), .IN4(n136), 
        .IN5(n135), .Q(N179) );
  MUX21X1 U136 ( .IN1(n15), .IN2(counter_mac[8]), .S(mac_time[8]), .Q(n141) );
  MUX21X1 U137 ( .IN1(n16), .IN2(counter_mac[10]), .S(mac_time[10]), .Q(n140)
         );
  MUX21X1 U138 ( .IN1(n45), .IN2(counter_mac[9]), .S(mac_time[9]), .Q(n139) );
  MUX21X1 U139 ( .IN1(n46), .IN2(counter_mac[5]), .S(mac_time[5]), .Q(n138) );
  NAND4X0 U140 ( .IN1(n141), .IN2(n140), .IN3(n139), .IN4(n138), .QN(n152) );
  MUX21X1 U141 ( .IN1(n47), .IN2(counter_mac[7]), .S(mac_time[7]), .Q(n145) );
  MUX21X1 U142 ( .IN1(n12), .IN2(counter_mac[6]), .S(mac_time[6]), .Q(n144) );
  MUX21X1 U143 ( .IN1(n10), .IN2(counter_mac[2]), .S(mac_time[2]), .Q(n143) );
  MUX21X1 U144 ( .IN1(n11), .IN2(counter_mac[4]), .S(mac_time[4]), .Q(n142) );
  NAND4X0 U145 ( .IN1(n145), .IN2(n144), .IN3(n143), .IN4(n142), .QN(n151) );
  MUX21X1 U146 ( .IN1(n48), .IN2(counter_mac[3]), .S(mac_time[3]), .Q(n149) );
  MUX21X1 U147 ( .IN1(n22), .IN2(counter_mac[0]), .S(mac_time[0]), .Q(n148) );
  MUX21X1 U148 ( .IN1(n50), .IN2(counter_mac[1]), .S(mac_time[1]), .Q(n147) );
  MUX21X1 U149 ( .IN1(n32), .IN2(counter_mac[11]), .S(mac_time[11]), .Q(n146)
         );
  NAND4X0 U150 ( .IN1(n149), .IN2(n148), .IN3(n147), .IN4(n146), .QN(n150) );
  NOR3X0 U151 ( .IN1(n152), .IN2(n151), .IN3(n150), .QN(n229) );
  INVX0 U152 ( .INP(ena_mac), .ZN(n153) );
  AND2X1 U153 ( .IN1(n22), .IN2(n168), .Q(N208) );
  INVX0 U154 ( .INP(n155), .ZN(n154) );
  OA221X1 U155 ( .IN1(counter_mac[2]), .IN2(n154), .IN3(n10), .IN4(n155), 
        .IN5(n168), .Q(N210) );
  NOR2X0 U156 ( .IN1(n10), .IN2(n155), .QN(n156) );
  INVX0 U157 ( .INP(n158), .ZN(n157) );
  OA221X1 U158 ( .IN1(counter_mac[4]), .IN2(n157), .IN3(n11), .IN4(n158), 
        .IN5(n168), .Q(N212) );
  NOR2X0 U159 ( .IN1(n11), .IN2(n158), .QN(n159) );
  INVX0 U160 ( .INP(n161), .ZN(n160) );
  OA221X1 U161 ( .IN1(counter_mac[6]), .IN2(n160), .IN3(n12), .IN4(n161), 
        .IN5(n168), .Q(N214) );
  NOR2X0 U162 ( .IN1(n12), .IN2(n161), .QN(n162) );
  INVX0 U163 ( .INP(n164), .ZN(n163) );
  OA221X1 U164 ( .IN1(counter_mac[8]), .IN2(n163), .IN3(n15), .IN4(n164), 
        .IN5(n168), .Q(N216) );
  NOR2X0 U165 ( .IN1(n15), .IN2(n164), .QN(n165) );
  NOR2X0 U166 ( .IN1(n16), .IN2(n166), .QN(n170) );
  INVX0 U167 ( .INP(n170), .ZN(n169) );
  AND3X1 U168 ( .IN1(n169), .IN2(n168), .IN3(n167), .Q(N218) );
  OA221X1 U169 ( .IN1(counter_mac[11]), .IN2(n170), .IN3(n32), .IN4(n169), 
        .IN5(n168), .Q(N219) );
  AND3X1 U170 ( .IN1(counter_mac_wait[1]), .IN2(counter_mac_wait[0]), .IN3(
        counter_mac_wait[2]), .Q(n177) );
  OR4X1 U171 ( .IN1(counter_mac_wait[7]), .IN2(counter_mac_wait[4]), .IN3(
        counter_mac_wait[6]), .IN4(counter_mac_wait[5]), .Q(n171) );
  NOR2X0 U172 ( .IN1(n179), .IN2(n171), .QN(n236) );
  NOR2X0 U173 ( .IN1(n236), .IN2(n176), .QN(n183) );
  INVX0 U174 ( .INP(n183), .ZN(n174) );
  NOR2X0 U175 ( .IN1(counter_mac_wait[0]), .IN2(n174), .QN(N239) );
  INVX0 U176 ( .INP(n172), .ZN(n173) );
  NOR2X0 U177 ( .IN1(counter_mac_wait[2]), .IN2(n173), .QN(n175) );
  NOR3X0 U178 ( .IN1(n175), .IN2(n177), .IN3(n174), .QN(N241) );
  INVX0 U179 ( .INP(n179), .ZN(n178) );
  OA221X1 U180 ( .IN1(n178), .IN2(counter_mac_wait[4]), .IN3(n179), .IN4(n30), 
        .IN5(n183), .Q(N243) );
  NOR2X0 U181 ( .IN1(n179), .IN2(n30), .QN(n180) );
  NOR2X0 U182 ( .IN1(n33), .IN2(n181), .QN(n185) );
  INVX0 U183 ( .INP(n185), .ZN(n184) );
  AND3X1 U184 ( .IN1(n184), .IN2(n183), .IN3(n182), .Q(N245) );
  OA221X1 U185 ( .IN1(counter_mac_wait[7]), .IN2(n185), .IN3(n53), .IN4(n184), 
        .IN5(n183), .Q(N246) );
  NOR2X0 U186 ( .IN1(counter_act_func[0]), .IN2(counter_act_func[1]), .QN(n188) );
  NOR4X0 U187 ( .IN1(counter_act_func[7]), .IN2(counter_act_func[2]), .IN3(
        counter_act_func[4]), .IN4(counter_act_func[6]), .QN(n187) );
  NAND4X0 U188 ( .IN1(n188), .IN2(counter_act_func[5]), .IN3(
        counter_act_func[3]), .IN4(n187), .QN(n231) );
  NOR2X0 U189 ( .IN1(counter_act_func[0]), .IN2(n191), .QN(N265) );
  AND2X1 U190 ( .IN1(counter_act_func[0]), .IN2(counter_act_func[1]), .Q(n189)
         );
  NOR3X0 U191 ( .IN1(n188), .IN2(n189), .IN3(n191), .QN(N266) );
  NOR2X0 U192 ( .IN1(n189), .IN2(counter_act_func[2]), .QN(n190) );
  AND3X1 U193 ( .IN1(counter_act_func[0]), .IN2(counter_act_func[1]), .IN3(
        counter_act_func[2]), .Q(n192) );
  NOR3X0 U194 ( .IN1(n190), .IN2(n192), .IN3(n191), .QN(N267) );
  INVX0 U195 ( .INP(n191), .ZN(n198) );
  INVX0 U196 ( .INP(n194), .ZN(n193) );
  OA221X1 U197 ( .IN1(counter_act_func[4]), .IN2(n193), .IN3(n28), .IN4(n194), 
        .IN5(n198), .Q(N269) );
  NOR2X0 U198 ( .IN1(n28), .IN2(n194), .QN(n195) );
  NOR2X0 U199 ( .IN1(n37), .IN2(n196), .QN(n200) );
  INVX0 U200 ( .INP(n200), .ZN(n199) );
  AND3X1 U201 ( .IN1(n199), .IN2(n198), .IN3(n197), .Q(N271) );
  OA221X1 U202 ( .IN1(counter_act_func[7]), .IN2(n200), .IN3(n52), .IN4(n199), 
        .IN5(n198), .Q(N272) );
  NOR2X0 U203 ( .IN1(counter_wr_int_mem[0]), .IN2(ena_wr_int_mem_BAR), .QN(
        N291) );
  OR4X1 U204 ( .IN1(counter_wr_int_mem[3]), .IN2(counter_wr_int_mem[4]), .IN3(
        counter_wr_int_mem[5]), .IN4(counter_wr_int_mem[6]), .Q(n201) );
  NOR4X0 U205 ( .IN1(counter_wr_int_mem[2]), .IN2(counter_wr_int_mem[7]), 
        .IN3(n202), .IN4(n201), .QN(n230) );
  NOR2X0 U206 ( .IN1(n230), .IN2(ena_wr_int_mem_BAR), .QN(n212) );
  OA222X1 U207 ( .IN1(counter_wr_int_mem[1]), .IN2(counter_wr_int_mem[0]), 
        .IN3(counter_wr_int_mem[1]), .IN4(n212), .IN5(N291), .IN6(n39), .Q(
        N292) );
  AND3X1 U208 ( .IN1(counter_wr_int_mem[1]), .IN2(counter_wr_int_mem[0]), 
        .IN3(counter_wr_int_mem[2]), .Q(n206) );
  AND2X1 U209 ( .IN1(counter_wr_int_mem[1]), .IN2(counter_wr_int_mem[0]), .Q(
        n203) );
  NOR2X0 U210 ( .IN1(counter_wr_int_mem[2]), .IN2(n203), .QN(n205) );
  INVX0 U211 ( .INP(n212), .ZN(n204) );
  NOR3X0 U212 ( .IN1(n206), .IN2(n205), .IN3(n204), .QN(N293) );
  INVX0 U213 ( .INP(n208), .ZN(n207) );
  OA221X1 U214 ( .IN1(counter_wr_int_mem[4]), .IN2(n207), .IN3(n27), .IN4(n208), .IN5(n212), .Q(N295) );
  NOR2X0 U215 ( .IN1(n27), .IN2(n208), .QN(n209) );
  NOR2X0 U216 ( .IN1(n34), .IN2(n210), .QN(n214) );
  INVX0 U217 ( .INP(n214), .ZN(n213) );
  AND3X1 U218 ( .IN1(n213), .IN2(n212), .IN3(n211), .Q(N297) );
  OA221X1 U219 ( .IN1(counter_wr_int_mem[7]), .IN2(n214), .IN3(n56), .IN4(n213), .IN5(n212), .Q(N298) );
  MUX21X1 U220 ( .IN1(node_counter[3]), .IN2(n41), .S(
        num_of_node_for_each_layer[3]), .Q(n223) );
  MUX21X1 U221 ( .IN1(node_counter[2]), .IN2(n40), .S(
        num_of_node_for_each_layer[2]), .Q(n222) );
  OAI22X1 U222 ( .IN1(num_of_node_for_each_layer[5]), .IN2(n38), .IN3(n8), 
        .IN4(num_of_node_for_each_layer[6]), .QN(n215) );
  AO221X1 U223 ( .IN1(n38), .IN2(num_of_node_for_each_layer[5]), .IN3(n8), 
        .IN4(num_of_node_for_each_layer[6]), .IN5(n215), .Q(n221) );
  MUX21X1 U224 ( .IN1(n17), .IN2(node_counter[1]), .S(
        num_of_node_for_each_layer[1]), .Q(n219) );
  MUX21X1 U225 ( .IN1(n6), .IN2(node_counter[0]), .S(
        num_of_node_for_each_layer[0]), .Q(n218) );
  MUX21X1 U226 ( .IN1(n20), .IN2(node_counter[4]), .S(
        num_of_node_for_each_layer[4]), .Q(n217) );
  MUX21X1 U227 ( .IN1(n31), .IN2(node_counter[7]), .S(
        num_of_node_for_each_layer[7]), .Q(n216) );
  NAND4X0 U228 ( .IN1(n219), .IN2(n218), .IN3(n217), .IN4(n216), .QN(n220) );
  NOR4X0 U229 ( .IN1(n223), .IN2(n222), .IN3(n221), .IN4(n220), .QN(n257) );
  INVX0 U230 ( .INP(n262), .ZN(n256) );
  AND2X1 U231 ( .IN1(n257), .IN2(n256), .Q(N320) );
  MUX21X1 U232 ( .IN1(layer_counter[0]), .IN2(n44), .S(num_of_layer[0]), .Q(
        n227) );
  MUX21X1 U233 ( .IN1(layer_counter[3]), .IN2(n24), .S(num_of_layer[3]), .Q(
        n226) );
  MUX21X1 U234 ( .IN1(layer_counter[1]), .IN2(n19), .S(num_of_layer[1]), .Q(
        n225) );
  MUX21X1 U235 ( .IN1(layer_counter[2]), .IN2(n7), .S(num_of_layer[2]), .Q(
        n224) );
  NOR4X0 U236 ( .IN1(n227), .IN2(n226), .IN3(n225), .IN4(n224), .QN(n228) );
  MUX21X1 U237 ( .IN1(n228), .IN2(is_last_layer), .S(n43), .Q(N334) );
  INVX0 U238 ( .INP(n230), .ZN(n232) );
  NAND3X0 U239 ( .IN1(n233), .IN2(n232), .IN3(n231), .QN(n234) );
  NOR4X0 U240 ( .IN1(n237), .IN2(n236), .IN3(n235), .IN4(n234), .QN(n245) );
  INVX0 U241 ( .INP(n245), .ZN(n247) );
  NAND3X0 U242 ( .IN1(state[1]), .IN2(n247), .IN3(n5), .QN(n238) );
  NAND2X0 U243 ( .IN1(n238), .IN2(state[2]), .QN(n239) );
  OAI21X1 U244 ( .IN1(n240), .IN2(n43), .IN3(n239), .QN(n124) );
  AO222X1 U245 ( .IN1(state[2]), .IN2(state[1]), .IN3(state[2]), .IN4(n245), 
        .IN5(state[1]), .IN6(n241), .Q(n242) );
  NOR2X0 U246 ( .IN1(n13), .IN2(n242), .QN(n243) );
  OA21X1 U247 ( .IN1(n13), .IN2(state[2]), .IN3(state[1]), .Q(n244) );
  OR2X1 U248 ( .IN1(state[1]), .IN2(state[2]), .Q(n246) );
  OA22X1 U249 ( .IN1(n243), .IN2(n244), .IN3(ena_neural), .IN4(n246), .Q(n123)
         );
  OAI22X1 U250 ( .IN1(ena_mac), .IN2(n244), .IN3(n5), .IN4(n247), .QN(n251) );
  AO21X1 U251 ( .IN1(ena_neural), .IN2(n5), .IN3(n246), .Q(n249) );
  AO221X1 U252 ( .IN1(n42), .IN2(change_layer), .IN3(n42), .IN4(n247), .IN5(
        n43), .Q(n248) );
  NAND4X0 U253 ( .IN1(n251), .IN2(n250), .IN3(n249), .IN4(n248), .QN(n122) );
  NOR2X0 U254 ( .IN1(n257), .IN2(n262), .QN(n269) );
  MUX21X1 U255 ( .IN1(n269), .IN2(n262), .S(node_counter[0]), .Q(n121) );
  INVX0 U256 ( .INP(n269), .ZN(n263) );
  NOR2X0 U257 ( .IN1(node_counter[1]), .IN2(n263), .QN(n255) );
  AO22X1 U258 ( .IN1(node_counter[1]), .IN2(n254), .IN3(node_counter[0]), 
        .IN4(n255), .Q(n120) );
  NOR4X0 U259 ( .IN1(node_counter[2]), .IN2(n17), .IN3(n6), .IN4(n263), .QN(
        n253) );
  AO221X1 U260 ( .IN1(node_counter[2]), .IN2(n255), .IN3(node_counter[2]), 
        .IN4(n254), .IN5(n253), .Q(n119) );
  AND3X1 U261 ( .IN1(node_counter[2]), .IN2(node_counter[1]), .IN3(
        node_counter[0]), .Q(n261) );
  OAI21X1 U262 ( .IN1(n257), .IN2(n261), .IN3(n256), .QN(n259) );
  NOR2X0 U263 ( .IN1(node_counter[3]), .IN2(n263), .QN(n260) );
  AO22X1 U264 ( .IN1(node_counter[3]), .IN2(n259), .IN3(n261), .IN4(n260), .Q(
        n118) );
  AND3X1 U265 ( .IN1(node_counter[3]), .IN2(n269), .IN3(n261), .Q(n258) );
  AO222X1 U266 ( .IN1(node_counter[4]), .IN2(n260), .IN3(node_counter[4]), 
        .IN4(n259), .IN5(n258), .IN6(n20), .Q(n117) );
  NAND3X0 U267 ( .IN1(node_counter[3]), .IN2(node_counter[4]), .IN3(n261), 
        .QN(n264) );
  AO21X1 U268 ( .IN1(n269), .IN2(n264), .IN3(n262), .Q(n266) );
  NOR2X0 U269 ( .IN1(node_counter[5]), .IN2(n263), .QN(n267) );
  INVX0 U270 ( .INP(n264), .ZN(n265) );
  AO22X1 U271 ( .IN1(node_counter[5]), .IN2(n266), .IN3(n267), .IN4(n265), .Q(
        n116) );
  AND3X1 U272 ( .IN1(node_counter[5]), .IN2(n269), .IN3(n265), .Q(n271) );
  OR2X1 U273 ( .IN1(n267), .IN2(n266), .Q(n268) );
  MUX21X1 U274 ( .IN1(n271), .IN2(n268), .S(node_counter[6]), .Q(n115) );
  AO21X1 U275 ( .IN1(n8), .IN2(n269), .IN3(n268), .Q(n270) );
  OA222X1 U276 ( .IN1(node_counter[7]), .IN2(node_counter[6]), .IN3(
        node_counter[7]), .IN4(n271), .IN5(n31), .IN6(n270), .Q(n114) );
  NAND2X0 U277 ( .IN1(change_layer), .IN2(layer_counter[0]), .QN(n272) );
  AO221X1 U278 ( .IN1(n272), .IN2(change_layer), .IN3(n272), .IN4(
        layer_counter[0]), .IN5(ena_neural), .Q(n113) );
  INVX0 U279 ( .INP(ena_neural), .ZN(n276) );
  NAND3X0 U280 ( .IN1(change_layer), .IN2(layer_counter[1]), .IN3(
        layer_counter[0]), .QN(n277) );
  NAND3X0 U281 ( .IN1(n273), .IN2(n276), .IN3(n277), .QN(n29) );
  INVX0 U282 ( .INP(n277), .ZN(n274) );
  OA221X1 U283 ( .IN1(layer_counter[2]), .IN2(n274), .IN3(n7), .IN4(n277), 
        .IN5(n276), .Q(n112) );
  AND3X1 U284 ( .IN1(layer_counter[2]), .IN2(layer_counter[1]), .IN3(
        layer_counter[0]), .Q(n275) );
  OA221X1 U285 ( .IN1(layer_counter[3]), .IN2(n275), .IN3(n24), .IN4(n7), 
        .IN5(change_layer), .Q(n278) );
  OA221X1 U286 ( .IN1(n278), .IN2(layer_counter[3]), .IN3(n278), .IN4(n277), 
        .IN5(n276), .Q(n111) );
  AO21X1 U287 ( .IN1(is_first_layer), .IN2(n18), .IN3(ena_neural), .Q(n110) );
  AO221X1 U288 ( .IN1(change_layer), .IN2(n21), .IN3(n18), .IN4(is_odd_layer), 
        .IN5(ena_neural), .Q(n109) );
endmodule


module para_controller ( clk, rst_n, ena_rd_user_para, is_first_layer, 
        para_addr, para_cof );
  output [19:0] para_addr;
  output [3:0] para_cof;
  input clk, rst_n, ena_rd_user_para, is_first_layer;
  wire   ena_rd_user_para_w1, N77, N78, N79, N80, n1, n2, n3, n5, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n4, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  DFFARX1 ena_rd_user_para_w1_reg ( .D(ena_rd_user_para), .CLK(clk), .RSTB(
        rst_n), .Q(ena_rd_user_para_w1), .QN(n3) );
  DFFARX1 para_addr_reg_9_ ( .D(n23), .CLK(clk), .RSTB(rst_n), .Q(para_addr[9]), .QN(n12) );
  DFFARX1 para_addr_reg_8_ ( .D(n24), .CLK(clk), .RSTB(rst_n), .Q(para_addr[8]) );
  DFFARX1 para_addr_reg_7_ ( .D(n25), .CLK(clk), .RSTB(rst_n), .Q(para_addr[7]), .QN(n6) );
  DFFARX1 para_addr_reg_6_ ( .D(n26), .CLK(clk), .RSTB(rst_n), .Q(para_addr[6]), .QN(n9) );
  DFFARX1 para_addr_reg_5_ ( .D(n27), .CLK(clk), .RSTB(rst_n), .Q(para_addr[5]), .QN(n4) );
  DFFARX1 para_addr_reg_4_ ( .D(n28), .CLK(clk), .RSTB(rst_n), .Q(para_addr[4]), .QN(n10) );
  DFFARX1 para_addr_reg_3_ ( .D(n29), .CLK(clk), .RSTB(rst_n), .Q(para_addr[3]), .QN(n7) );
  DFFARX1 para_addr_reg_2_ ( .D(n30), .CLK(clk), .RSTB(rst_n), .Q(para_addr[2]), .QN(n11) );
  DFFARX1 para_addr_reg_1_ ( .D(n31), .CLK(clk), .RSTB(rst_n), .Q(para_addr[1]), .QN(n8) );
  DFFARX1 para_addr_reg_0_ ( .D(n32), .CLK(clk), .RSTB(rst_n), .Q(para_addr[0]) );
  DFFASX1 ena_rd_user_para_w3_reg ( .D(n3), .CLK(clk), .SETB(rst_n), .Q(n2) );
  DFFASX1 ena_rd_user_para_w4_reg ( .D(n2), .CLK(clk), .SETB(rst_n), .Q(n1) );
  DFFASX1 ena_rd_user_para_w5_reg ( .D(n1), .CLK(clk), .SETB(rst_n), .Q(n5), 
        .QN(n14) );
  DFFARX1 para_cof_reg_0_ ( .D(N77), .CLK(clk), .RSTB(rst_n), .Q(para_cof[0])
         );
  DFFARX1 para_cof_reg_1_ ( .D(N78), .CLK(clk), .RSTB(rst_n), .Q(para_cof[1])
         );
  DFFARX1 para_cof_reg_2_ ( .D(N79), .CLK(clk), .RSTB(rst_n), .Q(para_cof[2])
         );
  DFFARX1 para_cof_reg_3_ ( .D(N80), .CLK(clk), .RSTB(rst_n), .Q(para_cof[3]), 
        .QN(n13) );
  NAND2X0 U3 ( .IN1(para_addr[0]), .IN2(n35), .QN(n20) );
  NAND2X0 U4 ( .IN1(n36), .IN2(n35), .QN(n38) );
  NAND2X0 U5 ( .IN1(para_addr[6]), .IN2(n39), .QN(n40) );
  NAND2X0 U6 ( .IN1(para_addr[8]), .IN2(n41), .QN(n42) );
  NAND2X0 U7 ( .IN1(n34), .IN2(n35), .QN(n22) );
  NOR2X0 U8 ( .IN1(n5), .IN2(para_cof[0]), .QN(N77) );
  NOR2X0 U9 ( .IN1(n5), .IN2(para_cof[1]), .QN(n15) );
  AO22X1 U10 ( .IN1(para_cof[1]), .IN2(N77), .IN3(n15), .IN4(para_cof[0]), .Q(
        N78) );
  AND3X1 U11 ( .IN1(para_cof[1]), .IN2(para_cof[0]), .IN3(n14), .Q(n19) );
  OR2X1 U12 ( .IN1(n15), .IN2(N77), .Q(n16) );
  MUX21X1 U13 ( .IN1(n19), .IN2(n16), .S(para_cof[2]), .Q(N79) );
  AND3X1 U14 ( .IN1(para_cof[2]), .IN2(para_cof[1]), .IN3(para_cof[0]), .Q(n17) );
  NOR2X0 U15 ( .IN1(n17), .IN2(n5), .QN(n18) );
  OA222X1 U16 ( .IN1(para_cof[3]), .IN2(para_cof[2]), .IN3(para_cof[3]), .IN4(
        n19), .IN5(n13), .IN6(n18), .Q(N80) );
  OA21X1 U17 ( .IN1(ena_rd_user_para_w1), .IN2(is_first_layer), .IN3(
        ena_rd_user_para), .Q(n35) );
  OA21X1 U18 ( .IN1(para_addr[0]), .IN2(n35), .IN3(n20), .Q(n32) );
  MUX21X1 U19 ( .IN1(n8), .IN2(para_addr[1]), .S(n20), .Q(n31) );
  NAND3X0 U20 ( .IN1(para_addr[1]), .IN2(para_addr[0]), .IN3(n35), .QN(n21) );
  MUX21X1 U21 ( .IN1(n11), .IN2(para_addr[2]), .S(n21), .Q(n30) );
  AND3X1 U22 ( .IN1(para_addr[2]), .IN2(para_addr[1]), .IN3(para_addr[0]), .Q(
        n34) );
  MUX21X1 U23 ( .IN1(n7), .IN2(para_addr[3]), .S(n22), .Q(n29) );
  NAND3X0 U24 ( .IN1(n34), .IN2(para_addr[3]), .IN3(n35), .QN(n33) );
  MUX21X1 U25 ( .IN1(n10), .IN2(para_addr[4]), .S(n33), .Q(n28) );
  AND3X1 U26 ( .IN1(n34), .IN2(para_addr[4]), .IN3(para_addr[3]), .Q(n36) );
  MUX21X1 U27 ( .IN1(n4), .IN2(para_addr[5]), .S(n38), .Q(n27) );
  OR2X1 U28 ( .IN1(n4), .IN2(n38), .Q(n37) );
  MUX21X1 U29 ( .IN1(n9), .IN2(para_addr[6]), .S(n37), .Q(n26) );
  NOR2X0 U30 ( .IN1(n4), .IN2(n38), .QN(n39) );
  MUX21X1 U31 ( .IN1(n6), .IN2(para_addr[7]), .S(n40), .Q(n25) );
  NOR2X0 U32 ( .IN1(n40), .IN2(n6), .QN(n41) );
  OA21X1 U33 ( .IN1(para_addr[8]), .IN2(n41), .IN3(n42), .Q(n24) );
  MUX21X1 U34 ( .IN1(n12), .IN2(para_addr[9]), .S(n42), .Q(n23) );
endmodule


module neural ( clk, rst_n, enable_neural, disable_neural, user_para_data, 
        user_para_addr, int_mem_addr_rd, input_mem_addr, w_addr, 
        int_mem_addr_wr, output_mem_addr, int_mem_data_rd, input_mem_data, 
        w_data, int_mem_data_wr, output_data, wr_ena_int_n_BAR, 
        wr_ena_out_n_BAR );
  input [31:0] user_para_data;
  output [19:0] user_para_addr;
  output [19:0] int_mem_addr_rd;
  output [19:0] input_mem_addr;
  output [19:0] w_addr;
  output [19:0] int_mem_addr_wr;
  output [19:0] output_mem_addr;
  input [31:0] int_mem_data_rd;
  input [31:0] input_mem_data;
  input [31:0] w_data;
  output [31:0] int_mem_data_wr;
  output [31:0] output_data;
  input clk, rst_n, enable_neural;
  output disable_neural, wr_ena_int_n_BAR, wr_ena_out_n_BAR;
  wire   ena_neural, end_neural, ena_wr_output_mem, ena_wr_int_mem,
         is_odd_layer, is_first_layer, ena_mac, ena_mac_wait, ena_mac_delay,
         ena_mul_add, input_or_int_mem_sel, N91, N92, N93, N94, N95, N96, N97,
         N98, N99, N100, N101, N102, N103, N104, N105, N106, N107, N108, N109,
         N110, N111, N112, N113, N114, N115, N116, N117, N118, N119, N120,
         N121, N122, N126, N127, N128, N129, N130, N131, N132, N133, N134,
         N135, N136, N137, N138, N139, N140, N141, N142, N143, N144, N145,
         N146, N147, N148, N149, N150, N151, N152, N153, N154, N155, N156,
         N157, refresh_mac, ena_act_func, N160, N161, N162, N163, N164, N165,
         N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176,
         N177, N178, N179, N180, N181, N182, N183, N184, N185, N186, N187,
         N188, N189, N190, N191, step_output_23_, N235, N236, N237, N238, N239,
         N240, N241, N242, N243, N244, N245, N246, N247, N248, N249, N250,
         N251, N252, N253, N254, N255, N256, N257, N258, N259, N260, N261,
         N262, N263, N264, N265, N266, change_layer, N272, N273, N274, N275,
         N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286,
         N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N307, N308, N309, N310, N311,
         N312, N313, N314, N315, N316, N317, N318, N319, N320, N321, N322,
         N323, N324, N325, N326, N327, N328, N329, N330, N331, N332, N333,
         N334, N335, N336, N337, N338, ena_rd_user_para, N347, N348, N349,
         N350, N351, N352, N353, N354, N355, N356, N357, N358, N359, N360,
         N361, N362, N363, N364, N365, N366, N367, N368, N369, N370, N371,
         N372, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22,
         SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24,
         SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26,
         SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28,
         SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30,
         SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32,
         SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34,
         SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36,
         SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38,
         SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40,
         SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42,
         SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44,
         SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46,
         SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48,
         SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50,
         SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52,
         SYNOPSYS_UNCONNECTED_53, SYNOPSYS_UNCONNECTED_54,
         SYNOPSYS_UNCONNECTED_55, SYNOPSYS_UNCONNECTED_56,
         SYNOPSYS_UNCONNECTED_57, SYNOPSYS_UNCONNECTED_58,
         SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_60,
         SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_62,
         SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_64,
         SYNOPSYS_UNCONNECTED_65, SYNOPSYS_UNCONNECTED_66,
         SYNOPSYS_UNCONNECTED_67, SYNOPSYS_UNCONNECTED_68,
         SYNOPSYS_UNCONNECTED_69, SYNOPSYS_UNCONNECTED_70,
         SYNOPSYS_UNCONNECTED_71, SYNOPSYS_UNCONNECTED_72;
  wire   [19:0] w_addr_w1;
  wire   [9:0] input_or_int_mem_addr;
  wire   [31:0] mac_input_01;
  wire   [31:0] mac_input_02;
  wire   [31:0] mac_output;
  wire   [31:0] input_act_func;
  wire   [31:0] linear_output;
  wire   [31:0] sigmoid_output;
  wire   [31:0] tansigmoid_output;
  wire   [1:0] act_function_sel;
  wire   [31:0] out_act_func;
  wire   [9:0] output_mem_addr_w1;
  wire   [9:0] int_mem_addr_wr_w1;
  wire   [11:0] mac_time;
  wire   [3:0] num_of_layer;
  wire   [7:0] num_of_node_for_each_layer;
  wire   [9:0] para_addr;
  wire   [3:0] para_cof;
  wire   [11:0] para_data;

  input_mac_controller input_mac_controller_01 ( .clk(clk), .rst_n(rst_n), 
        .is_odd_layer(is_odd_layer), .is_first_layer(is_first_layer), 
        .ena_mac(ena_mac), .ena_mac_wait(ena_mac_wait), .ena_mul_add(
        ena_mul_add), .ena_mac_delay(ena_mac_delay), .w_addr(w_addr_w1), 
        .input_or_int_mem_addr({SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, 
        SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, 
        SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, 
        SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10, input_or_int_mem_addr}) );
  mac mac_01 ( .clk(clk), .rst_n(rst_n), .refresh_mac(refresh_mac), .ena_mac(
        ena_mac_delay), .ena_mac_wait(ena_mac_wait), .ena_mul_add(ena_mul_add), 
        .mac_input_01(mac_input_01), .mac_input_02(mac_input_02), .mac_output(
        mac_output) );
  linear_function linear_function_01 ( .clk(clk), .rst_n(rst_n), 
        .linear_input(input_act_func), .linear_output({linear_output[31], 
        SYNOPSYS_UNCONNECTED_11, linear_output[29:0]}) );
  step_function step_function_01 ( .clk(clk), .rst_n(rst_n), .step_input({
        input_act_func[31], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .step_output({SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13, 
        SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, 
        SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17, 
        SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19, step_output_23_, 
        SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21, 
        SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_23, 
        SYNOPSYS_UNCONNECTED_24, SYNOPSYS_UNCONNECTED_25, 
        SYNOPSYS_UNCONNECTED_26, SYNOPSYS_UNCONNECTED_27, 
        SYNOPSYS_UNCONNECTED_28, SYNOPSYS_UNCONNECTED_29, 
        SYNOPSYS_UNCONNECTED_30, SYNOPSYS_UNCONNECTED_31, 
        SYNOPSYS_UNCONNECTED_32, SYNOPSYS_UNCONNECTED_33, 
        SYNOPSYS_UNCONNECTED_34, SYNOPSYS_UNCONNECTED_35, 
        SYNOPSYS_UNCONNECTED_36, SYNOPSYS_UNCONNECTED_37, 
        SYNOPSYS_UNCONNECTED_38, SYNOPSYS_UNCONNECTED_39, 
        SYNOPSYS_UNCONNECTED_40, SYNOPSYS_UNCONNECTED_41, 
        SYNOPSYS_UNCONNECTED_42}) );
  sigmoid_function sigmoid_function_01 ( .clk(clk), .rst_n(rst_n), 
        .sigmoid_input(input_act_func), .sigmoid_output(sigmoid_output) );
  tansigmoid_function tansigmoid_function_01 ( .clk(clk), .rst_n(rst_n), 
        .tansigmoid_input(input_act_func), .tansigmoid_output(
        tansigmoid_output) );
  wr_int_mem_controller wr_int_mem_controller_01 ( .clk(clk), .rst_n(rst_n), 
        .ena_wr_output_mem(ena_wr_output_mem), .is_odd_layer(is_odd_layer), 
        .is_first_layer(is_first_layer), .change_layer(change_layer), 
        .int_mem_addr_wr({SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44, 
        SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46, 
        SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48, 
        SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50, 
        SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52, int_mem_addr_wr_w1}), 
        .output_mem_addr({SYNOPSYS_UNCONNECTED_53, SYNOPSYS_UNCONNECTED_54, 
        SYNOPSYS_UNCONNECTED_55, SYNOPSYS_UNCONNECTED_56, 
        SYNOPSYS_UNCONNECTED_57, SYNOPSYS_UNCONNECTED_58, 
        SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_60, 
        SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_62, output_mem_addr_w1}), 
        .ena_wr_int_mem_BAR(ena_wr_int_mem) );
  network_control network_control_01 ( .clk(clk), .rst_n(rst_n), .ena_neural(
        ena_neural), .mac_time(mac_time), .num_of_layer(num_of_layer), 
        .num_of_node_for_each_layer(num_of_node_for_each_layer), 
        .ena_rd_user_para(ena_rd_user_para), .ena_mac(ena_mac), .ena_mac_wait(
        ena_mac_wait), .ena_act_func(ena_act_func), .input_or_int_mem_sel(
        input_or_int_mem_sel), .is_first_layer(is_first_layer), .is_odd_layer(
        is_odd_layer), .refresh_mac(refresh_mac), .change_layer(change_layer), 
        .ena_wr_output_mem(ena_wr_output_mem), .end_neural(end_neural), 
        .ena_wr_int_mem_BAR(ena_wr_int_mem) );
  para_controller para_controller_01 ( .clk(clk), .rst_n(rst_n), 
        .ena_rd_user_para(ena_rd_user_para), .is_first_layer(is_first_layer), 
        .para_addr({SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_64, 
        SYNOPSYS_UNCONNECTED_65, SYNOPSYS_UNCONNECTED_66, 
        SYNOPSYS_UNCONNECTED_67, SYNOPSYS_UNCONNECTED_68, 
        SYNOPSYS_UNCONNECTED_69, SYNOPSYS_UNCONNECTED_70, 
        SYNOPSYS_UNCONNECTED_71, SYNOPSYS_UNCONNECTED_72, para_addr}), 
        .para_cof(para_cof) );
  DFFARX1 ena_neural_reg ( .D(enable_neural), .CLK(clk), .RSTB(rst_n), .Q(
        ena_neural) );
  DFFARX1 para_data_reg_11_ ( .D(user_para_data[11]), .CLK(clk), .RSTB(rst_n), 
        .Q(para_data[11]) );
  DFFARX1 para_data_reg_10_ ( .D(user_para_data[10]), .CLK(clk), .RSTB(rst_n), 
        .Q(para_data[10]) );
  DFFARX1 para_data_reg_9_ ( .D(user_para_data[9]), .CLK(clk), .RSTB(rst_n), 
        .Q(para_data[9]) );
  DFFARX1 para_data_reg_8_ ( .D(user_para_data[8]), .CLK(clk), .RSTB(rst_n), 
        .Q(para_data[8]) );
  DFFARX1 para_data_reg_7_ ( .D(user_para_data[7]), .CLK(clk), .RSTB(rst_n), 
        .Q(para_data[7]) );
  DFFARX1 para_data_reg_6_ ( .D(user_para_data[6]), .CLK(clk), .RSTB(rst_n), 
        .Q(para_data[6]) );
  DFFARX1 para_data_reg_5_ ( .D(user_para_data[5]), .CLK(clk), .RSTB(rst_n), 
        .Q(para_data[5]) );
  DFFARX1 para_data_reg_4_ ( .D(user_para_data[4]), .CLK(clk), .RSTB(rst_n), 
        .Q(para_data[4]) );
  DFFARX1 para_data_reg_3_ ( .D(user_para_data[3]), .CLK(clk), .RSTB(rst_n), 
        .Q(para_data[3]) );
  DFFARX1 para_data_reg_2_ ( .D(user_para_data[2]), .CLK(clk), .RSTB(rst_n), 
        .Q(para_data[2]) );
  DFFARX1 para_data_reg_1_ ( .D(user_para_data[1]), .CLK(clk), .RSTB(rst_n), 
        .Q(para_data[1]) );
  DFFARX1 para_data_reg_0_ ( .D(user_para_data[0]), .CLK(clk), .RSTB(rst_n), 
        .Q(para_data[0]) );
  DFFARX1 num_of_layer_reg_0_ ( .D(N347), .CLK(clk), .RSTB(rst_n), .Q(
        num_of_layer[0]) );
  DFFARX1 disable_neural_reg ( .D(end_neural), .CLK(clk), .RSTB(rst_n), .Q(
        disable_neural) );
  DFFARX1 ena_wr_output_mem_w1_reg ( .D(ena_wr_output_mem), .CLK(clk), .RSTB(
        rst_n), .QN(n2) );
  DFFASX1 ena_wr_output_mem_w2_reg ( .D(n2), .CLK(clk), .SETB(rst_n), .Q(n3)
         );
  DFFASX1 wr_ena_out_n_reg ( .D(n3), .CLK(clk), .SETB(rst_n), .QN(
        wr_ena_out_n_BAR) );
  DFFARX1 ena_wr_int_mem_w1_reg ( .D(n13), .CLK(clk), .RSTB(rst_n), .QN(n1) );
  DFFASX1 ena_wr_int_mem_w2_reg ( .D(n1), .CLK(clk), .SETB(rst_n), .Q(n4) );
  DFFASX1 wr_ena_int_n_reg ( .D(n4), .CLK(clk), .SETB(rst_n), .QN(
        wr_ena_int_n_BAR) );
  DFFARX1 output_mem_addr_reg_0_ ( .D(output_mem_addr_w1[0]), .CLK(clk), 
        .RSTB(rst_n), .Q(output_mem_addr[0]) );
  DFFARX1 output_mem_addr_reg_1_ ( .D(output_mem_addr_w1[1]), .CLK(clk), 
        .RSTB(rst_n), .Q(output_mem_addr[1]) );
  DFFARX1 output_mem_addr_reg_2_ ( .D(output_mem_addr_w1[2]), .CLK(clk), 
        .RSTB(rst_n), .Q(output_mem_addr[2]) );
  DFFARX1 output_mem_addr_reg_3_ ( .D(output_mem_addr_w1[3]), .CLK(clk), 
        .RSTB(rst_n), .Q(output_mem_addr[3]) );
  DFFARX1 output_mem_addr_reg_4_ ( .D(output_mem_addr_w1[4]), .CLK(clk), 
        .RSTB(rst_n), .Q(output_mem_addr[4]) );
  DFFARX1 output_mem_addr_reg_5_ ( .D(output_mem_addr_w1[5]), .CLK(clk), 
        .RSTB(rst_n), .Q(output_mem_addr[5]) );
  DFFARX1 output_mem_addr_reg_6_ ( .D(output_mem_addr_w1[6]), .CLK(clk), 
        .RSTB(rst_n), .Q(output_mem_addr[6]) );
  DFFARX1 output_mem_addr_reg_7_ ( .D(output_mem_addr_w1[7]), .CLK(clk), 
        .RSTB(rst_n), .Q(output_mem_addr[7]) );
  DFFARX1 output_mem_addr_reg_8_ ( .D(output_mem_addr_w1[8]), .CLK(clk), 
        .RSTB(rst_n), .Q(output_mem_addr[8]) );
  DFFARX1 output_mem_addr_reg_9_ ( .D(output_mem_addr_w1[9]), .CLK(clk), 
        .RSTB(rst_n), .Q(output_mem_addr[9]) );
  DFFARX1 int_mem_addr_wr_reg_0_ ( .D(int_mem_addr_wr_w1[0]), .CLK(clk), 
        .RSTB(rst_n), .Q(int_mem_addr_wr[0]) );
  DFFARX1 int_mem_addr_wr_reg_1_ ( .D(int_mem_addr_wr_w1[1]), .CLK(clk), 
        .RSTB(rst_n), .Q(int_mem_addr_wr[1]) );
  DFFARX1 int_mem_addr_wr_reg_2_ ( .D(int_mem_addr_wr_w1[2]), .CLK(clk), 
        .RSTB(rst_n), .Q(int_mem_addr_wr[2]) );
  DFFARX1 int_mem_addr_wr_reg_3_ ( .D(int_mem_addr_wr_w1[3]), .CLK(clk), 
        .RSTB(rst_n), .Q(int_mem_addr_wr[3]) );
  DFFARX1 int_mem_addr_wr_reg_4_ ( .D(int_mem_addr_wr_w1[4]), .CLK(clk), 
        .RSTB(rst_n), .Q(int_mem_addr_wr[4]) );
  DFFARX1 int_mem_addr_wr_reg_5_ ( .D(int_mem_addr_wr_w1[5]), .CLK(clk), 
        .RSTB(rst_n), .Q(int_mem_addr_wr[5]) );
  DFFARX1 int_mem_addr_wr_reg_6_ ( .D(int_mem_addr_wr_w1[6]), .CLK(clk), 
        .RSTB(rst_n), .Q(int_mem_addr_wr[6]) );
  DFFARX1 int_mem_addr_wr_reg_7_ ( .D(int_mem_addr_wr_w1[7]), .CLK(clk), 
        .RSTB(rst_n), .Q(int_mem_addr_wr[7]) );
  DFFARX1 int_mem_addr_wr_reg_8_ ( .D(int_mem_addr_wr_w1[8]), .CLK(clk), 
        .RSTB(rst_n), .Q(int_mem_addr_wr[8]) );
  DFFARX1 int_mem_addr_wr_reg_9_ ( .D(int_mem_addr_wr_w1[9]), .CLK(clk), 
        .RSTB(rst_n), .Q(int_mem_addr_wr[9]) );
  DFFARX1 input_mem_addr_reg_0_ ( .D(input_or_int_mem_addr[0]), .CLK(clk), 
        .RSTB(rst_n), .Q(input_mem_addr[0]) );
  DFFARX1 input_mem_addr_reg_1_ ( .D(input_or_int_mem_addr[1]), .CLK(clk), 
        .RSTB(rst_n), .Q(input_mem_addr[1]) );
  DFFARX1 input_mem_addr_reg_2_ ( .D(input_or_int_mem_addr[2]), .CLK(clk), 
        .RSTB(rst_n), .Q(input_mem_addr[2]) );
  DFFARX1 input_mem_addr_reg_3_ ( .D(input_or_int_mem_addr[3]), .CLK(clk), 
        .RSTB(rst_n), .Q(input_mem_addr[3]) );
  DFFARX1 input_mem_addr_reg_4_ ( .D(input_or_int_mem_addr[4]), .CLK(clk), 
        .RSTB(rst_n), .Q(input_mem_addr[4]) );
  DFFARX1 input_mem_addr_reg_5_ ( .D(input_or_int_mem_addr[5]), .CLK(clk), 
        .RSTB(rst_n), .Q(input_mem_addr[5]) );
  DFFARX1 input_mem_addr_reg_6_ ( .D(input_or_int_mem_addr[6]), .CLK(clk), 
        .RSTB(rst_n), .Q(input_mem_addr[6]) );
  DFFARX1 input_mem_addr_reg_7_ ( .D(input_or_int_mem_addr[7]), .CLK(clk), 
        .RSTB(rst_n), .Q(input_mem_addr[7]) );
  DFFARX1 input_mem_addr_reg_8_ ( .D(input_or_int_mem_addr[8]), .CLK(clk), 
        .RSTB(rst_n), .Q(input_mem_addr[8]) );
  DFFARX1 input_mem_addr_reg_9_ ( .D(input_or_int_mem_addr[9]), .CLK(clk), 
        .RSTB(rst_n), .Q(input_mem_addr[9]) );
  DFFARX1 w_addr_reg_0_ ( .D(w_addr_w1[0]), .CLK(clk), .RSTB(rst_n), .Q(
        w_addr[0]) );
  DFFARX1 w_addr_reg_1_ ( .D(w_addr_w1[1]), .CLK(clk), .RSTB(rst_n), .Q(
        w_addr[1]) );
  DFFARX1 w_addr_reg_2_ ( .D(w_addr_w1[2]), .CLK(clk), .RSTB(rst_n), .Q(
        w_addr[2]) );
  DFFARX1 w_addr_reg_3_ ( .D(w_addr_w1[3]), .CLK(clk), .RSTB(rst_n), .Q(
        w_addr[3]) );
  DFFARX1 w_addr_reg_4_ ( .D(w_addr_w1[4]), .CLK(clk), .RSTB(rst_n), .Q(
        w_addr[4]) );
  DFFARX1 w_addr_reg_5_ ( .D(w_addr_w1[5]), .CLK(clk), .RSTB(rst_n), .Q(
        w_addr[5]) );
  DFFARX1 w_addr_reg_6_ ( .D(w_addr_w1[6]), .CLK(clk), .RSTB(rst_n), .Q(
        w_addr[6]) );
  DFFARX1 w_addr_reg_7_ ( .D(w_addr_w1[7]), .CLK(clk), .RSTB(rst_n), .Q(
        w_addr[7]) );
  DFFARX1 w_addr_reg_8_ ( .D(w_addr_w1[8]), .CLK(clk), .RSTB(rst_n), .Q(
        w_addr[8]) );
  DFFARX1 w_addr_reg_9_ ( .D(w_addr_w1[9]), .CLK(clk), .RSTB(rst_n), .Q(
        w_addr[9]) );
  DFFARX1 w_addr_reg_10_ ( .D(w_addr_w1[10]), .CLK(clk), .RSTB(rst_n), .Q(
        w_addr[10]) );
  DFFARX1 w_addr_reg_11_ ( .D(w_addr_w1[11]), .CLK(clk), .RSTB(rst_n), .Q(
        w_addr[11]) );
  DFFARX1 w_addr_reg_12_ ( .D(w_addr_w1[12]), .CLK(clk), .RSTB(rst_n), .Q(
        w_addr[12]) );
  DFFARX1 w_addr_reg_13_ ( .D(w_addr_w1[13]), .CLK(clk), .RSTB(rst_n), .Q(
        w_addr[13]) );
  DFFARX1 w_addr_reg_14_ ( .D(w_addr_w1[14]), .CLK(clk), .RSTB(rst_n), .Q(
        w_addr[14]) );
  DFFARX1 w_addr_reg_15_ ( .D(w_addr_w1[15]), .CLK(clk), .RSTB(rst_n), .Q(
        w_addr[15]) );
  DFFARX1 w_addr_reg_16_ ( .D(w_addr_w1[16]), .CLK(clk), .RSTB(rst_n), .Q(
        w_addr[16]) );
  DFFARX1 w_addr_reg_17_ ( .D(w_addr_w1[17]), .CLK(clk), .RSTB(rst_n), .Q(
        w_addr[17]) );
  DFFARX1 w_addr_reg_18_ ( .D(w_addr_w1[18]), .CLK(clk), .RSTB(rst_n), .Q(
        w_addr[18]) );
  DFFARX1 w_addr_reg_19_ ( .D(w_addr_w1[19]), .CLK(clk), .RSTB(rst_n), .Q(
        w_addr[19]) );
  DFFARX1 mac_input_01_reg_8_ ( .D(N99), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_01[8]) );
  DFFARX1 mac_input_01_reg_7_ ( .D(N98), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_01[7]) );
  DFFARX1 mac_input_01_reg_6_ ( .D(N97), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_01[6]) );
  DFFARX1 mac_input_01_reg_5_ ( .D(N96), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_01[5]) );
  DFFARX1 mac_input_01_reg_4_ ( .D(N95), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_01[4]) );
  DFFARX1 mac_input_01_reg_3_ ( .D(N94), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_01[3]) );
  DFFARX1 mac_input_01_reg_2_ ( .D(N93), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_01[2]) );
  DFFARX1 mac_input_01_reg_1_ ( .D(N92), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_01[1]) );
  DFFARX1 mac_input_01_reg_0_ ( .D(N91), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_01[0]) );
  DFFARX1 mac_input_01_reg_31_ ( .D(N122), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_01[31]) );
  DFFARX1 mac_input_01_reg_30_ ( .D(N121), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_01[30]) );
  DFFARX1 mac_input_01_reg_29_ ( .D(N120), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_01[29]) );
  DFFARX1 mac_input_01_reg_28_ ( .D(N119), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_01[28]) );
  DFFARX1 mac_input_01_reg_27_ ( .D(N118), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_01[27]) );
  DFFARX1 mac_input_01_reg_26_ ( .D(N117), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_01[26]) );
  DFFARX1 mac_input_01_reg_25_ ( .D(N116), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_01[25]) );
  DFFARX1 mac_input_01_reg_24_ ( .D(N115), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_01[24]) );
  DFFARX1 mac_input_01_reg_23_ ( .D(N114), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_01[23]) );
  DFFARX1 mac_input_01_reg_22_ ( .D(N113), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_01[22]) );
  DFFARX1 mac_input_01_reg_21_ ( .D(N112), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_01[21]) );
  DFFARX1 mac_input_01_reg_20_ ( .D(N111), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_01[20]) );
  DFFARX1 mac_input_01_reg_19_ ( .D(N110), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_01[19]) );
  DFFARX1 mac_input_01_reg_18_ ( .D(N109), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_01[18]) );
  DFFARX1 mac_input_01_reg_17_ ( .D(N108), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_01[17]) );
  DFFARX1 mac_input_01_reg_16_ ( .D(N107), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_01[16]) );
  DFFARX1 mac_input_01_reg_15_ ( .D(N106), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_01[15]) );
  DFFARX1 mac_input_01_reg_14_ ( .D(N105), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_01[14]) );
  DFFARX1 mac_input_01_reg_13_ ( .D(N104), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_01[13]) );
  DFFARX1 mac_input_01_reg_12_ ( .D(N103), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_01[12]) );
  DFFARX1 mac_input_01_reg_11_ ( .D(N102), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_01[11]) );
  DFFARX1 mac_input_01_reg_10_ ( .D(N101), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_01[10]) );
  DFFARX1 mac_input_01_reg_9_ ( .D(N100), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_01[9]) );
  DFFARX1 mac_input_02_reg_0_ ( .D(N126), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_02[0]) );
  DFFARX1 mac_input_02_reg_1_ ( .D(N127), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_02[1]) );
  DFFARX1 mac_input_02_reg_2_ ( .D(N128), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_02[2]) );
  DFFARX1 mac_input_02_reg_3_ ( .D(N129), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_02[3]) );
  DFFARX1 mac_input_02_reg_4_ ( .D(N130), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_02[4]) );
  DFFARX1 mac_input_02_reg_5_ ( .D(N131), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_02[5]) );
  DFFARX1 mac_input_02_reg_6_ ( .D(N132), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_02[6]) );
  DFFARX1 mac_input_02_reg_7_ ( .D(N133), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_02[7]) );
  DFFARX1 mac_input_02_reg_8_ ( .D(N134), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_02[8]) );
  DFFARX1 mac_input_02_reg_9_ ( .D(N135), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_02[9]) );
  DFFARX1 mac_input_02_reg_10_ ( .D(N136), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_02[10]) );
  DFFARX1 mac_input_02_reg_11_ ( .D(N137), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_02[11]) );
  DFFARX1 mac_input_02_reg_12_ ( .D(N138), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_02[12]) );
  DFFARX1 mac_input_02_reg_13_ ( .D(N139), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_02[13]) );
  DFFARX1 mac_input_02_reg_14_ ( .D(N140), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_02[14]) );
  DFFARX1 mac_input_02_reg_15_ ( .D(N141), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_02[15]) );
  DFFARX1 mac_input_02_reg_16_ ( .D(N142), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_02[16]) );
  DFFARX1 mac_input_02_reg_17_ ( .D(N143), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_02[17]) );
  DFFARX1 mac_input_02_reg_18_ ( .D(N144), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_02[18]) );
  DFFARX1 mac_input_02_reg_19_ ( .D(N145), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_02[19]) );
  DFFARX1 mac_input_02_reg_20_ ( .D(N146), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_02[20]) );
  DFFARX1 mac_input_02_reg_21_ ( .D(N147), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_02[21]) );
  DFFARX1 mac_input_02_reg_22_ ( .D(N148), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_02[22]) );
  DFFARX1 mac_input_02_reg_23_ ( .D(N149), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_02[23]) );
  DFFARX1 mac_input_02_reg_24_ ( .D(N150), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_02[24]) );
  DFFARX1 mac_input_02_reg_25_ ( .D(N151), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_02[25]) );
  DFFARX1 mac_input_02_reg_26_ ( .D(N152), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_02[26]) );
  DFFARX1 mac_input_02_reg_27_ ( .D(N153), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_02[27]) );
  DFFARX1 mac_input_02_reg_28_ ( .D(N154), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_02[28]) );
  DFFARX1 mac_input_02_reg_29_ ( .D(N155), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_02[29]) );
  DFFARX1 mac_input_02_reg_30_ ( .D(N156), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_02[30]) );
  DFFARX1 mac_input_02_reg_31_ ( .D(N157), .CLK(clk), .RSTB(rst_n), .Q(
        mac_input_02[31]) );
  DFFARX1 input_act_func_reg_0_ ( .D(N160), .CLK(clk), .RSTB(rst_n), .Q(
        input_act_func[0]) );
  DFFARX1 input_act_func_reg_1_ ( .D(N161), .CLK(clk), .RSTB(rst_n), .Q(
        input_act_func[1]) );
  DFFARX1 input_act_func_reg_2_ ( .D(N162), .CLK(clk), .RSTB(rst_n), .Q(
        input_act_func[2]) );
  DFFARX1 input_act_func_reg_4_ ( .D(N164), .CLK(clk), .RSTB(rst_n), .Q(
        input_act_func[4]) );
  DFFARX1 input_act_func_reg_6_ ( .D(N166), .CLK(clk), .RSTB(rst_n), .Q(
        input_act_func[6]) );
  DFFARX1 input_act_func_reg_7_ ( .D(N167), .CLK(clk), .RSTB(rst_n), .Q(
        input_act_func[7]) );
  DFFARX1 input_act_func_reg_8_ ( .D(N168), .CLK(clk), .RSTB(rst_n), .Q(
        input_act_func[8]) );
  DFFARX1 input_act_func_reg_10_ ( .D(N170), .CLK(clk), .RSTB(rst_n), .Q(
        input_act_func[10]) );
  DFFARX1 input_act_func_reg_12_ ( .D(N172), .CLK(clk), .RSTB(rst_n), .Q(
        input_act_func[12]) );
  DFFARX1 input_act_func_reg_14_ ( .D(N174), .CLK(clk), .RSTB(rst_n), .Q(
        input_act_func[14]) );
  DFFARX1 input_act_func_reg_16_ ( .D(N176), .CLK(clk), .RSTB(rst_n), .Q(
        input_act_func[16]) );
  DFFARX1 input_act_func_reg_18_ ( .D(N178), .CLK(clk), .RSTB(rst_n), .Q(
        input_act_func[18]) );
  DFFARX1 input_act_func_reg_20_ ( .D(N180), .CLK(clk), .RSTB(rst_n), .Q(
        input_act_func[20]) );
  DFFARX1 input_act_func_reg_21_ ( .D(N181), .CLK(clk), .RSTB(rst_n), .Q(
        input_act_func[21]) );
  DFFARX1 input_act_func_reg_22_ ( .D(N182), .CLK(clk), .RSTB(rst_n), .Q(
        input_act_func[22]) );
  DFFARX1 input_act_func_reg_23_ ( .D(N183), .CLK(clk), .RSTB(rst_n), .Q(
        input_act_func[23]) );
  DFFARX1 input_act_func_reg_24_ ( .D(N184), .CLK(clk), .RSTB(rst_n), .Q(
        input_act_func[24]) );
  DFFARX1 input_act_func_reg_25_ ( .D(N185), .CLK(clk), .RSTB(rst_n), .Q(
        input_act_func[25]) );
  DFFARX1 input_act_func_reg_26_ ( .D(N186), .CLK(clk), .RSTB(rst_n), .Q(
        input_act_func[26]) );
  DFFARX1 input_act_func_reg_27_ ( .D(N187), .CLK(clk), .RSTB(rst_n), .Q(
        input_act_func[27]) );
  DFFARX1 input_act_func_reg_28_ ( .D(N188), .CLK(clk), .RSTB(rst_n), .Q(
        input_act_func[28]) );
  DFFARX1 input_act_func_reg_29_ ( .D(N189), .CLK(clk), .RSTB(rst_n), .Q(
        input_act_func[29]) );
  DFFARX1 input_act_func_reg_30_ ( .D(N190), .CLK(clk), .RSTB(rst_n), .Q(
        input_act_func[30]) );
  DFFARX1 input_act_func_reg_31_ ( .D(N191), .CLK(clk), .RSTB(rst_n), .Q(
        input_act_func[31]) );
  DFFARX1 mac_time_reg_11_ ( .D(N362), .CLK(clk), .RSTB(rst_n), .Q(
        mac_time[11]) );
  DFFARX1 mac_time_reg_10_ ( .D(N361), .CLK(clk), .RSTB(rst_n), .Q(
        mac_time[10]) );
  DFFARX1 mac_time_reg_9_ ( .D(N360), .CLK(clk), .RSTB(rst_n), .Q(mac_time[9])
         );
  DFFARX1 mac_time_reg_8_ ( .D(N359), .CLK(clk), .RSTB(rst_n), .Q(mac_time[8])
         );
  DFFARX1 mac_time_reg_7_ ( .D(N358), .CLK(clk), .RSTB(rst_n), .Q(mac_time[7])
         );
  DFFARX1 mac_time_reg_6_ ( .D(N357), .CLK(clk), .RSTB(rst_n), .Q(mac_time[6])
         );
  DFFARX1 mac_time_reg_5_ ( .D(N356), .CLK(clk), .RSTB(rst_n), .Q(mac_time[5])
         );
  DFFARX1 mac_time_reg_4_ ( .D(N355), .CLK(clk), .RSTB(rst_n), .Q(mac_time[4])
         );
  DFFARX1 mac_time_reg_3_ ( .D(N354), .CLK(clk), .RSTB(rst_n), .Q(mac_time[3])
         );
  DFFARX1 mac_time_reg_2_ ( .D(N353), .CLK(clk), .RSTB(rst_n), .Q(mac_time[2])
         );
  DFFARX1 mac_time_reg_1_ ( .D(N352), .CLK(clk), .RSTB(rst_n), .Q(mac_time[1])
         );
  DFFARX1 mac_time_reg_0_ ( .D(N351), .CLK(clk), .RSTB(rst_n), .Q(mac_time[0])
         );
  DFFARX1 num_of_layer_reg_3_ ( .D(N350), .CLK(clk), .RSTB(rst_n), .Q(
        num_of_layer[3]) );
  DFFARX1 num_of_layer_reg_2_ ( .D(N349), .CLK(clk), .RSTB(rst_n), .Q(
        num_of_layer[2]) );
  DFFARX1 num_of_layer_reg_1_ ( .D(N348), .CLK(clk), .RSTB(rst_n), .Q(
        num_of_layer[1]) );
  DFFARX1 num_of_node_for_each_layer_reg_7_ ( .D(N370), .CLK(clk), .RSTB(rst_n), .Q(num_of_node_for_each_layer[7]) );
  DFFARX1 num_of_node_for_each_layer_reg_6_ ( .D(N369), .CLK(clk), .RSTB(rst_n), .Q(num_of_node_for_each_layer[6]) );
  DFFARX1 num_of_node_for_each_layer_reg_5_ ( .D(N368), .CLK(clk), .RSTB(rst_n), .Q(num_of_node_for_each_layer[5]) );
  DFFARX1 num_of_node_for_each_layer_reg_4_ ( .D(N367), .CLK(clk), .RSTB(rst_n), .Q(num_of_node_for_each_layer[4]) );
  DFFARX1 num_of_node_for_each_layer_reg_3_ ( .D(N366), .CLK(clk), .RSTB(rst_n), .Q(num_of_node_for_each_layer[3]) );
  DFFARX1 num_of_node_for_each_layer_reg_2_ ( .D(N365), .CLK(clk), .RSTB(rst_n), .Q(num_of_node_for_each_layer[2]) );
  DFFARX1 num_of_node_for_each_layer_reg_1_ ( .D(N364), .CLK(clk), .RSTB(rst_n), .Q(num_of_node_for_each_layer[1]) );
  DFFARX1 num_of_node_for_each_layer_reg_0_ ( .D(N363), .CLK(clk), .RSTB(rst_n), .Q(num_of_node_for_each_layer[0]) );
  DFFARX1 user_para_addr_reg_0_ ( .D(para_addr[0]), .CLK(clk), .RSTB(rst_n), 
        .Q(user_para_addr[0]) );
  DFFARX1 user_para_addr_reg_1_ ( .D(para_addr[1]), .CLK(clk), .RSTB(rst_n), 
        .Q(user_para_addr[1]) );
  DFFARX1 user_para_addr_reg_2_ ( .D(para_addr[2]), .CLK(clk), .RSTB(rst_n), 
        .Q(user_para_addr[2]) );
  DFFARX1 user_para_addr_reg_3_ ( .D(para_addr[3]), .CLK(clk), .RSTB(rst_n), 
        .Q(user_para_addr[3]) );
  DFFARX1 user_para_addr_reg_4_ ( .D(para_addr[4]), .CLK(clk), .RSTB(rst_n), 
        .Q(user_para_addr[4]) );
  DFFARX1 user_para_addr_reg_5_ ( .D(para_addr[5]), .CLK(clk), .RSTB(rst_n), 
        .Q(user_para_addr[5]) );
  DFFARX1 user_para_addr_reg_6_ ( .D(para_addr[6]), .CLK(clk), .RSTB(rst_n), 
        .Q(user_para_addr[6]) );
  DFFARX1 user_para_addr_reg_7_ ( .D(para_addr[7]), .CLK(clk), .RSTB(rst_n), 
        .Q(user_para_addr[7]) );
  DFFARX1 user_para_addr_reg_8_ ( .D(para_addr[8]), .CLK(clk), .RSTB(rst_n), 
        .Q(user_para_addr[8]) );
  DFFARX1 user_para_addr_reg_9_ ( .D(para_addr[9]), .CLK(clk), .RSTB(rst_n), 
        .Q(user_para_addr[9]) );
  DFFARX1 act_function_sel_reg_1_ ( .D(N372), .CLK(clk), .RSTB(rst_n), .Q(
        act_function_sel[1]) );
  DFFARX1 act_function_sel_reg_0_ ( .D(N371), .CLK(clk), .RSTB(rst_n), .Q(
        act_function_sel[0]), .QN(n8) );
  DFFARX1 out_act_func_reg_31_ ( .D(N266), .CLK(clk), .RSTB(rst_n), .Q(
        out_act_func[31]) );
  DFFARX1 int_mem_data_wr_reg_31_ ( .D(N303), .CLK(clk), .RSTB(rst_n), .Q(
        int_mem_data_wr[31]) );
  DFFARX1 output_data_reg_31_ ( .D(N338), .CLK(clk), .RSTB(rst_n), .Q(
        output_data[31]) );
  DFFARX1 out_act_func_reg_30_ ( .D(N265), .CLK(clk), .RSTB(rst_n), .Q(
        out_act_func[30]) );
  DFFARX1 int_mem_data_wr_reg_30_ ( .D(N302), .CLK(clk), .RSTB(rst_n), .Q(
        int_mem_data_wr[30]) );
  DFFARX1 output_data_reg_30_ ( .D(N337), .CLK(clk), .RSTB(rst_n), .Q(
        output_data[30]) );
  DFFARX1 out_act_func_reg_29_ ( .D(N264), .CLK(clk), .RSTB(rst_n), .Q(
        out_act_func[29]) );
  DFFARX1 int_mem_data_wr_reg_29_ ( .D(N301), .CLK(clk), .RSTB(rst_n), .Q(
        int_mem_data_wr[29]) );
  DFFARX1 output_data_reg_29_ ( .D(N336), .CLK(clk), .RSTB(rst_n), .Q(
        output_data[29]) );
  DFFARX1 out_act_func_reg_28_ ( .D(N263), .CLK(clk), .RSTB(rst_n), .Q(
        out_act_func[28]) );
  DFFARX1 int_mem_data_wr_reg_28_ ( .D(N300), .CLK(clk), .RSTB(rst_n), .Q(
        int_mem_data_wr[28]) );
  DFFARX1 output_data_reg_28_ ( .D(N335), .CLK(clk), .RSTB(rst_n), .Q(
        output_data[28]) );
  DFFARX1 out_act_func_reg_27_ ( .D(N262), .CLK(clk), .RSTB(rst_n), .Q(
        out_act_func[27]) );
  DFFARX1 int_mem_data_wr_reg_27_ ( .D(N299), .CLK(clk), .RSTB(rst_n), .Q(
        int_mem_data_wr[27]) );
  DFFARX1 output_data_reg_27_ ( .D(N334), .CLK(clk), .RSTB(rst_n), .Q(
        output_data[27]) );
  DFFARX1 out_act_func_reg_26_ ( .D(N261), .CLK(clk), .RSTB(rst_n), .Q(
        out_act_func[26]) );
  DFFARX1 int_mem_data_wr_reg_26_ ( .D(N298), .CLK(clk), .RSTB(rst_n), .Q(
        int_mem_data_wr[26]) );
  DFFARX1 output_data_reg_26_ ( .D(N333), .CLK(clk), .RSTB(rst_n), .Q(
        output_data[26]) );
  DFFARX1 out_act_func_reg_25_ ( .D(N260), .CLK(clk), .RSTB(rst_n), .Q(
        out_act_func[25]) );
  DFFARX1 int_mem_data_wr_reg_25_ ( .D(N297), .CLK(clk), .RSTB(rst_n), .Q(
        int_mem_data_wr[25]) );
  DFFARX1 output_data_reg_25_ ( .D(N332), .CLK(clk), .RSTB(rst_n), .Q(
        output_data[25]) );
  DFFARX1 out_act_func_reg_24_ ( .D(N259), .CLK(clk), .RSTB(rst_n), .Q(
        out_act_func[24]) );
  DFFARX1 int_mem_data_wr_reg_24_ ( .D(N296), .CLK(clk), .RSTB(rst_n), .Q(
        int_mem_data_wr[24]) );
  DFFARX1 output_data_reg_24_ ( .D(N331), .CLK(clk), .RSTB(rst_n), .Q(
        output_data[24]) );
  DFFARX1 out_act_func_reg_23_ ( .D(N258), .CLK(clk), .RSTB(rst_n), .Q(
        out_act_func[23]) );
  DFFARX1 int_mem_data_wr_reg_23_ ( .D(N295), .CLK(clk), .RSTB(rst_n), .Q(
        int_mem_data_wr[23]) );
  DFFARX1 output_data_reg_23_ ( .D(N330), .CLK(clk), .RSTB(rst_n), .Q(
        output_data[23]) );
  DFFARX1 out_act_func_reg_22_ ( .D(N257), .CLK(clk), .RSTB(rst_n), .Q(
        out_act_func[22]) );
  DFFARX1 int_mem_data_wr_reg_22_ ( .D(N294), .CLK(clk), .RSTB(rst_n), .Q(
        int_mem_data_wr[22]) );
  DFFARX1 output_data_reg_22_ ( .D(N329), .CLK(clk), .RSTB(rst_n), .Q(
        output_data[22]) );
  DFFARX1 out_act_func_reg_21_ ( .D(N256), .CLK(clk), .RSTB(rst_n), .Q(
        out_act_func[21]) );
  DFFARX1 int_mem_data_wr_reg_21_ ( .D(N293), .CLK(clk), .RSTB(rst_n), .Q(
        int_mem_data_wr[21]) );
  DFFARX1 output_data_reg_21_ ( .D(N328), .CLK(clk), .RSTB(rst_n), .Q(
        output_data[21]) );
  DFFARX1 out_act_func_reg_20_ ( .D(N255), .CLK(clk), .RSTB(rst_n), .Q(
        out_act_func[20]) );
  DFFARX1 int_mem_data_wr_reg_20_ ( .D(N292), .CLK(clk), .RSTB(rst_n), .Q(
        int_mem_data_wr[20]) );
  DFFARX1 output_data_reg_20_ ( .D(N327), .CLK(clk), .RSTB(rst_n), .Q(
        output_data[20]) );
  DFFARX1 out_act_func_reg_19_ ( .D(N254), .CLK(clk), .RSTB(rst_n), .Q(
        out_act_func[19]) );
  DFFARX1 int_mem_data_wr_reg_19_ ( .D(N291), .CLK(clk), .RSTB(rst_n), .Q(
        int_mem_data_wr[19]) );
  DFFARX1 output_data_reg_19_ ( .D(N326), .CLK(clk), .RSTB(rst_n), .Q(
        output_data[19]) );
  DFFARX1 out_act_func_reg_18_ ( .D(N253), .CLK(clk), .RSTB(rst_n), .Q(
        out_act_func[18]) );
  DFFARX1 int_mem_data_wr_reg_18_ ( .D(N290), .CLK(clk), .RSTB(rst_n), .Q(
        int_mem_data_wr[18]) );
  DFFARX1 output_data_reg_18_ ( .D(N325), .CLK(clk), .RSTB(rst_n), .Q(
        output_data[18]) );
  DFFARX1 out_act_func_reg_17_ ( .D(N252), .CLK(clk), .RSTB(rst_n), .Q(
        out_act_func[17]) );
  DFFARX1 int_mem_data_wr_reg_17_ ( .D(N289), .CLK(clk), .RSTB(rst_n), .Q(
        int_mem_data_wr[17]) );
  DFFARX1 output_data_reg_17_ ( .D(N324), .CLK(clk), .RSTB(rst_n), .Q(
        output_data[17]) );
  DFFARX1 out_act_func_reg_16_ ( .D(N251), .CLK(clk), .RSTB(rst_n), .Q(
        out_act_func[16]) );
  DFFARX1 int_mem_data_wr_reg_16_ ( .D(N288), .CLK(clk), .RSTB(rst_n), .Q(
        int_mem_data_wr[16]) );
  DFFARX1 output_data_reg_16_ ( .D(N323), .CLK(clk), .RSTB(rst_n), .Q(
        output_data[16]) );
  DFFARX1 out_act_func_reg_15_ ( .D(N250), .CLK(clk), .RSTB(rst_n), .Q(
        out_act_func[15]) );
  DFFARX1 int_mem_data_wr_reg_15_ ( .D(N287), .CLK(clk), .RSTB(rst_n), .Q(
        int_mem_data_wr[15]) );
  DFFARX1 output_data_reg_15_ ( .D(N322), .CLK(clk), .RSTB(rst_n), .Q(
        output_data[15]) );
  DFFARX1 out_act_func_reg_14_ ( .D(N249), .CLK(clk), .RSTB(rst_n), .Q(
        out_act_func[14]) );
  DFFARX1 int_mem_data_wr_reg_14_ ( .D(N286), .CLK(clk), .RSTB(rst_n), .Q(
        int_mem_data_wr[14]) );
  DFFARX1 output_data_reg_14_ ( .D(N321), .CLK(clk), .RSTB(rst_n), .Q(
        output_data[14]) );
  DFFARX1 out_act_func_reg_13_ ( .D(N248), .CLK(clk), .RSTB(rst_n), .Q(
        out_act_func[13]) );
  DFFARX1 int_mem_data_wr_reg_13_ ( .D(N285), .CLK(clk), .RSTB(rst_n), .Q(
        int_mem_data_wr[13]) );
  DFFARX1 output_data_reg_13_ ( .D(N320), .CLK(clk), .RSTB(rst_n), .Q(
        output_data[13]) );
  DFFARX1 out_act_func_reg_12_ ( .D(N247), .CLK(clk), .RSTB(rst_n), .Q(
        out_act_func[12]) );
  DFFARX1 int_mem_data_wr_reg_12_ ( .D(N284), .CLK(clk), .RSTB(rst_n), .Q(
        int_mem_data_wr[12]) );
  DFFARX1 output_data_reg_12_ ( .D(N319), .CLK(clk), .RSTB(rst_n), .Q(
        output_data[12]) );
  DFFARX1 out_act_func_reg_11_ ( .D(N246), .CLK(clk), .RSTB(rst_n), .Q(
        out_act_func[11]) );
  DFFARX1 int_mem_data_wr_reg_11_ ( .D(N283), .CLK(clk), .RSTB(rst_n), .Q(
        int_mem_data_wr[11]) );
  DFFARX1 output_data_reg_11_ ( .D(N318), .CLK(clk), .RSTB(rst_n), .Q(
        output_data[11]) );
  DFFARX1 out_act_func_reg_10_ ( .D(N245), .CLK(clk), .RSTB(rst_n), .Q(
        out_act_func[10]) );
  DFFARX1 int_mem_data_wr_reg_10_ ( .D(N282), .CLK(clk), .RSTB(rst_n), .Q(
        int_mem_data_wr[10]) );
  DFFARX1 output_data_reg_10_ ( .D(N317), .CLK(clk), .RSTB(rst_n), .Q(
        output_data[10]) );
  DFFARX1 out_act_func_reg_9_ ( .D(N244), .CLK(clk), .RSTB(rst_n), .Q(
        out_act_func[9]) );
  DFFARX1 int_mem_data_wr_reg_9_ ( .D(N281), .CLK(clk), .RSTB(rst_n), .Q(
        int_mem_data_wr[9]) );
  DFFARX1 output_data_reg_9_ ( .D(N316), .CLK(clk), .RSTB(rst_n), .Q(
        output_data[9]) );
  DFFARX1 out_act_func_reg_8_ ( .D(N243), .CLK(clk), .RSTB(rst_n), .Q(
        out_act_func[8]) );
  DFFARX1 int_mem_data_wr_reg_8_ ( .D(N280), .CLK(clk), .RSTB(rst_n), .Q(
        int_mem_data_wr[8]) );
  DFFARX1 output_data_reg_8_ ( .D(N315), .CLK(clk), .RSTB(rst_n), .Q(
        output_data[8]) );
  DFFARX1 out_act_func_reg_7_ ( .D(N242), .CLK(clk), .RSTB(rst_n), .Q(
        out_act_func[7]) );
  DFFARX1 int_mem_data_wr_reg_7_ ( .D(N279), .CLK(clk), .RSTB(rst_n), .Q(
        int_mem_data_wr[7]) );
  DFFARX1 output_data_reg_7_ ( .D(N314), .CLK(clk), .RSTB(rst_n), .Q(
        output_data[7]) );
  DFFARX1 out_act_func_reg_6_ ( .D(N241), .CLK(clk), .RSTB(rst_n), .Q(
        out_act_func[6]) );
  DFFARX1 int_mem_data_wr_reg_6_ ( .D(N278), .CLK(clk), .RSTB(rst_n), .Q(
        int_mem_data_wr[6]) );
  DFFARX1 output_data_reg_6_ ( .D(N313), .CLK(clk), .RSTB(rst_n), .Q(
        output_data[6]) );
  DFFARX1 out_act_func_reg_5_ ( .D(N240), .CLK(clk), .RSTB(rst_n), .Q(
        out_act_func[5]) );
  DFFARX1 int_mem_data_wr_reg_5_ ( .D(N277), .CLK(clk), .RSTB(rst_n), .Q(
        int_mem_data_wr[5]) );
  DFFARX1 output_data_reg_5_ ( .D(N312), .CLK(clk), .RSTB(rst_n), .Q(
        output_data[5]) );
  DFFARX1 out_act_func_reg_4_ ( .D(N239), .CLK(clk), .RSTB(rst_n), .Q(
        out_act_func[4]) );
  DFFARX1 int_mem_data_wr_reg_4_ ( .D(N276), .CLK(clk), .RSTB(rst_n), .Q(
        int_mem_data_wr[4]) );
  DFFARX1 output_data_reg_4_ ( .D(N311), .CLK(clk), .RSTB(rst_n), .Q(
        output_data[4]) );
  DFFARX1 out_act_func_reg_3_ ( .D(N238), .CLK(clk), .RSTB(rst_n), .Q(
        out_act_func[3]) );
  DFFARX1 int_mem_data_wr_reg_3_ ( .D(N275), .CLK(clk), .RSTB(rst_n), .Q(
        int_mem_data_wr[3]) );
  DFFARX1 output_data_reg_3_ ( .D(N310), .CLK(clk), .RSTB(rst_n), .Q(
        output_data[3]) );
  DFFARX1 out_act_func_reg_2_ ( .D(N237), .CLK(clk), .RSTB(rst_n), .Q(
        out_act_func[2]) );
  DFFARX1 int_mem_data_wr_reg_2_ ( .D(N274), .CLK(clk), .RSTB(rst_n), .Q(
        int_mem_data_wr[2]) );
  DFFARX1 output_data_reg_2_ ( .D(N309), .CLK(clk), .RSTB(rst_n), .Q(
        output_data[2]) );
  DFFARX1 out_act_func_reg_1_ ( .D(N236), .CLK(clk), .RSTB(rst_n), .Q(
        out_act_func[1]) );
  DFFARX1 int_mem_data_wr_reg_1_ ( .D(N273), .CLK(clk), .RSTB(rst_n), .Q(
        int_mem_data_wr[1]) );
  DFFARX1 output_data_reg_1_ ( .D(N308), .CLK(clk), .RSTB(rst_n), .Q(
        output_data[1]) );
  DFFARX1 out_act_func_reg_0_ ( .D(N235), .CLK(clk), .RSTB(rst_n), .Q(
        out_act_func[0]) );
  DFFARX1 int_mem_data_wr_reg_0_ ( .D(N272), .CLK(clk), .RSTB(rst_n), .Q(
        int_mem_data_wr[0]) );
  DFFARX1 output_data_reg_0_ ( .D(N307), .CLK(clk), .RSTB(rst_n), .Q(
        output_data[0]) );
  DFFARX1 input_act_func_reg_9_ ( .D(N169), .CLK(clk), .RSTB(rst_n), .Q(
        input_act_func[9]) );
  DFFARX1 input_act_func_reg_5_ ( .D(N165), .CLK(clk), .RSTB(rst_n), .Q(
        input_act_func[5]) );
  DFFARX1 input_act_func_reg_3_ ( .D(N163), .CLK(clk), .RSTB(rst_n), .Q(
        input_act_func[3]) );
  DFFARX1 input_act_func_reg_11_ ( .D(N171), .CLK(clk), .RSTB(rst_n), .Q(
        input_act_func[11]) );
  DFFARX1 input_act_func_reg_13_ ( .D(N173), .CLK(clk), .RSTB(rst_n), .Q(
        input_act_func[13]) );
  DFFARX1 input_act_func_reg_17_ ( .D(N177), .CLK(clk), .RSTB(rst_n), .Q(
        input_act_func[17]) );
  DFFARX1 input_act_func_reg_15_ ( .D(N175), .CLK(clk), .RSTB(rst_n), .Q(
        input_act_func[15]) );
  DFFARX1 input_act_func_reg_19_ ( .D(N179), .CLK(clk), .RSTB(rst_n), .Q(
        input_act_func[19]) );
  NAND2X0 U3 ( .IN1(n43), .IN2(linear_output[23]), .QN(n20) );
  NAND2X0 U4 ( .IN1(n42), .IN2(tansigmoid_output[23]), .QN(n21) );
  NAND2X0 U5 ( .IN1(n7), .IN2(sigmoid_output[23]), .QN(n22) );
  NAND2X0 U6 ( .IN1(n43), .IN2(linear_output[24]), .QN(n23) );
  NAND2X0 U7 ( .IN1(n42), .IN2(tansigmoid_output[24]), .QN(n24) );
  NAND2X0 U8 ( .IN1(n7), .IN2(sigmoid_output[24]), .QN(n25) );
  NAND2X0 U9 ( .IN1(n43), .IN2(linear_output[25]), .QN(n26) );
  NAND2X0 U10 ( .IN1(n42), .IN2(tansigmoid_output[25]), .QN(n27) );
  NAND2X0 U11 ( .IN1(n7), .IN2(sigmoid_output[25]), .QN(n28) );
  NAND2X0 U12 ( .IN1(n43), .IN2(linear_output[26]), .QN(n29) );
  NAND2X0 U13 ( .IN1(n42), .IN2(tansigmoid_output[26]), .QN(n30) );
  NAND2X0 U14 ( .IN1(n7), .IN2(sigmoid_output[26]), .QN(n31) );
  NAND2X0 U15 ( .IN1(n43), .IN2(linear_output[27]), .QN(n32) );
  NAND2X0 U16 ( .IN1(n42), .IN2(tansigmoid_output[27]), .QN(n33) );
  NAND2X0 U17 ( .IN1(n7), .IN2(sigmoid_output[27]), .QN(n34) );
  NAND2X0 U18 ( .IN1(n43), .IN2(linear_output[28]), .QN(n35) );
  NAND2X0 U19 ( .IN1(n42), .IN2(tansigmoid_output[28]), .QN(n36) );
  NAND2X0 U20 ( .IN1(n7), .IN2(sigmoid_output[28]), .QN(n37) );
  NAND2X0 U21 ( .IN1(n43), .IN2(linear_output[29]), .QN(n38) );
  NAND2X0 U22 ( .IN1(n42), .IN2(tansigmoid_output[29]), .QN(n39) );
  NAND2X0 U23 ( .IN1(n7), .IN2(sigmoid_output[29]), .QN(n40) );
  NAND2X0 U24 ( .IN1(n9), .IN2(n10), .QN(N265) );
  NAND2X0 U25 ( .IN1(n42), .IN2(tansigmoid_output[30]), .QN(n10) );
  NAND2X0 U26 ( .IN1(n7), .IN2(sigmoid_output[30]), .QN(n9) );
  NBUFFX8 U27 ( .INP(ena_act_func), .Z(n14) );
  NBUFFX8 U28 ( .INP(n53), .Z(n13) );
  NBUFFX8 U29 ( .INP(n44), .Z(n12) );
  NAND2X0 U30 ( .IN1(ena_wr_output_mem), .IN2(n13), .QN(n44) );
  INVX0 U31 ( .INP(ena_wr_int_mem), .ZN(n53) );
  NAND3X0 U32 ( .IN1(para_cof[1]), .IN2(n47), .IN3(n50), .QN(n46) );
  NOR2X0 U33 ( .IN1(input_or_int_mem_sel), .IN2(n15), .QN(n6) );
  AND2X1 U34 ( .IN1(n11), .IN2(input_or_int_mem_sel), .Q(n5) );
  AND3X1 U35 ( .IN1(act_function_sel[1]), .IN2(act_function_sel[0]), .IN3(n18), 
        .Q(n42) );
  AND2X1 U36 ( .IN1(act_function_sel[0]), .IN2(n19), .Q(n43) );
  NOR2X0 U37 ( .IN1(act_function_sel[0]), .IN2(n16), .QN(n7) );
  NAND2X0 U38 ( .IN1(act_function_sel[1]), .IN2(n18), .QN(n16) );
  INVX0 U39 ( .INP(n15), .ZN(n11) );
  NOR2X0 U40 ( .IN1(ena_mac_wait), .IN2(ena_mac), .QN(n15) );
  AO22X1 U42 ( .IN1(n5), .IN2(input_mem_data[9]), .IN3(n6), .IN4(
        int_mem_data_rd[9]), .Q(N100) );
  AO22X1 U43 ( .IN1(n5), .IN2(input_mem_data[10]), .IN3(n6), .IN4(
        int_mem_data_rd[10]), .Q(N101) );
  AO22X1 U44 ( .IN1(n5), .IN2(input_mem_data[11]), .IN3(n6), .IN4(
        int_mem_data_rd[11]), .Q(N102) );
  AO22X1 U45 ( .IN1(n5), .IN2(input_mem_data[12]), .IN3(n6), .IN4(
        int_mem_data_rd[12]), .Q(N103) );
  AO22X1 U46 ( .IN1(n5), .IN2(input_mem_data[13]), .IN3(n6), .IN4(
        int_mem_data_rd[13]), .Q(N104) );
  AO22X1 U47 ( .IN1(n5), .IN2(input_mem_data[14]), .IN3(n6), .IN4(
        int_mem_data_rd[14]), .Q(N105) );
  AO22X1 U48 ( .IN1(n5), .IN2(input_mem_data[15]), .IN3(n6), .IN4(
        int_mem_data_rd[15]), .Q(N106) );
  AO22X1 U49 ( .IN1(n5), .IN2(input_mem_data[16]), .IN3(n6), .IN4(
        int_mem_data_rd[16]), .Q(N107) );
  AO22X1 U50 ( .IN1(n5), .IN2(input_mem_data[17]), .IN3(n6), .IN4(
        int_mem_data_rd[17]), .Q(N108) );
  AO22X1 U51 ( .IN1(n5), .IN2(input_mem_data[18]), .IN3(n6), .IN4(
        int_mem_data_rd[18]), .Q(N109) );
  AO22X1 U52 ( .IN1(n5), .IN2(input_mem_data[19]), .IN3(n6), .IN4(
        int_mem_data_rd[19]), .Q(N110) );
  AO22X1 U53 ( .IN1(n5), .IN2(input_mem_data[20]), .IN3(n6), .IN4(
        int_mem_data_rd[20]), .Q(N111) );
  AO22X1 U54 ( .IN1(n5), .IN2(input_mem_data[21]), .IN3(n6), .IN4(
        int_mem_data_rd[21]), .Q(N112) );
  AO22X1 U55 ( .IN1(n5), .IN2(input_mem_data[22]), .IN3(n6), .IN4(
        int_mem_data_rd[22]), .Q(N113) );
  AO22X1 U56 ( .IN1(n5), .IN2(input_mem_data[23]), .IN3(n6), .IN4(
        int_mem_data_rd[23]), .Q(N114) );
  AO22X1 U57 ( .IN1(n5), .IN2(input_mem_data[24]), .IN3(n6), .IN4(
        int_mem_data_rd[24]), .Q(N115) );
  AO22X1 U58 ( .IN1(n5), .IN2(input_mem_data[25]), .IN3(n6), .IN4(
        int_mem_data_rd[25]), .Q(N116) );
  AO22X1 U59 ( .IN1(n5), .IN2(input_mem_data[26]), .IN3(n6), .IN4(
        int_mem_data_rd[26]), .Q(N117) );
  AO22X1 U60 ( .IN1(n5), .IN2(input_mem_data[27]), .IN3(n6), .IN4(
        int_mem_data_rd[27]), .Q(N118) );
  AO22X1 U61 ( .IN1(n5), .IN2(input_mem_data[28]), .IN3(n6), .IN4(
        int_mem_data_rd[28]), .Q(N119) );
  AO22X1 U62 ( .IN1(n5), .IN2(input_mem_data[29]), .IN3(n6), .IN4(
        int_mem_data_rd[29]), .Q(N120) );
  AO22X1 U63 ( .IN1(n5), .IN2(input_mem_data[30]), .IN3(n6), .IN4(
        int_mem_data_rd[30]), .Q(N121) );
  AO22X1 U64 ( .IN1(n5), .IN2(input_mem_data[31]), .IN3(n6), .IN4(
        int_mem_data_rd[31]), .Q(N122) );
  AND2X1 U65 ( .IN1(w_data[0]), .IN2(n11), .Q(N126) );
  AND2X1 U66 ( .IN1(w_data[1]), .IN2(n11), .Q(N127) );
  AND2X1 U67 ( .IN1(w_data[2]), .IN2(n11), .Q(N128) );
  AND2X1 U68 ( .IN1(w_data[3]), .IN2(n11), .Q(N129) );
  AND2X1 U69 ( .IN1(w_data[4]), .IN2(n11), .Q(N130) );
  AND2X1 U70 ( .IN1(w_data[5]), .IN2(n11), .Q(N131) );
  AND2X1 U71 ( .IN1(w_data[6]), .IN2(n11), .Q(N132) );
  AND2X1 U72 ( .IN1(w_data[7]), .IN2(n11), .Q(N133) );
  AND2X1 U73 ( .IN1(w_data[8]), .IN2(n11), .Q(N134) );
  AND2X1 U74 ( .IN1(w_data[9]), .IN2(n11), .Q(N135) );
  AND2X1 U75 ( .IN1(w_data[10]), .IN2(n11), .Q(N136) );
  AND2X1 U76 ( .IN1(w_data[11]), .IN2(n11), .Q(N137) );
  AND2X1 U77 ( .IN1(w_data[12]), .IN2(n11), .Q(N138) );
  AND2X1 U78 ( .IN1(w_data[13]), .IN2(n11), .Q(N139) );
  AND2X1 U79 ( .IN1(w_data[14]), .IN2(n11), .Q(N140) );
  AND2X1 U80 ( .IN1(w_data[15]), .IN2(n11), .Q(N141) );
  AND2X1 U81 ( .IN1(w_data[16]), .IN2(n11), .Q(N142) );
  AND2X1 U82 ( .IN1(w_data[17]), .IN2(n11), .Q(N143) );
  AND2X1 U83 ( .IN1(w_data[18]), .IN2(n11), .Q(N144) );
  AND2X1 U84 ( .IN1(w_data[19]), .IN2(n11), .Q(N145) );
  AND2X1 U85 ( .IN1(w_data[20]), .IN2(n11), .Q(N146) );
  AND2X1 U86 ( .IN1(w_data[21]), .IN2(n11), .Q(N147) );
  AND2X1 U87 ( .IN1(w_data[22]), .IN2(n11), .Q(N148) );
  AND2X1 U88 ( .IN1(w_data[23]), .IN2(n11), .Q(N149) );
  AND2X1 U89 ( .IN1(w_data[24]), .IN2(n11), .Q(N150) );
  AND2X1 U90 ( .IN1(w_data[25]), .IN2(n11), .Q(N151) );
  AND2X1 U91 ( .IN1(w_data[26]), .IN2(n11), .Q(N152) );
  AND2X1 U92 ( .IN1(w_data[27]), .IN2(n11), .Q(N153) );
  AND2X1 U93 ( .IN1(w_data[28]), .IN2(n11), .Q(N154) );
  AND2X1 U94 ( .IN1(w_data[29]), .IN2(n11), .Q(N155) );
  AND2X1 U95 ( .IN1(w_data[30]), .IN2(n11), .Q(N156) );
  AND2X1 U96 ( .IN1(w_data[31]), .IN2(n11), .Q(N157) );
  MUX21X1 U97 ( .IN1(input_act_func[0]), .IN2(mac_output[0]), .S(ena_act_func), 
        .Q(N160) );
  MUX21X1 U98 ( .IN1(input_act_func[1]), .IN2(mac_output[1]), .S(ena_act_func), 
        .Q(N161) );
  MUX21X1 U99 ( .IN1(input_act_func[2]), .IN2(mac_output[2]), .S(ena_act_func), 
        .Q(N162) );
  MUX21X1 U100 ( .IN1(input_act_func[3]), .IN2(mac_output[3]), .S(ena_act_func), .Q(N163) );
  MUX21X1 U101 ( .IN1(input_act_func[4]), .IN2(mac_output[4]), .S(ena_act_func), .Q(N164) );
  MUX21X1 U102 ( .IN1(input_act_func[5]), .IN2(mac_output[5]), .S(n14), .Q(
        N165) );
  MUX21X1 U103 ( .IN1(input_act_func[6]), .IN2(mac_output[6]), .S(ena_act_func), .Q(N166) );
  MUX21X1 U104 ( .IN1(input_act_func[7]), .IN2(mac_output[7]), .S(ena_act_func), .Q(N167) );
  MUX21X1 U105 ( .IN1(input_act_func[8]), .IN2(mac_output[8]), .S(ena_act_func), .Q(N168) );
  MUX21X1 U106 ( .IN1(input_act_func[9]), .IN2(mac_output[9]), .S(ena_act_func), .Q(N169) );
  MUX21X1 U107 ( .IN1(input_act_func[10]), .IN2(mac_output[10]), .S(
        ena_act_func), .Q(N170) );
  MUX21X1 U108 ( .IN1(input_act_func[11]), .IN2(mac_output[11]), .S(n14), .Q(
        N171) );
  MUX21X1 U109 ( .IN1(input_act_func[12]), .IN2(mac_output[12]), .S(
        ena_act_func), .Q(N172) );
  MUX21X1 U110 ( .IN1(input_act_func[13]), .IN2(mac_output[13]), .S(n14), .Q(
        N173) );
  MUX21X1 U111 ( .IN1(input_act_func[14]), .IN2(mac_output[14]), .S(n14), .Q(
        N174) );
  MUX21X1 U112 ( .IN1(input_act_func[15]), .IN2(mac_output[15]), .S(
        ena_act_func), .Q(N175) );
  MUX21X1 U113 ( .IN1(input_act_func[16]), .IN2(mac_output[16]), .S(
        ena_act_func), .Q(N176) );
  MUX21X1 U114 ( .IN1(input_act_func[17]), .IN2(mac_output[17]), .S(
        ena_act_func), .Q(N177) );
  MUX21X1 U115 ( .IN1(input_act_func[18]), .IN2(mac_output[18]), .S(
        ena_act_func), .Q(N178) );
  MUX21X1 U116 ( .IN1(input_act_func[19]), .IN2(mac_output[19]), .S(n14), .Q(
        N179) );
  MUX21X1 U117 ( .IN1(input_act_func[20]), .IN2(mac_output[20]), .S(n14), .Q(
        N180) );
  MUX21X1 U118 ( .IN1(input_act_func[21]), .IN2(mac_output[21]), .S(n14), .Q(
        N181) );
  MUX21X1 U119 ( .IN1(input_act_func[22]), .IN2(mac_output[22]), .S(
        ena_act_func), .Q(N182) );
  MUX21X1 U120 ( .IN1(input_act_func[23]), .IN2(mac_output[23]), .S(
        ena_act_func), .Q(N183) );
  MUX21X1 U121 ( .IN1(input_act_func[24]), .IN2(mac_output[24]), .S(n14), .Q(
        N184) );
  MUX21X1 U122 ( .IN1(input_act_func[25]), .IN2(mac_output[25]), .S(n14), .Q(
        N185) );
  MUX21X1 U123 ( .IN1(input_act_func[26]), .IN2(mac_output[26]), .S(n14), .Q(
        N186) );
  MUX21X1 U124 ( .IN1(input_act_func[27]), .IN2(mac_output[27]), .S(n14), .Q(
        N187) );
  MUX21X1 U125 ( .IN1(input_act_func[28]), .IN2(mac_output[28]), .S(n14), .Q(
        N188) );
  MUX21X1 U126 ( .IN1(input_act_func[29]), .IN2(mac_output[29]), .S(n14), .Q(
        N189) );
  MUX21X1 U127 ( .IN1(input_act_func[30]), .IN2(mac_output[30]), .S(n14), .Q(
        N190) );
  MUX21X1 U128 ( .IN1(input_act_func[31]), .IN2(mac_output[31]), .S(n14), .Q(
        N191) );
  NOR2X0 U129 ( .IN1(n14), .IN2(n13), .QN(n17) );
  INVX0 U130 ( .INP(n17), .ZN(n18) );
  NOR2X0 U131 ( .IN1(act_function_sel[1]), .IN2(n17), .QN(n19) );
  AO222X1 U132 ( .IN1(n7), .IN2(sigmoid_output[0]), .IN3(n43), .IN4(
        linear_output[0]), .IN5(n42), .IN6(tansigmoid_output[0]), .Q(N235) );
  AO222X1 U133 ( .IN1(n7), .IN2(sigmoid_output[1]), .IN3(n43), .IN4(
        linear_output[1]), .IN5(n42), .IN6(tansigmoid_output[1]), .Q(N236) );
  AO222X1 U134 ( .IN1(n7), .IN2(sigmoid_output[2]), .IN3(n43), .IN4(
        linear_output[2]), .IN5(n42), .IN6(tansigmoid_output[2]), .Q(N237) );
  AO222X1 U135 ( .IN1(n7), .IN2(sigmoid_output[3]), .IN3(n43), .IN4(
        linear_output[3]), .IN5(n42), .IN6(tansigmoid_output[3]), .Q(N238) );
  AO222X1 U136 ( .IN1(n7), .IN2(sigmoid_output[4]), .IN3(n43), .IN4(
        linear_output[4]), .IN5(n42), .IN6(tansigmoid_output[4]), .Q(N239) );
  AO222X1 U137 ( .IN1(n7), .IN2(sigmoid_output[5]), .IN3(n43), .IN4(
        linear_output[5]), .IN5(n42), .IN6(tansigmoid_output[5]), .Q(N240) );
  AO222X1 U138 ( .IN1(n7), .IN2(sigmoid_output[6]), .IN3(n43), .IN4(
        linear_output[6]), .IN5(n42), .IN6(tansigmoid_output[6]), .Q(N241) );
  AO222X1 U139 ( .IN1(n7), .IN2(sigmoid_output[7]), .IN3(n43), .IN4(
        linear_output[7]), .IN5(n42), .IN6(tansigmoid_output[7]), .Q(N242) );
  AO222X1 U140 ( .IN1(n7), .IN2(sigmoid_output[8]), .IN3(n43), .IN4(
        linear_output[8]), .IN5(n42), .IN6(tansigmoid_output[8]), .Q(N243) );
  AO222X1 U141 ( .IN1(n7), .IN2(sigmoid_output[9]), .IN3(n43), .IN4(
        linear_output[9]), .IN5(n42), .IN6(tansigmoid_output[9]), .Q(N244) );
  AO222X1 U142 ( .IN1(n7), .IN2(sigmoid_output[10]), .IN3(n43), .IN4(
        linear_output[10]), .IN5(n42), .IN6(tansigmoid_output[10]), .Q(N245)
         );
  AO222X1 U143 ( .IN1(n7), .IN2(sigmoid_output[11]), .IN3(n43), .IN4(
        linear_output[11]), .IN5(n42), .IN6(tansigmoid_output[11]), .Q(N246)
         );
  AO222X1 U144 ( .IN1(n7), .IN2(sigmoid_output[12]), .IN3(n43), .IN4(
        linear_output[12]), .IN5(n42), .IN6(tansigmoid_output[12]), .Q(N247)
         );
  AO222X1 U145 ( .IN1(n7), .IN2(sigmoid_output[13]), .IN3(n43), .IN4(
        linear_output[13]), .IN5(n42), .IN6(tansigmoid_output[13]), .Q(N248)
         );
  AO222X1 U146 ( .IN1(n7), .IN2(sigmoid_output[14]), .IN3(n43), .IN4(
        linear_output[14]), .IN5(n42), .IN6(tansigmoid_output[14]), .Q(N249)
         );
  AO222X1 U147 ( .IN1(n7), .IN2(sigmoid_output[15]), .IN3(n43), .IN4(
        linear_output[15]), .IN5(n42), .IN6(tansigmoid_output[15]), .Q(N250)
         );
  AO222X1 U148 ( .IN1(n7), .IN2(sigmoid_output[16]), .IN3(n43), .IN4(
        linear_output[16]), .IN5(n42), .IN6(tansigmoid_output[16]), .Q(N251)
         );
  AO222X1 U149 ( .IN1(n7), .IN2(sigmoid_output[17]), .IN3(n43), .IN4(
        linear_output[17]), .IN5(n42), .IN6(tansigmoid_output[17]), .Q(N252)
         );
  AO222X1 U150 ( .IN1(n7), .IN2(sigmoid_output[18]), .IN3(n43), .IN4(
        linear_output[18]), .IN5(n42), .IN6(tansigmoid_output[18]), .Q(N253)
         );
  AO222X1 U151 ( .IN1(n7), .IN2(sigmoid_output[19]), .IN3(n43), .IN4(
        linear_output[19]), .IN5(n42), .IN6(tansigmoid_output[19]), .Q(N254)
         );
  AO222X1 U152 ( .IN1(n7), .IN2(sigmoid_output[20]), .IN3(n43), .IN4(
        linear_output[20]), .IN5(n42), .IN6(tansigmoid_output[20]), .Q(N255)
         );
  AO222X1 U153 ( .IN1(n7), .IN2(sigmoid_output[21]), .IN3(n43), .IN4(
        linear_output[21]), .IN5(n42), .IN6(tansigmoid_output[21]), .Q(N256)
         );
  AO222X1 U154 ( .IN1(n7), .IN2(sigmoid_output[22]), .IN3(n43), .IN4(
        linear_output[22]), .IN5(n42), .IN6(tansigmoid_output[22]), .Q(N257)
         );
  NAND3X0 U155 ( .IN1(n19), .IN2(step_output_23_), .IN3(n8), .QN(n41) );
  NAND4X0 U156 ( .IN1(n41), .IN2(n22), .IN3(n21), .IN4(n20), .QN(N258) );
  NAND4X0 U157 ( .IN1(n41), .IN2(n25), .IN3(n24), .IN4(n23), .QN(N259) );
  NAND4X0 U158 ( .IN1(n41), .IN2(n28), .IN3(n27), .IN4(n26), .QN(N260) );
  NAND4X0 U159 ( .IN1(n41), .IN2(n31), .IN3(n30), .IN4(n29), .QN(N261) );
  NAND4X0 U160 ( .IN1(n41), .IN2(n34), .IN3(n33), .IN4(n32), .QN(N262) );
  NAND4X0 U161 ( .IN1(n41), .IN2(n37), .IN3(n36), .IN4(n35), .QN(N263) );
  NAND4X0 U162 ( .IN1(n41), .IN2(n40), .IN3(n39), .IN4(n38), .QN(N264) );
  AO222X1 U163 ( .IN1(n7), .IN2(sigmoid_output[31]), .IN3(n43), .IN4(
        linear_output[31]), .IN5(n42), .IN6(tansigmoid_output[31]), .Q(N266)
         );
  MUX21X1 U164 ( .IN1(int_mem_data_wr[0]), .IN2(out_act_func[0]), .S(n13), .Q(
        N272) );
  MUX21X1 U165 ( .IN1(int_mem_data_wr[1]), .IN2(out_act_func[1]), .S(n13), .Q(
        N273) );
  MUX21X1 U166 ( .IN1(int_mem_data_wr[2]), .IN2(out_act_func[2]), .S(n13), .Q(
        N274) );
  MUX21X1 U167 ( .IN1(int_mem_data_wr[3]), .IN2(out_act_func[3]), .S(n13), .Q(
        N275) );
  MUX21X1 U168 ( .IN1(int_mem_data_wr[4]), .IN2(out_act_func[4]), .S(n13), .Q(
        N276) );
  MUX21X1 U169 ( .IN1(int_mem_data_wr[5]), .IN2(out_act_func[5]), .S(n13), .Q(
        N277) );
  MUX21X1 U170 ( .IN1(int_mem_data_wr[6]), .IN2(out_act_func[6]), .S(n13), .Q(
        N278) );
  MUX21X1 U171 ( .IN1(int_mem_data_wr[7]), .IN2(out_act_func[7]), .S(n13), .Q(
        N279) );
  MUX21X1 U172 ( .IN1(int_mem_data_wr[8]), .IN2(out_act_func[8]), .S(n53), .Q(
        N280) );
  MUX21X1 U173 ( .IN1(int_mem_data_wr[9]), .IN2(out_act_func[9]), .S(n53), .Q(
        N281) );
  MUX21X1 U174 ( .IN1(int_mem_data_wr[10]), .IN2(out_act_func[10]), .S(n53), 
        .Q(N282) );
  MUX21X1 U175 ( .IN1(int_mem_data_wr[11]), .IN2(out_act_func[11]), .S(n53), 
        .Q(N283) );
  MUX21X1 U176 ( .IN1(int_mem_data_wr[12]), .IN2(out_act_func[12]), .S(n53), 
        .Q(N284) );
  MUX21X1 U177 ( .IN1(int_mem_data_wr[13]), .IN2(out_act_func[13]), .S(n53), 
        .Q(N285) );
  MUX21X1 U178 ( .IN1(int_mem_data_wr[14]), .IN2(out_act_func[14]), .S(n53), 
        .Q(N286) );
  MUX21X1 U179 ( .IN1(int_mem_data_wr[15]), .IN2(out_act_func[15]), .S(n53), 
        .Q(N287) );
  MUX21X1 U180 ( .IN1(int_mem_data_wr[16]), .IN2(out_act_func[16]), .S(n53), 
        .Q(N288) );
  MUX21X1 U181 ( .IN1(int_mem_data_wr[17]), .IN2(out_act_func[17]), .S(n53), 
        .Q(N289) );
  MUX21X1 U182 ( .IN1(int_mem_data_wr[18]), .IN2(out_act_func[18]), .S(n53), 
        .Q(N290) );
  MUX21X1 U183 ( .IN1(int_mem_data_wr[19]), .IN2(out_act_func[19]), .S(n13), 
        .Q(N291) );
  MUX21X1 U184 ( .IN1(int_mem_data_wr[20]), .IN2(out_act_func[20]), .S(n13), 
        .Q(N292) );
  MUX21X1 U185 ( .IN1(int_mem_data_wr[21]), .IN2(out_act_func[21]), .S(n13), 
        .Q(N293) );
  MUX21X1 U186 ( .IN1(int_mem_data_wr[22]), .IN2(out_act_func[22]), .S(n13), 
        .Q(N294) );
  MUX21X1 U187 ( .IN1(int_mem_data_wr[23]), .IN2(out_act_func[23]), .S(n13), 
        .Q(N295) );
  MUX21X1 U188 ( .IN1(int_mem_data_wr[24]), .IN2(out_act_func[24]), .S(n13), 
        .Q(N296) );
  MUX21X1 U189 ( .IN1(int_mem_data_wr[25]), .IN2(out_act_func[25]), .S(n53), 
        .Q(N297) );
  MUX21X1 U190 ( .IN1(int_mem_data_wr[26]), .IN2(out_act_func[26]), .S(n53), 
        .Q(N298) );
  MUX21X1 U191 ( .IN1(int_mem_data_wr[27]), .IN2(out_act_func[27]), .S(n53), 
        .Q(N299) );
  MUX21X1 U192 ( .IN1(int_mem_data_wr[28]), .IN2(out_act_func[28]), .S(n53), 
        .Q(N300) );
  MUX21X1 U193 ( .IN1(int_mem_data_wr[29]), .IN2(out_act_func[29]), .S(n53), 
        .Q(N301) );
  MUX21X1 U194 ( .IN1(int_mem_data_wr[30]), .IN2(out_act_func[30]), .S(n53), 
        .Q(N302) );
  MUX21X1 U195 ( .IN1(int_mem_data_wr[31]), .IN2(out_act_func[31]), .S(n53), 
        .Q(N303) );
  MUX21X1 U196 ( .IN1(out_act_func[0]), .IN2(output_data[0]), .S(n44), .Q(N307) );
  MUX21X1 U197 ( .IN1(out_act_func[1]), .IN2(output_data[1]), .S(n44), .Q(N308) );
  MUX21X1 U198 ( .IN1(out_act_func[2]), .IN2(output_data[2]), .S(n44), .Q(N309) );
  MUX21X1 U199 ( .IN1(out_act_func[3]), .IN2(output_data[3]), .S(n44), .Q(N310) );
  MUX21X1 U200 ( .IN1(out_act_func[4]), .IN2(output_data[4]), .S(n44), .Q(N311) );
  MUX21X1 U201 ( .IN1(out_act_func[5]), .IN2(output_data[5]), .S(n44), .Q(N312) );
  MUX21X1 U202 ( .IN1(out_act_func[6]), .IN2(output_data[6]), .S(n44), .Q(N313) );
  MUX21X1 U203 ( .IN1(out_act_func[7]), .IN2(output_data[7]), .S(n44), .Q(N314) );
  MUX21X1 U204 ( .IN1(out_act_func[8]), .IN2(output_data[8]), .S(n44), .Q(N315) );
  MUX21X1 U205 ( .IN1(out_act_func[9]), .IN2(output_data[9]), .S(n12), .Q(N316) );
  MUX21X1 U206 ( .IN1(out_act_func[10]), .IN2(output_data[10]), .S(n12), .Q(
        N317) );
  MUX21X1 U207 ( .IN1(out_act_func[11]), .IN2(output_data[11]), .S(n12), .Q(
        N318) );
  MUX21X1 U208 ( .IN1(out_act_func[12]), .IN2(output_data[12]), .S(n12), .Q(
        N319) );
  MUX21X1 U209 ( .IN1(out_act_func[13]), .IN2(output_data[13]), .S(n12), .Q(
        N320) );
  MUX21X1 U210 ( .IN1(out_act_func[14]), .IN2(output_data[14]), .S(n12), .Q(
        N321) );
  MUX21X1 U211 ( .IN1(out_act_func[15]), .IN2(output_data[15]), .S(n12), .Q(
        N322) );
  MUX21X1 U212 ( .IN1(out_act_func[16]), .IN2(output_data[16]), .S(n12), .Q(
        N323) );
  MUX21X1 U213 ( .IN1(out_act_func[17]), .IN2(output_data[17]), .S(n12), .Q(
        N324) );
  MUX21X1 U214 ( .IN1(out_act_func[18]), .IN2(output_data[18]), .S(n12), .Q(
        N325) );
  MUX21X1 U215 ( .IN1(out_act_func[19]), .IN2(output_data[19]), .S(n12), .Q(
        N326) );
  MUX21X1 U216 ( .IN1(out_act_func[20]), .IN2(output_data[20]), .S(n12), .Q(
        N327) );
  MUX21X1 U217 ( .IN1(out_act_func[21]), .IN2(output_data[21]), .S(n12), .Q(
        N328) );
  MUX21X1 U218 ( .IN1(out_act_func[22]), .IN2(output_data[22]), .S(n12), .Q(
        N329) );
  MUX21X1 U219 ( .IN1(out_act_func[23]), .IN2(output_data[23]), .S(n12), .Q(
        N330) );
  MUX21X1 U220 ( .IN1(out_act_func[24]), .IN2(output_data[24]), .S(n12), .Q(
        N331) );
  MUX21X1 U221 ( .IN1(out_act_func[25]), .IN2(output_data[25]), .S(n12), .Q(
        N332) );
  MUX21X1 U222 ( .IN1(out_act_func[26]), .IN2(output_data[26]), .S(n12), .Q(
        N333) );
  MUX21X1 U223 ( .IN1(out_act_func[27]), .IN2(output_data[27]), .S(n12), .Q(
        N334) );
  MUX21X1 U224 ( .IN1(out_act_func[28]), .IN2(output_data[28]), .S(n12), .Q(
        N335) );
  MUX21X1 U225 ( .IN1(out_act_func[29]), .IN2(output_data[29]), .S(n12), .Q(
        N336) );
  MUX21X1 U226 ( .IN1(out_act_func[30]), .IN2(output_data[30]), .S(n12), .Q(
        N337) );
  MUX21X1 U227 ( .IN1(out_act_func[31]), .IN2(output_data[31]), .S(n12), .Q(
        N338) );
  NOR2X0 U228 ( .IN1(para_cof[3]), .IN2(para_cof[2]), .QN(n47) );
  INVX0 U229 ( .INP(para_cof[1]), .ZN(n51) );
  NAND4X0 U230 ( .IN1(input_or_int_mem_sel), .IN2(para_cof[0]), .IN3(n47), 
        .IN4(n51), .QN(n45) );
  MUX21X1 U231 ( .IN1(para_data[0]), .IN2(num_of_layer[0]), .S(n45), .Q(N347)
         );
  MUX21X1 U232 ( .IN1(para_data[1]), .IN2(num_of_layer[1]), .S(n45), .Q(N348)
         );
  MUX21X1 U233 ( .IN1(para_data[2]), .IN2(num_of_layer[2]), .S(n45), .Q(N349)
         );
  MUX21X1 U234 ( .IN1(para_data[3]), .IN2(num_of_layer[3]), .S(n45), .Q(N350)
         );
  INVX0 U235 ( .INP(para_cof[0]), .ZN(n50) );
  MUX21X1 U236 ( .IN1(para_data[0]), .IN2(mac_time[0]), .S(n46), .Q(N351) );
  MUX21X1 U237 ( .IN1(para_data[1]), .IN2(mac_time[1]), .S(n46), .Q(N352) );
  MUX21X1 U238 ( .IN1(para_data[2]), .IN2(mac_time[2]), .S(n46), .Q(N353) );
  MUX21X1 U239 ( .IN1(para_data[3]), .IN2(mac_time[3]), .S(n46), .Q(N354) );
  MUX21X1 U240 ( .IN1(para_data[4]), .IN2(mac_time[4]), .S(n46), .Q(N355) );
  MUX21X1 U241 ( .IN1(para_data[5]), .IN2(mac_time[5]), .S(n46), .Q(N356) );
  MUX21X1 U242 ( .IN1(para_data[6]), .IN2(mac_time[6]), .S(n46), .Q(N357) );
  MUX21X1 U243 ( .IN1(para_data[7]), .IN2(mac_time[7]), .S(n46), .Q(N358) );
  MUX21X1 U244 ( .IN1(para_data[8]), .IN2(mac_time[8]), .S(n46), .Q(N359) );
  MUX21X1 U245 ( .IN1(para_data[9]), .IN2(mac_time[9]), .S(n46), .Q(N360) );
  MUX21X1 U246 ( .IN1(para_data[10]), .IN2(mac_time[10]), .S(n46), .Q(N361) );
  MUX21X1 U247 ( .IN1(para_data[11]), .IN2(mac_time[11]), .S(n46), .Q(N362) );
  NAND3X0 U248 ( .IN1(para_cof[1]), .IN2(para_cof[0]), .IN3(n47), .QN(n48) );
  MUX21X1 U249 ( .IN1(para_data[0]), .IN2(num_of_node_for_each_layer[0]), .S(
        n48), .Q(N363) );
  MUX21X1 U250 ( .IN1(para_data[1]), .IN2(num_of_node_for_each_layer[1]), .S(
        n48), .Q(N364) );
  MUX21X1 U251 ( .IN1(para_data[2]), .IN2(num_of_node_for_each_layer[2]), .S(
        n48), .Q(N365) );
  MUX21X1 U252 ( .IN1(para_data[3]), .IN2(num_of_node_for_each_layer[3]), .S(
        n48), .Q(N366) );
  MUX21X1 U253 ( .IN1(para_data[4]), .IN2(num_of_node_for_each_layer[4]), .S(
        n48), .Q(N367) );
  MUX21X1 U254 ( .IN1(para_data[5]), .IN2(num_of_node_for_each_layer[5]), .S(
        n48), .Q(N368) );
  MUX21X1 U255 ( .IN1(para_data[6]), .IN2(num_of_node_for_each_layer[6]), .S(
        n48), .Q(N369) );
  MUX21X1 U256 ( .IN1(para_data[7]), .IN2(num_of_node_for_each_layer[7]), .S(
        n48), .Q(N370) );
  INVX0 U257 ( .INP(para_cof[3]), .ZN(n49) );
  NAND4X0 U258 ( .IN1(para_cof[2]), .IN2(n51), .IN3(n50), .IN4(n49), .QN(n52)
         );
  MUX21X1 U259 ( .IN1(para_data[0]), .IN2(act_function_sel[0]), .S(n52), .Q(
        N371) );
  MUX21X1 U260 ( .IN1(para_data[1]), .IN2(act_function_sel[1]), .S(n52), .Q(
        N372) );
  AO22X1 U261 ( .IN1(n5), .IN2(input_mem_data[0]), .IN3(n6), .IN4(
        int_mem_data_rd[0]), .Q(N91) );
  AO22X1 U262 ( .IN1(n5), .IN2(input_mem_data[1]), .IN3(n6), .IN4(
        int_mem_data_rd[1]), .Q(N92) );
  AO22X1 U263 ( .IN1(n5), .IN2(input_mem_data[2]), .IN3(n6), .IN4(
        int_mem_data_rd[2]), .Q(N93) );
  AO22X1 U264 ( .IN1(n5), .IN2(input_mem_data[3]), .IN3(n6), .IN4(
        int_mem_data_rd[3]), .Q(N94) );
  AO22X1 U265 ( .IN1(n5), .IN2(input_mem_data[4]), .IN3(n6), .IN4(
        int_mem_data_rd[4]), .Q(N95) );
  AO22X1 U266 ( .IN1(n5), .IN2(input_mem_data[5]), .IN3(n6), .IN4(
        int_mem_data_rd[5]), .Q(N96) );
  AO22X1 U267 ( .IN1(n5), .IN2(input_mem_data[6]), .IN3(n6), .IN4(
        int_mem_data_rd[6]), .Q(N97) );
  AO22X1 U268 ( .IN1(n5), .IN2(input_mem_data[7]), .IN3(n6), .IN4(
        int_mem_data_rd[7]), .Q(N98) );
  AO22X1 U269 ( .IN1(n5), .IN2(input_mem_data[8]), .IN3(n6), .IN4(
        int_mem_data_rd[8]), .Q(N99) );
endmodule


module top ( clk_sys, rst_n, ena_regconize, ena_checker, w_data, w_addr );
  input [31:0] w_data;
  output [19:0] w_addr;
  input clk_sys, rst_n, ena_regconize;
  output ena_checker;
  wire   wr_ena_n, wr_ena_out_n, SYNOPSYS_UNCONNECTED_1,
         SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3,
         SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5,
         SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7,
         SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9,
         SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11,
         SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13,
         SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15,
         SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17,
         SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19,
         SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21,
         SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_23,
         SYNOPSYS_UNCONNECTED_24, SYNOPSYS_UNCONNECTED_25,
         SYNOPSYS_UNCONNECTED_26, SYNOPSYS_UNCONNECTED_27,
         SYNOPSYS_UNCONNECTED_28, SYNOPSYS_UNCONNECTED_29,
         SYNOPSYS_UNCONNECTED_30, SYNOPSYS_UNCONNECTED_31,
         SYNOPSYS_UNCONNECTED_32, SYNOPSYS_UNCONNECTED_33,
         SYNOPSYS_UNCONNECTED_34, SYNOPSYS_UNCONNECTED_35,
         SYNOPSYS_UNCONNECTED_36, SYNOPSYS_UNCONNECTED_37,
         SYNOPSYS_UNCONNECTED_38, SYNOPSYS_UNCONNECTED_39,
         SYNOPSYS_UNCONNECTED_40, SYNOPSYS_UNCONNECTED_41,
         SYNOPSYS_UNCONNECTED_42, SYNOPSYS_UNCONNECTED_43,
         SYNOPSYS_UNCONNECTED_44, SYNOPSYS_UNCONNECTED_45,
         SYNOPSYS_UNCONNECTED_46, SYNOPSYS_UNCONNECTED_47,
         SYNOPSYS_UNCONNECTED_48, SYNOPSYS_UNCONNECTED_49,
         SYNOPSYS_UNCONNECTED_50, SYNOPSYS_UNCONNECTED_51,
         SYNOPSYS_UNCONNECTED_52, SYNOPSYS_UNCONNECTED_53,
         SYNOPSYS_UNCONNECTED_54, SYNOPSYS_UNCONNECTED_55,
         SYNOPSYS_UNCONNECTED_56, SYNOPSYS_UNCONNECTED_57,
         SYNOPSYS_UNCONNECTED_58, SYNOPSYS_UNCONNECTED_59,
         SYNOPSYS_UNCONNECTED_60, SYNOPSYS_UNCONNECTED_61,
         SYNOPSYS_UNCONNECTED_62, SYNOPSYS_UNCONNECTED_63,
         SYNOPSYS_UNCONNECTED_64, SYNOPSYS_UNCONNECTED_65,
         SYNOPSYS_UNCONNECTED_66, SYNOPSYS_UNCONNECTED_67,
         SYNOPSYS_UNCONNECTED_68, SYNOPSYS_UNCONNECTED_69,
         SYNOPSYS_UNCONNECTED_70, SYNOPSYS_UNCONNECTED_71,
         SYNOPSYS_UNCONNECTED_72, SYNOPSYS_UNCONNECTED_73,
         SYNOPSYS_UNCONNECTED_74, SYNOPSYS_UNCONNECTED_75,
         SYNOPSYS_UNCONNECTED_76, SYNOPSYS_UNCONNECTED_77,
         SYNOPSYS_UNCONNECTED_78, SYNOPSYS_UNCONNECTED_79,
         SYNOPSYS_UNCONNECTED_80;
  wire   [9:0] input_mem_addr;
  wire   [31:0] int_data;
  wire   [9:0] int_mem_wr_addr;
  wire   [31:0] int_mem_data_wr;
  wire   [9:0] para_addr;
  wire   [11:0] para_data;
  wire   [9:0] mem_out_addr;
  wire   [31:0] output_data;
  wire   [31:0] mfcc_data;

  mem_int mem_int_01 ( .clk(clk_sys), .addr_rd({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, input_mem_addr}), .wr_ena(wr_ena_n), 
        .data_rd(int_data), .addr_wr({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, int_mem_wr_addr}), .data_wr(int_mem_data_wr) );
  mem_interface mem_interface_01 ( .clk(clk_sys), .addr_rd({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, para_addr}), .wr_ena(
        wr_ena_out_n), .data_rd({SYNOPSYS_UNCONNECTED_1, 
        SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4, 
        SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, 
        SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, 
        SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11, 
        SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13, 
        SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, 
        SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17, 
        SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19, 
        SYNOPSYS_UNCONNECTED_20, para_data}), .addr_wr({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mem_out_addr}), .data_wr(
        output_data) );
  mem_mfcc mem_mfcc_01 ( .clk(clk_sys), .addr({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, input_mem_addr[8:0]}), .wr_ena(
        1'b0), .data(mfcc_data) );
  neural neural_01 ( .clk(clk_sys), .rst_n(rst_n), .enable_neural(
        ena_regconize), .disable_neural(ena_checker), .user_para_data({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, para_data}), 
        .user_para_addr({SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22, 
        SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24, 
        SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26, 
        SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28, 
        SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30, para_addr}), 
        .int_mem_addr_rd({SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32, 
        SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34, 
        SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36, 
        SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38, 
        SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40, 
        SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42, 
        SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44, 
        SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46, 
        SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48, 
        SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50}), .input_mem_addr({
        SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52, 
        SYNOPSYS_UNCONNECTED_53, SYNOPSYS_UNCONNECTED_54, 
        SYNOPSYS_UNCONNECTED_55, SYNOPSYS_UNCONNECTED_56, 
        SYNOPSYS_UNCONNECTED_57, SYNOPSYS_UNCONNECTED_58, 
        SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_60, input_mem_addr}), 
        .w_addr(w_addr), .int_mem_addr_wr({SYNOPSYS_UNCONNECTED_61, 
        SYNOPSYS_UNCONNECTED_62, SYNOPSYS_UNCONNECTED_63, 
        SYNOPSYS_UNCONNECTED_64, SYNOPSYS_UNCONNECTED_65, 
        SYNOPSYS_UNCONNECTED_66, SYNOPSYS_UNCONNECTED_67, 
        SYNOPSYS_UNCONNECTED_68, SYNOPSYS_UNCONNECTED_69, 
        SYNOPSYS_UNCONNECTED_70, int_mem_wr_addr}), .output_mem_addr({
        SYNOPSYS_UNCONNECTED_71, SYNOPSYS_UNCONNECTED_72, 
        SYNOPSYS_UNCONNECTED_73, SYNOPSYS_UNCONNECTED_74, 
        SYNOPSYS_UNCONNECTED_75, SYNOPSYS_UNCONNECTED_76, 
        SYNOPSYS_UNCONNECTED_77, SYNOPSYS_UNCONNECTED_78, 
        SYNOPSYS_UNCONNECTED_79, SYNOPSYS_UNCONNECTED_80, mem_out_addr}), 
        .int_mem_data_rd(int_data), .input_mem_data(mfcc_data), .w_data(w_data), .int_mem_data_wr(int_mem_data_wr), .output_data(output_data), 
        .wr_ena_int_n_BAR(wr_ena_n), .wr_ena_out_n_BAR(wr_ena_out_n) );
endmodule


module vr ( RST_N, PLL_CLOCK, ENA_RECOGNIZE, SRAM_DQ0, SRAM_DQ1, SRAM_DQ2, 
        SRAM_DQ3, SRAM_DQ4, SRAM_DQ5, SRAM_DQ6, SRAM_DQ7, SRAM_DQ8, SRAM_DQ9, 
        SRAM_DQ10, SRAM_DQ11, SRAM_DQ12, SRAM_DQ13, SRAM_DQ14, SRAM_DQ15, 
        SRAM_DQ16, SRAM_DQ17, SRAM_DQ18, SRAM_DQ19, SRAM_DQ20, SRAM_DQ21, 
        SRAM_DQ22, SRAM_DQ23, SRAM_DQ24, SRAM_DQ25, SRAM_DQ26, SRAM_DQ27, 
        SRAM_DQ28, SRAM_DQ29, SRAM_DQ30, SRAM_DQ31, SRAM_ADDR0, SRAM_ADDR1, 
        SRAM_ADDR2, SRAM_ADDR3, SRAM_ADDR4, SRAM_ADDR5, SRAM_ADDR6, SRAM_ADDR7, 
        SRAM_ADDR8, SRAM_ADDR9, SRAM_ADDR10, SRAM_ADDR11, SRAM_ADDR12, 
        SRAM_ADDR13, SRAM_ADDR14, SRAM_ADDR15, SRAM_ADDR16, SRAM_ADDR17, 
        SRAM_ADDR18, SRAM_ADDR19, ENA_CHECKER );
  input RST_N, PLL_CLOCK, ENA_RECOGNIZE, SRAM_DQ0, SRAM_DQ1, SRAM_DQ2,
         SRAM_DQ3, SRAM_DQ4, SRAM_DQ5, SRAM_DQ6, SRAM_DQ7, SRAM_DQ8, SRAM_DQ9,
         SRAM_DQ10, SRAM_DQ11, SRAM_DQ12, SRAM_DQ13, SRAM_DQ14, SRAM_DQ15,
         SRAM_DQ16, SRAM_DQ17, SRAM_DQ18, SRAM_DQ19, SRAM_DQ20, SRAM_DQ21,
         SRAM_DQ22, SRAM_DQ23, SRAM_DQ24, SRAM_DQ25, SRAM_DQ26, SRAM_DQ27,
         SRAM_DQ28, SRAM_DQ29, SRAM_DQ30, SRAM_DQ31;
  output SRAM_ADDR0, SRAM_ADDR1, SRAM_ADDR2, SRAM_ADDR3, SRAM_ADDR4,
         SRAM_ADDR5, SRAM_ADDR6, SRAM_ADDR7, SRAM_ADDR8, SRAM_ADDR9,
         SRAM_ADDR10, SRAM_ADDR11, SRAM_ADDR12, SRAM_ADDR13, SRAM_ADDR14,
         SRAM_ADDR15, SRAM_ADDR16, SRAM_ADDR17, SRAM_ADDR18, SRAM_ADDR19,
         ENA_CHECKER;
  wire   pll_clock, reset, ena_regconize, ena_checker;
  wire   [31:0] w_data;
  wire   [19:0] w_addr;
  tri   SRAM_ADDR0;
  tri   SRAM_ADDR1;
  tri   SRAM_ADDR2;
  tri   SRAM_ADDR3;
  tri   SRAM_ADDR4;
  tri   SRAM_ADDR5;
  tri   SRAM_ADDR6;
  tri   SRAM_ADDR7;
  tri   SRAM_ADDR8;
  tri   SRAM_ADDR9;
  tri   SRAM_ADDR10;
  tri   SRAM_ADDR11;
  tri   SRAM_ADDR12;
  tri   SRAM_ADDR13;
  tri   SRAM_ADDR14;
  tri   SRAM_ADDR15;
  tri   SRAM_ADDR16;
  tri   SRAM_ADDR17;
  tri   SRAM_ADDR18;
  tri   SRAM_ADDR19;
  tri   ENA_CHECKER;

  top top_01 ( .clk_sys(pll_clock), .rst_n(reset), .ena_regconize(
        ena_regconize), .ena_checker(ena_checker), .w_data(w_data), .w_addr(
        w_addr) );
  D2I1025 D2I1025_ENA_CHECKER ( .DIN(ena_checker), .EN(1'b1), .PADIO(
        ENA_CHECKER) );
  ISH1025 ISH1025_ENA_REG ( .PADIO(ENA_RECOGNIZE), .R_EN(1'b1), .DOUT(
        ena_regconize) );
  ISH1025 ISH1025_PRST_N ( .PADIO(RST_N), .R_EN(1'b1), .DOUT(reset) );
  ISH1025 ISH1025_PLL_CLOCK ( .PADIO(PLL_CLOCK), .R_EN(1'b1), .DOUT(pll_clock)
         );
  D2I1025 D2I1025_SRAM_ADD19 ( .DIN(w_addr[19]), .EN(1'b1), .PADIO(SRAM_ADDR19) );
  D2I1025 D2I1025_SRAM_ADD18 ( .DIN(w_addr[18]), .EN(1'b1), .PADIO(SRAM_ADDR18) );
  D2I1025 D2I1025_SRAM_ADD17 ( .DIN(w_addr[17]), .EN(1'b1), .PADIO(SRAM_ADDR17) );
  D2I1025 D2I1025_SRAM_ADD16 ( .DIN(w_addr[16]), .EN(1'b1), .PADIO(SRAM_ADDR16) );
  D2I1025 D2I1025_SRAM_ADD15 ( .DIN(w_addr[15]), .EN(1'b1), .PADIO(SRAM_ADDR15) );
  D2I1025 D2I1025_SRAM_ADD14 ( .DIN(w_addr[14]), .EN(1'b1), .PADIO(SRAM_ADDR14) );
  D2I1025 D2I1025_SRAM_ADD13 ( .DIN(w_addr[13]), .EN(1'b1), .PADIO(SRAM_ADDR13) );
  D2I1025 D2I1025_SRAM_ADD12 ( .DIN(w_addr[12]), .EN(1'b1), .PADIO(SRAM_ADDR12) );
  D2I1025 D2I1025_SRAM_ADD11 ( .DIN(w_addr[11]), .EN(1'b1), .PADIO(SRAM_ADDR11) );
  D2I1025 D2I1025_SRAM_ADD10 ( .DIN(w_addr[10]), .EN(1'b1), .PADIO(SRAM_ADDR10) );
  D2I1025 D2I1025_SRAM_ADD9 ( .DIN(w_addr[9]), .EN(1'b1), .PADIO(SRAM_ADDR9)
         );
  D2I1025 D2I1025_SRAM_ADD8 ( .DIN(w_addr[8]), .EN(1'b1), .PADIO(SRAM_ADDR8)
         );
  D2I1025 D2I1025_SRAM_ADD7 ( .DIN(w_addr[7]), .EN(1'b1), .PADIO(SRAM_ADDR7)
         );
  D2I1025 D2I1025_SRAM_ADD6 ( .DIN(w_addr[6]), .EN(1'b1), .PADIO(SRAM_ADDR6)
         );
  D2I1025 D2I1025_SRAM_ADD5 ( .DIN(w_addr[5]), .EN(1'b1), .PADIO(SRAM_ADDR5)
         );
  D2I1025 D2I1025_SRAM_ADD4 ( .DIN(w_addr[4]), .EN(1'b1), .PADIO(SRAM_ADDR4)
         );
  D2I1025 D2I1025_SRAM_ADD3 ( .DIN(w_addr[3]), .EN(1'b1), .PADIO(SRAM_ADDR3)
         );
  D2I1025 D2I1025_SRAM_ADD2 ( .DIN(w_addr[2]), .EN(1'b1), .PADIO(SRAM_ADDR2)
         );
  D2I1025 D2I1025_SRAM_ADD1 ( .DIN(w_addr[1]), .EN(1'b1), .PADIO(SRAM_ADDR1)
         );
  D2I1025 D2I1025_SRAM_ADD0 ( .DIN(w_addr[0]), .EN(1'b1), .PADIO(SRAM_ADDR0)
         );
  ISH1025 ISH1025_SRAM_DQ31 ( .PADIO(SRAM_DQ31), .R_EN(1'b1), .DOUT(w_data[31]) );
  ISH1025 ISH1025_SRAM_DQ30 ( .PADIO(SRAM_DQ30), .R_EN(1'b1), .DOUT(w_data[30]) );
  ISH1025 ISH1025_SRAM_DQ29 ( .PADIO(SRAM_DQ29), .R_EN(1'b1), .DOUT(w_data[29]) );
  ISH1025 ISH1025_SRAM_DQ28 ( .PADIO(SRAM_DQ28), .R_EN(1'b1), .DOUT(w_data[28]) );
  ISH1025 ISH1025_SRAM_DQ27 ( .PADIO(SRAM_DQ27), .R_EN(1'b1), .DOUT(w_data[27]) );
  ISH1025 ISH1025_SRAM_DQ26 ( .PADIO(SRAM_DQ26), .R_EN(1'b1), .DOUT(w_data[26]) );
  ISH1025 ISH1025_SRAM_DQ25 ( .PADIO(SRAM_DQ25), .R_EN(1'b1), .DOUT(w_data[25]) );
  ISH1025 ISH1025_SRAM_DQ24 ( .PADIO(SRAM_DQ24), .R_EN(1'b1), .DOUT(w_data[24]) );
  ISH1025 ISH1025_SRAM_DQ23 ( .PADIO(SRAM_DQ23), .R_EN(1'b1), .DOUT(w_data[23]) );
  ISH1025 ISH1025_SRAM_DQ22 ( .PADIO(SRAM_DQ22), .R_EN(1'b1), .DOUT(w_data[22]) );
  ISH1025 ISH1025_SRAM_DQ21 ( .PADIO(SRAM_DQ21), .R_EN(1'b1), .DOUT(w_data[21]) );
  ISH1025 ISH1025_SRAM_DQ20 ( .PADIO(SRAM_DQ20), .R_EN(1'b1), .DOUT(w_data[20]) );
  ISH1025 ISH1025_SRAM_DQ19 ( .PADIO(SRAM_DQ19), .R_EN(1'b1), .DOUT(w_data[19]) );
  ISH1025 ISH1025_SRAM_DQ18 ( .PADIO(SRAM_DQ18), .R_EN(1'b1), .DOUT(w_data[18]) );
  ISH1025 ISH1025_SRAM_DQ17 ( .PADIO(SRAM_DQ17), .R_EN(1'b1), .DOUT(w_data[17]) );
  ISH1025 ISH1025_SRAM_DQ16 ( .PADIO(SRAM_DQ16), .R_EN(1'b1), .DOUT(w_data[16]) );
  ISH1025 ISH1025_SRAM_DQ15 ( .PADIO(SRAM_DQ15), .R_EN(1'b1), .DOUT(w_data[15]) );
  ISH1025 ISH1025_SRAM_DQ14 ( .PADIO(SRAM_DQ14), .R_EN(1'b1), .DOUT(w_data[14]) );
  ISH1025 ISH1025_SRAM_DQ13 ( .PADIO(SRAM_DQ13), .R_EN(1'b1), .DOUT(w_data[13]) );
  ISH1025 ISH1025_SRAM_DQ12 ( .PADIO(SRAM_DQ12), .R_EN(1'b1), .DOUT(w_data[12]) );
  ISH1025 ISH1025_SRAM_DQ11 ( .PADIO(SRAM_DQ11), .R_EN(1'b1), .DOUT(w_data[11]) );
  ISH1025 ISH1025_SRAM_DQ10 ( .PADIO(SRAM_DQ10), .R_EN(1'b1), .DOUT(w_data[10]) );
  ISH1025 ISH1025_SRAM_DQ9 ( .PADIO(SRAM_DQ9), .R_EN(1'b1), .DOUT(w_data[9])
         );
  ISH1025 ISH1025_SRAM_DQ8 ( .PADIO(SRAM_DQ8), .R_EN(1'b1), .DOUT(w_data[8])
         );
  ISH1025 ISH1025_SRAM_DQ7 ( .PADIO(SRAM_DQ7), .R_EN(1'b1), .DOUT(w_data[7])
         );
  ISH1025 ISH1025_SRAM_DQ6 ( .PADIO(SRAM_DQ6), .R_EN(1'b1), .DOUT(w_data[6])
         );
  ISH1025 ISH1025_SRAM_DQ5 ( .PADIO(SRAM_DQ5), .R_EN(1'b1), .DOUT(w_data[5])
         );
  ISH1025 ISH1025_SRAM_DQ4 ( .PADIO(SRAM_DQ4), .R_EN(1'b1), .DOUT(w_data[4])
         );
  ISH1025 ISH1025_SRAM_DQ3 ( .PADIO(SRAM_DQ3), .R_EN(1'b1), .DOUT(w_data[3])
         );
  ISH1025 ISH1025_SRAM_DQ2 ( .PADIO(SRAM_DQ2), .R_EN(1'b1), .DOUT(w_data[2])
         );
  ISH1025 ISH1025_SRAM_DQ1 ( .PADIO(SRAM_DQ1), .R_EN(1'b1), .DOUT(w_data[1])
         );
  ISH1025 ISH1025_SRAM_DQ0 ( .PADIO(SRAM_DQ0), .R_EN(1'b1), .DOUT(w_data[0])
         );
endmodule

